��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_I
y��������k%̜S���9('�X�@�'�X��m+��G������g��d�:]�<'� F��-!�k(�M�u�=X͝c���/���A�l�8��'?nZ�]�,�u�������k��ᚘYڏ㑠ڲ]��L���s��F�N��o3KK�+^_o;�_3B���'���f��jI��j��ŪD����8��3֓��p�O�P�hD�����ץtT��Wp��ZӰ]1�b��#�A�H��,�n�ʫ�I|�_T#{i;��5�$mX��b�"�(���<�B��p�J�O"R���Cr�7몈K����r��K��ΐ*W�`� �s���2q���k1wA#���k�b>����8��0~XӋ�ub����?�\;VQ��!�o�U��u_3��7��"�o r��-�ڙ �j��}��q�4(��jbu�h�b)h:������d!$_���E��FH� �%��?�V��o��[M#ߕ�>*8N�5DIba��lm[����������)w�3����#Gk��y��~�*�s3��£�9�eC��>��U���.S���u�_��D��1#�����\'��v���O!��M�,$�* dM��Me쎶��ʧ<��p�9:�`��[5�^�`�e#5{���% [��Dnî�]���3^&�'���l�z�t3�B�Y�ׅ����r��Rc���O;#��#B�j�R�&@3|N'h���Jޒ�1��j���%�
�on�{�����}��.|"�R��.�ڮ�6��J���ℳ�l�\�jS�f=��LI�gh�k� ����4kUϮoe_�8������e�'vSO��Oh$'�8�`�y]5�lL�����w�Hb�%�u�B�:��dL�>N`k�\������Ǘ���'K.Rr��
�yIe��   խ��tW���b+^�U��`���wK�WMn
�Nf�ص�w�o߹/|{�Ƈ�
Uf$)1tF}�P̳ ��E�4ֶ?��v���$�wy~]����zY����DQA�1�j��e��A�����9K��-�Ms���U^v��V�������Y���4��]z5�N�,���F��[T���L��4]����$�|&ڿf�Җ�`��*s֗ n�����x.� C�+HM@=��ޞYS!��P�HK�f>���=�S��a-�MY���0�?����=
Pv�Y�$Ov5$�m���#'��W4��$o-X�ڱ�
�ew	H��C9�^Vo��C����
)�JM'3�&�N�z���Pbo�=6��>�$0�o*IP�f�q���P!�Bn��p��ؾ�~���������'��:X~v�1� ��Zc_�˹�H�<��pk��vK�$A��ڍ��y4� ���P��PX����:�z'[̊f��?!`]Z�o�sh,���<����;Z����q��?`	���(���� �4E�:)P��I ���l��(f*ͮ6�����������)�9��វ.�g��;j��o��3�ʭ"�I����lž�3y���K��>��#\P-�(,�	�qo�*@kS�	�v E��Em`���Ґhk���G�iŸ	���x?h�(�K��B��FdO��]�2�����4s߽�*�ysO.K*G.��w����p���/�`�������"h���@�Z��p��sSn���B����W{�7^��k�Lnc���X4��My����J�U顺�r��q ��$��5�3 ��+�=s	G�wN��>�B�a����?[�X�3��[��6:up����,���̈ߧL�Ô�m��r0���qϩ��a���PzU8��n�ڲp�:RS%u�j2����	�+X�3]9�aE ����$�m%9}ڣ<�2��0�m<D�	*��b�DB!&���=hs���)7l{r+v���𵍡5������H�ES�k���2C����%oV9C���	dU��-��ܵ+��_ݕ�"6��ǅ{�eɂ���-�k�u�.A���Y��Hjپ��y���rr�*Y������1��Vpz�k�Ρ�~�E��sEA+�k��V���Ͷ����O�WjA �ﭛ�KԱ
1X�?$$��@��-I���vTF��i򶘒�qlFB���'sYN�a��A#��Y�V恣J�Bz,�C���-�2g\1�D���.V�JWq���:����:9S��y!x��d��S �����`���Y��>��
 ��F���K˘䱠#'oemw�#�M�����H*( ��?o��uD����|pjxP�ˡbjfʞ��5��o[ܲ��?o��(�u�-�M����Ri�H+�%�g)^��}o��L�^�ɐ��� E�W�`܂<M�s(�t����[u՗`j��i�e�
w!�I�rf~��{��kL�^Ϝ��Rh:��D�\�.��u�q��!R�Aw��3��&�\�%���s/�E��.¥{�[�����9W�P���=�@/�<���_�Ղ(�h�_���wb� �{��;q�~��C������r�A'1A�1�g�y�=�w���R���Ȥ��/��OL���|��w
�oiR]���M�ˬ��ҦG�+�'r�nKؖ��A|�0�뢈䫄ӂ� �Id�����Ѥ��D�T1e- �G��\�����E�d�7�0�J���J�8�6�e��Kg���" ![횾��Xǃ�3��s�a+�?��EC_��ιhn����1��I�1�12-W�j�NT�LL��*Ip��6x�}�c۲o�`]Qữ���!3j�yf�Ȕ*w�d	�C���`F�S��p�gE���7�\|m�e�Bj0c��Y1���?�~��B���ksyK��i���3Z6�?����[����EޡWS�/w�?��U��c����B�!R֤��?��#�M�8�؜���F�;ybH�[:� ya�c;��.]�?#�%彆%��� ����¡�3�5��0��+�m��V�A3(��0�B�ږ?��2-рq]����!B�*+x�P�:ǫ�`&P傗�2�ꮺ���>X���XT�f�ݭ/XBD��_卷���J�v;�X-1�6?�##��.>tz/�bx�G�nij#C�����D��:7��������k\��Y��9X{�,��m�^ѩ�4��Z�����*�)��P��c��
�oe�z'��]q,fOqSg|!Q�ʐ[˙I�L�/SJ���"-��:. K�[�Y!2O�V2���C����FI��0ד@�WL<�@�\i�
���-O��&|V�ٍU�t��ȝ��8k�~����	��ql�&���4�����N}R���;H\M���/��䡂 ��p|Ѹf@���	��:��WV��ukwXU� �D��~G`B�� (b{mO�qi�.�'��	9i:Yp���bF�o�� Q��/��&�5�H��R(� �8�W���5�Dp������p�<ǩ�k�4ԧ�C*.��G��&�ENL�Ӽ���&��t�:���ߚ-&��r'&��U�ݷ>���@�������e�z���ݱx�-G�6�uqGE��^ƶI�>E�t�1Y��|��A�m�=�bg�
���d?)P$�^Tj�CӒ�QМ��I����#���>�NW�]?
 b��
��%�%F8C�C�a�I7UѲ��[���E�w�ҞH���TMqJN`x�+	S@��Ɍ2�~~8��a�%RKxW=�^f;�pm-�G&���ߩ��@Rs)����g��J�ý�.K���,p�rU����e�h,x!�tdi�:�%=iu�E޹�V�W2+B�2&�beE�X����A�r����QM���C�FMVx�/Mek$RxMu� �ED�o��T:�v������-���;��y��?���-$�"M0`F��-�x�HN��uvu�cP�j�F���w���xF���q(�6`���|�"��엣?�$	w�B̒�Q� �)��y}y��FiO���q>��L_�����p�l ��	O=�)����i�?K\�P���8Hꎈ�u��/$l�/�!�	�g�����X��
s٠\W�ia$�hT�^�׌k�V�iU�B{�k�\\����Fe&pj9���=ٓ3�d���YQ��qk-lD�Ȋ#���`^��R+�O!�tɡ"���Dp��+��O����&� �Q���f�Q�"Щ�j��te,P�2�"�f�c��5�a&Bf[����4U�h��0����.��?�-����|��ź ������9�[�h.��X�
�W�
�=�.m��B*�*�N��4Ɠ�?G�j׷'��ɞϠBR�|���	͹���)	��	zb�z�KI����X)~�]_R��q	
Z���S=;/�0TW��3�$i5o�􂲉��iV��X����
?E�K���_[�&2&���5t"
���e�֪���Ψ���Hn�!�u��Ġ��,�R�5tF{�-w�
\\b�MS����Jh�pi�0�#6����Z=T4�L��m|:ީ��X�:Gkc13hG���Ε`z�_��Ŏ'E�*���E������a�Ӱ�I�9e��R=�(KT'�)� ��D�r�����ɚ��X�bJR<��qG�=z�X+A�A��,��ʀA��ax��ۘO|���/÷ ��l��	θ��|	*@d�h����8����ޅ�AB#��?�ټ�[��^�4Dh�y���V�U��L��D�H��H}���a��|�)>�8�>��D��D~ݥ�(˾���m�lL����"�����\��fo���7l֞�c�`�DP�3�Q�����㡅d�� k�t��q�ܱ��/T��-�gsG>�c���;z��$�ʣVx�Η��,��G溵�Ib�����^n��Z� --���lDp�1�́EEOk7rm͇����ve`�$V~}�xH;��U�U��5�7�f>p������;G@ИM~[����pE�t+��+��*$4G�^v�1��GO��H��9ՙ������uz���_S��� ���F�-xb�T��(�g��FB������gQ3s�7\����%�0���|�?Y�t�a�7^o��\my����#m�[`�O��A'NbA��"z2i{��X��X�W���qL���0y�õ�ɯ՗р[ac���seA���*�*0f�9 &�|x�ޗ������#�m�M6��q�Ŀ��;Od�Ӟ�=I����[���y�K����;dv�M#�(�l��e �;7p̓'qL ��&�-�x(6��Fi��L&�t����Ưe��c�Z<R�9}�L�UsaЌhPF���~�勦�e��Zl���N�T<#:b8	�;���]�ۈ�T�
�h,�5��q�>Zy�ؤ����Rc����?]$D�x������U}��`�p���đ ݯ{�H�ΐP����+��Z.G1F[�%	���%LL
�Du�V�Y�uX��|��(cA�q���X�7�������}Rc�v"��V�q�z��R�!?;B_�*�T�!�}��F�ԟ_ULSet�dj��٧�㍤�&by��0��VN�4�޹��6��2�~=�e�R�f0���Ǥ�3������;���TF�b�*%�̐"�Zp�g\4��=�4E`eB��[FTv} �7\��m`�ɷuNy�G�AѤM-?�������N���"���B��I7-U��%�Ճ�73lCJ�-	�#r����E�>8L���Kj��V��7z�#C�M��Cb�'��l�V��H/_�o����Y�-O�m��n�k�.3�I��OV���!�PШԑ���j�׉m�9}S�ȓ�Ǎ�a�	9 �Y�4�-I�HP���xK�s��`���0w9$b�ܷެ֦�S"�E9��0ǽ�ua���w�|I?:@�*�p�#��a|�l Gգ��\�=b��W��{"w���_�����X��'��M�)���U,����s��ؚΘ�4�~��N��5���h�.cI�k �ZF}/&�ZW=���j�=\�F�H� �@n7��k�� qE����Q���r��.b��[��r�z��:]��o��:��N1#� q��W{��d��Y�q��{_�]�	��8�Cs;K�ҏ.ң$����y
�7�Z$��QE#������Q�s�U���#�,퓫�O���^�q�:*g�G=ψ�<_����H��ת��-1fA�B�&hI�7�:#w���d��9��l$�?4C�'*�C�թ�.�d��������b�]�ty��k��0�311p�������Q&V�#8��7��wf�
���Lf"?��ByMR�����2fJ&ϩ;#]Ge���$1o�h\,Tf*��-�U�Dw�C�h�'�Ԩ/X
h�� �9(��=��H���.�Ӭ�W���I�v�$�W�x@w��'�q��H�!��̆���¡J���xR6ZQ9�Ļ%�)]��3��[}�s^3�@��!y"V
&(���$CY��#A�$�z�$�"t�㷬\�x�1�	���.9��ȮBR�ο�k�߽
���~Xx\n� *�k��3n���?�;i�Aktb�Xm�MK�flHWUY���!�@*���nhݺ��◲N8M�d
t�o��f|I�&ڡ�'��[����0�;�����hh�pڥ�
�b�	&�B�]a�V��1.m9�
ں04�2C��c���~X��F���>��!RU��$��;of&��g��`�S��Y]�DTȚ��i�W�-��
�f�1�z[M'	B�U���{��ж�H�������NjY�����:	۳:�0�͛�%�Z�Ύ��I�4��O;�G��~���I�"w�~���U,��f?S����Q�(�~P��l����"�i��]�Z���^a�so�>��#���o���5�S�!ֺ
1��=���*�rJ��R��e��Ѷ߃��F
	�	<���o�mא��ٝp<Չ��W��;�H��;L�M�Q��N�bgc�t��=�:�x���dA�"
҆�5�o�:����{2�NT͒���I��]��-���4���?}C܍+��u��B�Jt���{��K������r寴���p��:��|8"+��������;�������9����GD��q�j4���D�L%�{�^����l-�~���;��n���0��<�C}ll	����R\��<~�
Jdn��/0�n�*���=iS(,`�Nafa��7�U@䇃����<�̅NȚ�?.W��ہ����,7�q	1ʁ�^�VWs? �D�8$�/8���.c���*�^�WY���+�~�7oQ0���QV�͎+������v�p (�㊜\�E%����"��)E�7;�[-�d�B�2�\73ưdW�k���� ��y���,�P���D�u���u ���G�����,g O��$�v�S�:���y�AYxp(ؖ#U~}.hI2!"��Ӭ�$u���3�=͋���CyL]�Dۂ����O6-��V���j������d�dJe�&2�g��8H.�����WW�-t��v[�~��Y�C����H��2���gs���u��G�^�*"g�ǭ�]�c�#忺>w��R�h��bA� ��̗�ŻrPC��墜A\�:����(�� 98k��e��'c�L���d�r���m�Ģ��
�k� ���@m��s��r�~�8��ٜ�@ߕao���4u��2!{�Mf ϒ����%�|hҁ�ɸD��h�gPݠ�B�YĄ�~���p:ۂn]cl�CU0-�V�*pMiǬ�/K��.��y&o@ʊ��TCl��N��/���l3h�}Q��t����,QW
��D��B��]��T�%��M+����}v o{��Ұ'[H�k7Πר�!���cO�ܱ�Pe�YK��>ٛ�V�Ƅ�8�Ӭ�7q�BJ�G
�O@Y}x���*�r�Ȼ	w��2�Z��8F� ��?.�"j���Ά|zk��=zV��Uy�x8��<��*|�1�y�2ݵ�b����+��ݲ��	5�3+s�8,��a�����Zn�_</�yo�UʐC���m�ڱ��^�5et�dРT,��{)ԗSĔ���N �\�
p�����ߘ�1	�fYX�Ol��ݵל����#5j��)��	,��ܔ�[�e�1�W��bw��sxm�=:~I�iP�'���؍Qjs�m��e�
���� �&�Y��F���v�7�>v�1
�ux��$��s�3N�V��컺�Uw$P(uP�^���pPd�@0���E	�P�^V���n:��)��eh�I�F�ן�t�j췸�M���>������B�@M�i�p�V#�~�X4���)��o�����iGK���5�B
]�#�/f���͟�O�Iv )xzu�Ox �.�/�Wr����uF�Cw�}N�+�W�\��K�����#'D��!zJ�A(���X�\�LDr��52 �iVDp�Aݘ�`�J?�Ph(-�^�^jE�'r���,�8�|
��H �2j�}~�WK�#�eA첦$�sD.3Y�,�=9�mb��������K�ك�A��[�I�h��U��ZSc��_�����8y,C�0u{{�_�����bX�q{V���2m���̒lX�W�j7�/��`�GW)z1��W��2<
~�����W��A�J�{|�\@&b�� ��Ǉ�x{̀�?'�����LQ�B�3��v��dı+&hWF��gT�m��9~��lqt�d�M#�>�	��
��V>�����g�Dw�?�����Q�h�1�x[��~�����s�+�<��c8����k�X
���\[` �O��.�y������2 �T�0�j�|�9p���=jR�s����q��/c����WM����,c[��gF
n?����U2Me�(�M�:�z!ʲ��~{K6�љ��i�S�(�}��{��O����u9����~!f�ʙ�:4�i�vE��Rd$�$F:�d$ȑ�Ñ�l��/	F�eٕ$o�*�N�n�V�4}Rn��s�x�.�c]}&���.[�*��N����`0��1��)�e�����F���Mr\n��Э��"�>n#���'5��B0���w��g;JIàO˵��"����������{��s�8�pX��}Cסfʂ���d$U����q	�y����{W� $ {��8����<�4�Vp#E]��JX��'ź���Ɔ�Z�$�GO���9�l#$��d�|Q��m���Os3D��̶a�|���ɝ_�_[t�G�O�6g������r�;9��\�\�~]����a9�����h��H�Ә�r���u,	��հ�RR���Ƨ��}b�����/�T�؟�"*�5��KV�a���g���B���l�3(���1ޜAd�z��CkV�\B^��f5���x�^&E���y6�y-�l�,'a�S��U�v��m�A�\�?hp�t_64{����^�2���bqA`�Os|���Z ����AC ��=�O׋?����O�i�ֺ�}Vt(�R���k�T�7�H	��v��G��@�ض*�R�^��q&�-��;۹��{��^ݕ<��j����و#6�-p�����.��$�9P)���XH6���l�Um:�f#S=B�G�yb �$U�aKԭ�
�3�&���n
�#��g�������nM��]�v'
_�ְ�q:G�U�h{���a�[t��!�!��D�'��9�Lnv?;�:%�^ֺ�����"�:K��W{��yMa���m;~�	k���VN<�@�Rh 4zq97�{sR�.�)�~�(~��ʤ�ݒ�"ɢ�¿]�j��V=}�k��"+_#�	>]�hU]�!��g��>�	
�>z:^*ڐ�ͩ��O/w�Q��B�~]o�A՘�_d�P����g�JIP���@1�4��>�E���Ǉ�(Չ���4A�e��m����	���9P��	k�y����B[X�?d-Sn6��9�����|�U�fA����΍��?�my�Q��'�6�Q�F#�������n)L5+�;v�:E�u7s�	tu�b��Ĕ|�<r��J}�(�-�O��A�=۱ffC�Y�:os�%�p�q��fv���/#�ڟ��L�a�B9�,��x"~�%�5d���;��4ִA%xO��d�ހș������m:��T�Ʉ�&3��A��at;޼V��=̻m�r��������!*�n�,m41�[��ρ��pQH���$�MruƢ`p�cpt �N1{�eՓ�R}�(b@T�m�M������5/�:��Qى�w���yR�v)��s#40Y������쨬����� ����k!��`�aU.Q����[O�ӞSi�	q��=�����y����S�����N|y��5��%��}�,ٖ���ْjJ���6.J�%���K�:�[Nm�`<i��,Da`U��,�uޠ<c?��[Ԋ�����\�Jʪ=�N/�|�_%�D?���p���3ͅ���-)�e�@���������#¨fY���UglUŭ�P��'.�m���)�r������e�
3���n����M�&�mg,�xW:�xضPt���7�]V�����R:ˁ�+�4y/J�vF#�E"	�3������j&�m���;ž�l:h����Ay&��w����N�T�ŷ��{rf�8��q�"g�����|��[��_����p"b�͏Y~A�d!Xg$X���"�w��*���j����J0͞�Z:D�<�k�N?���L���r�ѝV�ʽ���H;\A}
h�D�奚�W����{��l�R��nF6����lhD?�"������#"w�15|W�BB��7,�0d�h3�e=�� ^��ZĆ�n&TtP�-�V��]����;�1�?2v�S�"t�V�~j���xK���n�-ޕ��C����[,sL�];v=-ҷ�Ŏ�v�A�gV��~��0	,��������x{>��_j9Kˇ�N<��Y��7�HY꿟������5Æ~󪚏d����ehK�bo����$�YWm?�:u�}��,N:��}G*��dI���Da0��Kg���~���������j�2�x����	.�N�YQF���B4��Ѥg?�x�z���[g�k�PoN����U��E��4�^Y�H����}Ta��N��3�"�6�5$p��i�H0:�Q�@Ո�EB^���=�>�,
&0����nc�fv�]�0�;��$�]ej/̥y�&�/ �#
��8�j
�2^NFv\#TH���ފ'���0�߸��]����o���xNx�R�y�7�=YL���0潐������g�C��>�)���/p*^�Һ.T<����X�FNX�j�3`<0��ĄE?�j��[��J	�B�ZİX�z�J�ry�/�a	�Dʹ�[�L3%�������~�e�ِ��@Wu������̫�p_Ý�oh���Q����X�rx����� ���Zr-[�o|�"��^�F��Ó!	P i��
͏��:	��w�(l�D�M �u\`|��	߳������K�.m|�{S���?���5f��a_|��(]t�u�4�E����t�y��~���&Į�T��.
��V0�����2@�+�mrx9�.��A�{4**� ���Tø5� v�ܦ��D��~XcQ����&�k��V9wv\2���-�zcI�/e��C���г�]@�Y�m��\+����Q��7��o;�6L�'���4�� ��yO�#F���,��t����g�� �EQ>(DO�sq't�����Nm�ѹϸo_���r�6c*��#8<{a>v��@/u[���7��R�p�϶�j�x�_����/�3׬���&�0'[)�f#Ea�s4d𮂁o� �� ����{��T!`������{�{s��v���q3;W7���r���#�2� ����@K��M�H5�;M�)��t9�ʠ��@�%�J�jHt�uҨ�J3��'�q+#���^�׽$5�d_q��˟�3�?���^�51Oi�%��0S�H:��v���Kg������|�[{T`�&o�(w��g:ȕ�-�9L��7 �o�e+��'�����|N��1G/�//ը/�����Q��N�w�Ձ�	H'��衉5 ԣRQ]�	4��q7�����Xy蒋��9���d�aY����^��=����o�W����O��c�no%Ƃ[�/n���"�nj�7�\kbu&��G/1o1�(ƏR�N�m����E��ޞ��Q�i�U�nk�$��PH�7t���:S�Ct��ɹ1�)�/����]g<YD�_�m�Fg5�3� �}՜���Qaᑱ@_����Ѝ��L��*� ����_X֬��gj�+��>h���"�-��M4����ܟb�.�5�'{����R�Q���xr=s0Q�B��&A�ΈM�NV�^��b�r���B���i�[��R�qap���FT2y?��i�:p~�eK�#=f,�2�]��&��*��2���ݜ�D�{��@LJl"	^Rc�$���S"��p)�"�[3�sK�0,�+��:
Hb�����hM����7=er����E���9�T�-rhk啾�V�p y�z2��#;���>���L5`N����o��y��j�o}�Ha���e�H �L�dά���v������W��o�-Teaꈋ��F�_���Z��sX�Vq
����
�-dr���	}�ݏ�Ƽ�~����fSPD�.!.�=�O�Q�����~ÿ�X"H�1 �Q�T10*��G�*������ٛ��=gғ��)� 3q��R�j�`�oIYԅ +G���BZ�N*V��4pTR*zn1��j{ ���![�w�W<J)o
�K��_b�VpSjo���>�*��u�y���?#yx;i�<�n�!-B��+<�r%'�a�:N;�)�-WJhXu��̾K�=�i$"����iE���@6ΰ�u\�Z$gƗg�܉j͹�<IZQ�W%���.��7o;�F�%�����?t\�2{Q���E;��k��M-^���$�C^
.go
�y��^]^ W�jJ5�>�����3�b͒�n�g�٠N�K�����! �D�q�q/?��i���ז�Aa2��o��[%�Tx"�� �7�G�= �l�D쥦Rt�}Y��d�J��[�;����D#���I}B���&����!�(��	�� [+���8��:'�V%���{��E�Y\a�۟�5Y��XLҍ�5M��G��z��#뵬�5ú�Dl�g@��ʆ��Iȁ;(I̟̙�nM,�	�Q�"�Qn,tYb�����`l�����)\a�9��)Q�Wu���F�d������}U��_�ɴ�w�5�`�8���]HVx2�{5�n˂�ǔ��R2�_��;�i��f��V��-pg��Z�������0������dרf��]1ߎ��$:\��/�����[94�R�ﶚ�S,�i�ᵅ'7����іGq He�rl��cȓ�
�CΪ�j$G�2�&J͘I�h�j4���DQ!�1x6g�p.%��Bj\ܸ�J`��Tq�c�'��Cw�l���e��?fC��<f��F�o$e�fH�vR �bS�YX<��r%�r��^%�ü^
�L焙��H�wq�
�nHJ�"�Iz=|��%"eG�a-ĒA��}NG4|j���F1A:���,+2&�n������cܻf=�Y=k��Y���*�@���{���J���+Fq��\w��b���!�5�q*!G@���DUgPV��#������=�ϑ���m�?
������X���b&��W�L�0.@�����},j���̴/f��h!�f����^���*�����{�o��%$p��/�lXkf��ms
FB/�;�DNO���ף.�bn�S�&��0~�rL)!G���5`Gx���>�Xq��;��ٌH��<���Ct\7'�;fPE�Ⱥ��^K��e�|+�PQz��p���&#GJ���ax�-gv�T'w������)_��B�m�3n��7]4F�U�~��S�f`wg{hN�:�b)���z�b�C�R��MC���H�E���&>>��q�Z��CB��K�S�H9��à�0�UN��QC�_�uHe���`��:�5�m�����J8�E�m4�4K�w����e�#�.L��>��r�~79��N����7ԫ6͹�U^vX���̚�����ܛNy��̜4'�4���t&-�T"U�@o��yu�X@(�3?3�L��Eމ�vǝ=4i�)^�q���r+���+�ШJ^(���+`�KG]o�9g}o��A_�}���4~�J�"h�n���Iv��ytb 8��g@ �l�I��f����Hk'� �O�i:B�R�dBJ�'���"�y�f�)��t��M�jwЌ�ܭ��J��R,�O��n�-���V�������fG~G@�̒C+��G�G���8�"7������_$�{��S#So ^�TaJ�u!7H�6�b�x�kl�/n~�1Yl��*�i�.��q�,�X�so������߫�b�t,�9E��UӢ���[��z�F^4G�AS-OS�%�+L�׺k�f����~hM���Ffu�e٫Ob�
�������/-�������a���t���d���אʻ��I�}鱋����%�}���ߝ�x.[��1hQ��[[B0?X�D8����w��`#����v��b���D ��j����^1��	�����C�N��σ�>V�@��Г���'k<o��ŭ�2:uYz��H��D����c	'ok�މZ|5ۖÑDMQ�鿸�s����R���ͦ|��v0T��ۆ�e���>�7?��g)(��:�f���px���(e��ᴦ�>�fX��K:���UҮ"ߗ��X�fF<&\G�Z��~׹�/�G��T�-n(dJo�/�ͱ́#���!���ъm�Y���M�Hnk��	|Ao��e�mM>�	�=�&��5���7�^�t�e:K�!L��MVu!9YǤ��rqp�0�I`����mS�>]���(ȶ���.:0����s$�(�yF��
�K�Z;��4�JZΨ��{��<�N�	��$B��%N�Ĕo���&E�Zǹ�&)��u�SST�)�q��ـ���b�*\Zm��%�e~'�*��b���q��������$�%Eb��	�)�X9�Uo-7���A0�6ڕ'�Zs��iU(�o8t����At35�i�=?�~�����=J�5v��t�~E}x�P���m
ȑ�M:������"���!T���?�mO��Q��{�a��9�(��2m�@�PQ��Q���ge��9��]�C��dI����^�y�t�(6d��B"�}�7�R-�n^���.�XRz�tѶR�>Q�P�\��J$�z$�\�U�FJ����;�f����{�(F�{+�B<�w�H���c|,J��H8�E+�K������r��|���Ki���C�Ci��x��f~`���N��:���G���x��}2K]y��8k�&aǽz����~+�e��dC�"ʬ��Z/���.��p��x�W��)�(��[���7~zw����<h�8��*�3�EX�s����&טN_�qh�:�߂�I|ٿ�"�W�TF�%/�搤��?H��##�8�z֣4uOg��)�Q�M�'��a�iuD�t]Ҿ$]ob��r�%����? ��c�s���P9H���+����[L���R~���.�p{� X'� ��
�U��`��U�%b�GYo -����Pkf���@��S�W�|��%J&>ǐDżWU<��`��LE��>�g��/��A(���M����R��6kY��@���-��V�_Zk\}�?0�|��6+����q�@�}�4K.����"a<�6O��������fN��7��.6�EB`� ��LU��	����(b圫��Ҥ��)R�"�[��Ú�yx?�Y�K'_����F�!4����(�t�WV.�[2�B(�K�O%*�X�ϠrK`�]^F=2yv&һ7i-�{\Tx��۰��ll��VJ_ww��<�[�Q��덻�b�3��P���T�ͼ�%�-����6OE'��R���A�*����k�c �>��S� ���R(R�'�#;�߉��0�#Dw6��e�'j����GB�����`i���'k�?�f���O���U��a���%�����S��E�]�
��۲��7Q�{/�B�i9������I��wF[�=d���+9�}H�Q�ahN��� �h�$��7����~c���$�$�����[���BȖ���<l5�Dސ�Giz�y�'�j�����n��Ⱥȿ'�+�域Р���E��W2�ݘ��,9��&�5�KMjOegW2�h0�|5s�gB���LP�`��:�1�}hh�{'G~sV���X��X��UIJV�b����*�B�!��!��7��n�[�J�{Ix��b:��w��R[��N�-��/�E�'y]*Z,�&3$MJ�EBh7 �c/����;�wC0�DMG��}����7ڷ�C3�����F�G�X�dX��[�3'S��{������P0Ó�ҫ�������d��O�3�Q�:w�W�D�s)�w؈���ZInK��d��1n���'3RI�4p_�[DC��JŇ2�3֍9�'Ip�<���Y���Մ�d������B�}��»Ȑ{��t��Ov*�sP�c�s_E�=�1p�,R�����s�b���.�4�-o�$������u���rm�A�R�c�p"�)�*`L^�L�p������wk��C���{�̒�����5JFz��BP	Ӹs��-���	��t
����L	L���	[�eo�g`��X�&�;H2c�J��cק���g�v��Pسv��V�8�a��k7���)VE�]l����/��I�&��o
 ����( �/��Z�D8#��s)	�X��wc�EV3 �BO��hr�y��V_��EU��#���Y���z�&����s���F�NȮ��Ǳ�L�s~Ab�Cb���4�����&���q�jL��hN��u�/zbjĸ!������J��.R��^a��z�Y��\�*8�D�5ȶ}J�d�����|s�C2/=o��)IL7o$�ޥ�H�QMy.0O��J���L�f�)�/�z��T9-�Љ�����O�X�ͺ`�6�q`�u{��FJ®[s3���c}^T��\�WX2ʬZ3�GE��~����z>�j�����Psȑ���3)\`�a����Ǎj�2�+����p7cML��Fu�%y���Ʊ�#��A7�i���A�\&XQ�1�cz �������D�e���1$�69��M��&"�jc��܏���'Mg�JU+Wm�u����z�\G������nMd�'_���w���z��`y呁t�Ī�����r�(���3�i"�3}���D\�2��<}5v07:{ռ�5.�H�����y�X)��L��D��8�(���қb�t��y�E�[&2Jr�V�@+ t��!��:�G�Kh�(<�rBI��6f�����D6������E��+������YW���6��cu�yqy����xJ� ���QUUמ���n��F�f�Ĕ$d�J�ޖ�	ݞ�/�g��%j$��;@r<�w�}�@���3|�CeW ^/&P+��@By,?2�ϯ�3s�5Ep��_�5d�~��x)6=?	��"F�$nӫ�5XQ�`��7)(ݟ'�UX$�-!mq��)OvG�
�z����/@̊��O-�Ǉ#�a�2����.*��I��*k2_n��2��O�I̔ �-m�h��Ռ��6�$�NT[�O>Ȍ7���5ϟt����Q0�,���\I��)DNXs���9<�!��Y Ƕ���&�F���j�i��3^�nѯ�s�)�מۂ1��¬�1��^fsl� ~�C½g%;VE���y�䗟5����f6�A9Mҭ�e�[�����׏o4�c�a:Q&#��`Bi+����:���o_0[wd[27���%{/�}��*����S��3Qs	8���Ӳd�,v6�Y T��@Y��
H=��>��o�?�&8�Og�J��F�»�ы� 9�]JSv��L�z�3�����h�u'�[�G�Ӿ�7.l���@D���q�:�����T�L�'�+`>NB|�@���p[���Fo�.�����-�^�m�;O1	e�`16��,Ce�շ=�����#@��#j21�vwV
_�G{�ke�2���W� �>0<��Ш\<��� 0�qy�-I~����m��x0��u���c�XK��@��0� �F�y���8��\��-�^r³�	,�1�o*�!H�����v�W��*��by]� ���|����B��O��V�j3�Ns���
��#A��>�13������=�W��!���*~�􏺻Tٛ�1�b?H��������8��#�]��vE��kM�2\6]�A�����OK��1p�~��;��b^j\�M�=ѕ�vz�n��K*��),�{�Q�L~�E2�{=�_�� M8c!z��C�
�� lu�dH��soH���T�NB�gin���3'��_�nH{Z� ��{��������vW8��8�P(���$��5AHr���{m� ]�pD��w�?��%íg�We%�AF$=��BOTWm���AH�x��+B,�#�檈-9�!"���}C�'�ӽTAS��t?\X��E��Q��	��Υ=wDd	�B��z��{ӖGŭ?s2����Ջ�ŋ?.dy&�g�iAi������ɰ;z2\6�C�M�U�lP����nkK�p����}���lh�a�4�7�H���3�_񮃓4�bVM��V�pef�)T��h��a�AI�B�7ar?('$̞��PD�mA|�n/br����N�y�2��ĝbU
X��Z�F����g�6@�YӞz�XO�Ƀu%�DZ��}��ʇ��7��17�W�o;<����[n}Z29"���^�\�2��\k�|��9Y �����zo����򥯽������;a�u� r��i���"ɧ#��v�3Z���b�zW� K��� ��'�{��}����ٳ0���'d_���/�Ѽ�c��A�!����۫�ތo/�$��ƛ�}�V�1J������[Iհ�h7J�G'��e�j,}WW��C���$]���#�&E_u'u�<顝1�hO �\�r����Wr4��[.x'�?�� ��7�"��}ߍ�`�V���\j�n������.Ov�C� ��Ů�#%��|�g�K���~��1!�uf��o�Y���K��ٌ�ݧ�=�p�f��[3�2Os�[�n���-q1�����G�6�L���\.C�Uj�L�:���(��K��U�=m]�X�~����\B�a\l%
(I$ˣ��yA���ݑ<��Spp��5�b��0ܪ`�8ȯy����В*F�D���.�ҽgWv��k���I]�o���kk%Ek4�{��A���6��ۃg8\��u�V����m�q��@���(��26`"�g6�0��(�!j��r���I����@�?��y��4�=��&�#wscA�S-��Y֋���=%6�r��x��#9�<#�'�\&�7�{��G�Ԟ�V�$JBpT\ēT��gvѓ
�~ٍQO�R*�@�_�b��-��Y<,w_�.)�b�d�lq�(ٖs���P̵�i���/��|�Ja*%�����56>����<}��$:�{�	�Σ�>��?Y^Ab�.���~՗{�с��wb)��;o6kyj����]c_r#���+����A�g�Abo���vz\+{R���"Q�芨�$���_A��2ϩ@w�6�.4�@��@��ڮN�|�y"mҀ4Q���>o�n��g~��k=v>yb���_��$4�_y���Z$�n���d=��v���%�p�]h���κ�qX��P�hٮB���!Ʌ#�5
fV�ks��<!���I�(�x8��o7C��5 ���Gx�j�G ��m������~E���6����b�Lx�@ D׉H��ѷ�F�i���yg?��Q��Ҥt���̡x�T���.yߟi��ע�������o��4GR����Ժ�=��Յ|"�S��W�nF��1'�s�l<7������#J	gUF&X�3�Y���GY���m�8�bNM����%��70;رg��ɡv�2##��e�U[�ƽp�Tz?~�iϻ�I��׼���
yv�d#��~�e���6w����W1����07i+�
��r�zħ�_��d�N+�NgWR�[�QE�jۘX����Q���O�OVy����[�n���0����6�T�h�v�4s��z����уm�o(�%j�ro���蕡W�#���H�� /Bg ��T� ,�iv���]��p�[l�5��f�s^Cꗆ�%8*0��ۆ�r�!�<[�S�>l�˻;��+_qd��M ���n�d
���H�Ko:mbu�Q � �$5%�Κ�˧'JR�ݫ8�O1��5\��,#�pp�
a!�*�_��b��zs\���9:�%��N��&q?�U����e��%��I���Z�B���cM��U�fVH
{c�}�$4�7�ώ�}L��u����Ik�V�����k	���g�==��CX[f�:&C�t��}~�4�hݘ�~f\
2Ğ���.�<�n6�?W��1A�X�����ʄ�|_UmJ�F}r�4�[2��5�����*�f����'Ƞr ��u���+u��M�w���F�Jx��]�B�qi���/�r``v���3�ˏN,^&l���pؙA`�ݑ)�~o���š|fG[e�-��|��.���^D����V�/ʎ�z5��B�EV�}�䛩�?E��ë�湍Lw��ϫ�i�e�e��F�_�f�2�o�[`N��{���
J�ܥ�S���O�6zjd�څq��'U? �����06�N����a3�Q� X5¤�)���y�'�����5b[pNv���a6��1Ʀ���Ƙ��v������8�[&�.�6.���	M���m$ș�ч�Z���+����O������)� �3ήP��f&T��i�R�ʤA��g0C�;g&�j�~��z�گԵ��r�.hk9�eb�ڶ�'/�>C�2���+P�f�.)?q�^��5��ҭ�_Ek�0���\�5@�	��1�?��+
�>r���~�;$��>���������(��{V�ȑ�,�Kz?�,DF��Z�OSTfZ+Zp�Ev�]�eP�N�^��\w�$!k�(v�(����� B0���5|�X_ܕZo��Ӌx9�䃰/�m.��Xu�n����AN���Q���~ly��r� �����ٮ��¢��`���8��Xugc;�!^��%��'2D32e�J��P��Oƨ�&��@;���ň`^Y���'6l',�Fg�	3����B��1���ɿ �!$�{Z�����kdz"�Hʀ��H'�3��	Q�L[+c_w�-�h���!"`-��aD�E�y�����]�D���[/�ݮ��<A���0Lm�I#e�.&�.tX��'����ț�.˾�vAjQ>���-�o�o^�l����I�����B"`���/�~�౑h	���G��B���5'I@o�?��7�D����ً��0=D����K8Y��c��
�i�{:>x�����������ڛ=W�' �$r�U>��OL��d�L�( }7�=a��뤀(�]N�?\\:��&�v�ߘ0 �J��t~���΋^$+M	T���l���dPղ�j���i;38ݩü��F>!�7�eHI�z�|E󞫕~�\�>G�t��}�=|���.���t7�zs�M0Ր���I�v�ΰ�5��0��#;�%Ў&�Q97����l����X*h��--��l� �?t�� �%%]�{�.�>��wd*����#���t!J�|xЦoe��q�-��D��aO��4/��}����0��O���w�;�F%7�t��C�-���䎚�3+��Lb��$��$�ݍD���*�ֳ't��o8gg�-K7A&(b;���[zֽ�Њ��Lwy\��h���;�0R2�bbW�庌���m���6`��MeY���>�ۍJ�����t�</}$�A`YRn~�:���t�/!a�c��I�sq�������*�.��:c�Zs�p���N��(��nOs�W:Փ�̓���*	#h�kFAU��^����%V*������}\�1_�*�	]�׫-q(%�2��&����\FnE����(�����NSN]�2�ܵs��6�E���C!�;��[���}ڻ|hI�
L?-ƵX�h��p���B�ק��7���_Ā�Q�g���n��l��X&�m�	����߱��h�f�sM�ͼD-ؒ���kg��%�*n�τ��Ql,e�C�r��ɮ�w�qK�e�<j��@�����gM,W����O����}�P~�L����U�ފ��D".k���n����;��lI�Tz�]Y8"$F��D�	�R������x��1�i�J3\?4TPC&⭎f�-#�af4�Gmv��{�1q)+�!�>$pĀO"���_X�A���5~c�M�+�|�Ƶ'1���I������@&8i��v�+mnL���木��q�+���4�hc�����L���썶��R�W@�b-���4��V����п2����]�Cc����d�g���|c�(Xxp��#0H�Z(aψKk��~�[�vo��XV�b�㉔��S�~,�݃��T��Ҡdx�T�_�v�Le~]�ʟG�~��� 6�G_�p4�5D;�n�L$5+��G~q�UDX�-�9OeF�
Cjq����&���pQ�Y2�=�U1(��fm����q��ZmHA�*]l����Z���~�x��@��. 'T9H\�a����~򛚫~�~­�G�W������i��A�
8
�)H�5��5~�B�y�㜞���%�3���\ӀW�q��K����
�3 +Xt�&FUm,@�qyޓ�A��gV�v�&���,W�@��ފ���ݸ���l�Jh���l b�Ak7��/(8�9���ʭ�Ď���{�W�����Ç�Q\�(����֫���PQZ�>L���<~�3�A�QH�̇�����c�"mUP7�� z4+(��K��(T��R���<K@
,Qax��c� w���	�m�=�z�.�˥Nu"��ԿD��`B�"��`e2c5���ԺD���4�t�
�0��Cg4G.9cb?������Ǔ+Y�;x^I+�?���;�pYa���Y�=ԙ���=�Ys�k��q���+rZ4^��Ȭm��s��<��s|j0�*f4_�<���>���2��wL�y���4�л7�&�6z24��r���-�M��k�q�ڿ�'"��d�=N�d?�.��2H�w|Ёo'gl��0l=�OP�]����GA��(���n�)Nm%MV ѽ@V��J�(�;,#�P7���{�[�ҩ��ϵ��I���f|�Gz���K_���9K���T��}�e(K�X�^od9����j���_�_�C..+�^���iw|��!���)e�����V��6|�3= �}X�`�7�|��.�ct���(��}7j�lY,�ڤ�8���U�p�t&RM�*�&��˝8�iA�l��RCZVuj����Hs�>|n+ӘV`58�a�6�L��ds��� �t��	�����ן�\&_/����F{#\��H#�������1�E 싒�R�9?��(�&7�<@'�p
:n�(�['��}��	�ʢ���z�H)���� ���w�I���5ga�Va�4�"	�=�ՀT�?T�Gȷ�O�tiF`c��r#���(���1=�-9m���;�F�o2�Tӽ2�U`�H���E�sz�f� �Wp]8���;K��/��z�<ώWjc���L1^w&D&�d�$;��) �|G_��a�qL���S�-�<c�et�U�a�I�`���#a���E~� �K��gW_m�r��m4-��b9Ң������C�Ĺ�7.�ᢆ�z
L��B.���S� �vP��"��8�D�=�m'��'p�]���<����YrRZ}����O O�6��ca���L�Yw�N&v�0vHu�r��ݵ�]q��8��=_��e���D@ ub�U�e���1w���m�����x����F,8�����qk{Q����_Ģem�O��֓93�d;��I���&ƛ���������R~6� ����*}���g�J$�u̔��zZ�6~�t�g����;�t�J������ ��%�2�GS�6,f �?^v�\jTd-������	��	����+� twЬM:��aHa+4��t�(�*�_
ũ0��U�E�L�y�����ş��.v��M�FZ����;��iahF�Ѥ
6�3���3w�tˬU�n�)�O�yS?"�	���Mh�l���T-�a�y�u�
{bN���<Ω�� ����B���1�z�_>�b-�bc�.>̋^LE{�B�=��t�&��V-�y�!��26_���= ��FJ���E7�E�]<���(�]*O1iP�X��Ex�)x�"�IAg����Jt�\)5��X�'��Bʰa�?`���N����w�:#�����bQ�,�w�&+:�)��D�&��?^�N�����
�fPV��<!V���g<�$�n�T:��*�K$.?Rq�ܛY�Z�
z��UP����DQB\=Qv�VG?�l�>�� ����k�����բk$��k�t��^/f;i�QS���G�>~Ȣ�3�_$�wb!}���z����x#��e�҅���eC!ʼ��5��R �	T���}��7�������
ӥ��ԉ�+|��ΖaD��H�=m�qX\ʦvg�w��q0.��<��&V98�4{ $vF��,�����`��K�3�*�ʷ���E811A|�x6Ӕ�^����M#!B�;_$W��N�'�s��,Qz!.:/���C�K���w��.w�1S	���߆Ol<�J.�%��#��eT=&�z��OnPF?�&�2���紾�'�<`�K�ܺ�t63\�A\�;zڕ�\�n�(�������~��f�?/��*}Oy�a��sF�/��-�˒ud>뽹����~
ȩ��!����%���n9N(y��A&��E���˜�U����&@�ua����d0�&L�xM���S�<q�������{A�kti�{��|��s�_v-�r?��M8{}.� _Kr������[5B]�L])v��A/`�i��'ri"YD侕����j)��۹�^+dT���J�Ӑ�i̤a��GԚ������|#��[��yS�K��FFu����7����O��u���K�ź"1��ږmk��J�,�V�E������t4�n�_'@����a���O� �ed��%��|�a�/N"��i�sU��㺟�&��T��۫�C�o�(=�V��ڥ��ˬ!%X]�G��k5-�oe�Q�Ж�ԍ�����L��
�%o�j�۔_�9���e�.�grNv��m�o�Z#~:D�.���x٬�F���٘O�{*��]�5W�V2��e�K�+E^��Qл�n4ʪ	�vf_d-��S��4k�C�"0x)����\��&KHw}<�E��L�v��ᄱTbwQ�����P�mU�*��!� АK5�^1(hU�upkd�ͺ����~��,��������+	���D��$&�@�C�
����L���p@҈� \�/����~5���4�[���sm�G�����\W�z�S�װ�g��ݒ�����IhT�u��E�O4۷k�T(�Ӂ����g��+���^����<ଇ��ƽв�W�Ze)���/
Գ)�a�׮��3�{
��Q`�'�}��;駘�ʹ�;�Q|vM� t�]��
��m27�+ԯ���oF���C��t_=%���+�h���e��!�	��S���d��|'����pU"�0�Pf���PIcH�b��3���@wv��?�ބێې���		J���z_�gw����y�,k�I]�_��f���Z.���$OG�ɤs�7U�
�0E��
��9@��)��&N2Or?�̓���i�n�B%�0^�p�U�&^���f,�Ɓi���r���\����B.4`��ڍICO/��/��9��ݤq>Uܑ��"T"��EM�ýq]�����@E*����^cu��}h��ڇ�"��e0c�Q��������#�B:(�th�~nk*�~�׳�f=���4S��]�I�b�y��\�í�j<�8Sы(t��K�8�Dj%B�'/��d|�+3)H8��	?5.>KG�	�e֍����۬B'�?��9&1%����ȰZ�fغ����^"b�`��#�k6���c��r��3�x�m�_,V�ǈ����}gG����� ���
Z��A����s�~:�*�������؁?�q�Y����* T|�W!h���c�T�n&���d&���)��"D����V��x���
��m���d�D��{f*�^��k7�݃�)��߇��V��@�vE?�H��s�Sli'�Ja8Z1?Χ )��X��l�˞���a�¾J|k[@t v9e�pı��+�����Q�:@��*�Jf��^l���G׍9o�����I���c��UPLL� /�:D�����2	N�E�,е�i*����d�9��ݺ/��m��ؽd��6xuw���[$T�Y����N-���U-Q_�1ĵ����یN�m�pmeN7d����� 鷚�	����0A�_��wz�8ٹ��<���Q��W)�Db�Ů���Y��-_�i� ����q7�Z|�^X484�9t,	%�S�|E���Z=ΐ9e�IC�ᶹ`���/OMQz��Ã��z�3y!�-�[[���t#���A��0��AH|s��	��Q+��`��z��D<�iLE'�e�1 �)!�oo*��Q��9��4%��-Z�]M�~�Kǉ�S�:��A��>L˺$
�c�$��'��E)�+�����F	�_���iGRh���@k1e1ȑ�M�Bp ���.��� �$�|�r�c=��'
��F���V��P1��������h���]9��v|^����葯�߃$d0���g2K�x\���O2���%T ١e�V��nu �8��)��~���`����鹒��
�H�js#rrWB8����)�����M9�#��E�R��wz�ݣ�+��)|b�@V�������
�t�8��E{cNx��IU�e]�cD�h���خ��R�,�&��w��m���@�K���d�qj��V�?�nj
�Frψ���_x����1�1<J�{�/�����i݄�y�x[�f"a�c۷�bv����Y�D�$͝��������Tb�+4�#dW�U\����M���W^�ҥ7�sAjV��J_�?C��/�.�}�/�o���^�$���nW�Ml�@Ѱ��;�E��Q����B�4�}ԅ�ܗp� ��nn�81��O��N/��W������^#��Z����  \p&ɣԑ^B���|���Ft�<�2�Ҡ9ʊ_�����JFͬG�a'���Iɀ���qV��R�er��9\k��&��I�����F<s���?gD�)~~��R-���Jv.dXP'���)�E/O<�NB�p0Q�R��%�h��dF�p����;Q3��2���)Q#ҫ�|����K��X�����V�Ǝ=�N���o����5'��ˣ&v9{������[�0�m
vv֌�7δ���9������;���~ZV��A�uni��8)�8�غW���E�d�ڬY���]&ɝ������M=�}�s��s�4MHAp��鉫K���G��L��Q���	\wӉ�/�xن^��ƾ"*2�F/�r�`pW��tc���Sx�`��6Y���#R����p�=Ġ�Z@#"3���M�8���c�s��V81�yv���ߔ3����sN����smn�[69Y)�?��*u�������,T���Rg��śa��vz=��*�����A WA���.F���X#�����7C�kZ74�E֤��2�M����@!�gM�]2��x�{#t���|����}��i9�
�.�^�0�z@eЉ~5�v�Ά��7�X�j�#�@.Ab��^�}�cP��@9���&�'b^?����:u� �w��bx�Ō�.�(J�����l�����)�E4Ռr���+bՕ��օzά"�2���EU�7�w���E�3˿r�źmeD;�uxI7��k�O��H>Ū��X|� <�	�>����&.���� �����]�-�܌�4�J���҆�%`��ܣeU�i���s�A�_�3+9�$(��8��ؾM�+\O8?v!�%�����e
M~R����/*�B��Fz�|��a13�l���y���k���J��s�>nu�6}e3���U.,��ｯ&�X���M�3RT��A�������`g�5�1�m�q��/�r���kC��&|��nAL���|��1`�❔������\�ܘ���\���bs��,�ZH�
Yz�l�����!W���8r�
�u�wwg��&&�?Ȉ�B
~6Ոe��%+�T/^��4�e�J��k��:��H �0�Bv���G1+�o.�z��ڱ���5�`�(�
6�1*�S&M����yO����F�<$��Kv�w�u(�6H��|O5A_0�긋\H�w�1��\�*$ �＞c���%��^���u8`9�A�9DG��,������98����{d��������6������}Z:��Kڐ���Ŷ
�N����J�G3&�"�pq =�b0;]aT�������8�."�z�+mz,ݱO?m�5�e����ns_�n~q����C׊(|�4d��B'�����;<�;*	����]@�|�U��&rqt(�����W��~R�V'�#<�����#��#����@/ФL��w�{��Xk�#�ؗ( e߭�����&S^�QlqzaC�f_��ա��j�c+h݋4��3 hgZm����v� ��M��̀������P=����ni�������Fk���5���!SlP�h�A=X4�j�<މ��@�%*�3�t��_���
=Æ`��:txU�A�9��=UK�g�� �-�=�bi �[�
�~喘�����<�=���9��N�rCDi���
�`o�l��Y���T�7�v���wJ @����ַ<0A��I���;�%1c�t���Q���ޕKR����#��.e�)�S!�Q���,B�a��m��X�t�����>�4C�c$L�O$�}+p��$�4��G��\1������W��Ț�Ũ���~J+j��Vh���De0N�o� g��qE`�n#/��(ъ�l�Y�Y5��[�&)��!Xh3�]�}U74'Cd%�xDG/y͒�H.f������s+�Y��f�(�p�� ����EW�g��4��ͦe��w��f�!|����@�}a��Q8As�S���][[��p�@���lh��aKzz�p�v�r���uG��F��o�a"񰱂|�����i�U\s>Sy�G���nZ�n�7y��Z.�p�%�SE���rP�I�}{P��sYt@j�]�
D����`L��Q$e?C�G)�;��qj�g�Ԉ2��]�U�\�裕��N�<(1�l�}��CW��zДM��p �ٰ۷5�g��.��wA�6re��ѣȏ�A���1��g/���J��?��C�BG�A u*��eeh*y�����B	!H���s���퇘\�RR�� �#"y��;*��z?m��]��=#o`�Нd��J�2������~�h7�/�HE�˭&��:�"��x:�� K#^]�#-t3"�� ��/��G�g�aq�չbc�ʠ��6� �
�
+P��P����s1� s{���ݍ��..���������p�ҘS��u��^'1��S�X]��q���(cvB���.�QV̟4R��0�s>��������d�Ï�6S�7퉽:sƁ����p��C�Chf�l�aX�Tf�k6lS"[������*�u�x槁��ϊu��i\�4Y��'���Se��!�!�rκ�,��z���<�0c��yk�cJ52j6�%-��qb����h�Ӫ�F��Tϟ�e��晳���bkӨ�B���Dy�!R�k�R��)�q��ԊAb!�M`���eE�m��5'+!�y�+�Ka�ϯ�߱���J�>�����BY�q�_q���Tera��Rg��8��86]7���cx<��F�w �x�y1�R} ��g>	�X�U3.9bݹ�� �{o�A��7n.��� ���z�m�� ¨�!���������U��T�ޤ)����{���ɲ4�)� ���6SL�|c
lp��,G8c^�]�;h�_�<\/�<?ZY��[�c��I3���GW�"���{�a-7�a��CĚ#�@t�K���^'���〇F��n�����V��/tg)�Ō��ၗ!ˈ/��Ĉ#���ݩV4F
�qvp�>�L���®Ea�F΀y(&%�wJ�u��]�qה�N��-Gn'�(���;h�S�/Ϋ�bi�CF�g�h7�6����������=���E����D�<^�]-�|���q�
�=�!��C��< >뿹�v�Y��0j\���]f�=Z�
�ڥ��(�
I���KU�|zj��yz����;E�r�g�m�G�樧T [+O��(#���=�u7�|+�ۥ��d��L��)�T
R����J�5`3"�&sy-y=�a��ڭ�UC�D��
m:��Xu��o��wT�?���g�,�u�h�+]��6.@��:w��x]>ϔ\�~���Yeb�"�f�r��j�p�uغ���˫����+�q�tĎX���v8�vJ�3�
,^`��W���*��k|?
�.2��k6�YtaZl�;�U��}V���j��j��!g�>6�S
z?f[���b�a���'ߘv��Fty���H~�"u��D�i1_[/���Β�V�"`Q�SZn�#��> ]�g� �n�ic�=����&�W�`؈���d5��2��k��J�$l}�p6�SF��I.@-�oJ�mW��B#��Q(>7g�����i��� �2���	�b��5!J;�	�u���S�f���եAa�W���6���D>*2=�o�>2W,���'c7(�l����E��c��G;�����f䂞����H������<��U�qeY�G�	xwd�u�{]����Ͻ����'G#�p�����C���ԡ��f?��(��Ǉ��.:r$l���p ���U�����յWÄ 
�,��î ]ͪɥ�ţ��B"f*��Fp ��A C�x@���Y g6.�]
9�_���w.����Px�h�AD���/�"�6��#�c�IvtI�i��OMˋ�����E��c��cb��k��E�L�}]+�q�{_�T��(���w�D��Iắ�oݺJ�ߺWE �E�.�Q�Tu�h�#�S%��V��A^���@��X}�Ã/j��at�T�j�@/g�or�j�y�W~����&� ���U�kn���h1�GtZ)y�k���*�en$wvF��DĀ��
�e3[�$���R_s�=��6U�Yx*LD�����~ԏ��\&�0j����mxq�s���%�������<��<ۦ���G��Q}ZP��:Z�tyJz����F&�:i.7�ft)I��yGԅ���A�����!�"�X����`�cs��y�WA`؅	��d�e�$�'��	~�2B�/tXu;�-���s)���� ��)w)���"�ZNl�t,�ӖG���La���G��V���mؐ�;i��� 7�����y�E�kT��V��vZ�k�\u*7O瓳�HП��.�(kA�����	��ǽx�C�,����L�V�\�D�-w���=��znn,�,��P�Lo��o�U��s�FMer�?~�?�ƥQ:+����ç;���ʑ�"�.�"�-����|���ƣ�1GZ/�)e
2. C�� ��C^�v*�!���v#��lz�ه)z�|���<.X$Q,��F	�1S��r��|p�dP��2���]���:a8>#ɐ�⧾�R�y�m-�D��B�Vֆ�(|s����؉��ʽ�V�mrt���a�+1U-(�����(T�������!e��#�:Q�{H^���٩��-[���4��P�a�/X���إ���w�^y�|��ϡ���H{��d>�W*��8����{�ea���	��4;��<m��<�������-6�U+�80��3�U��2�%��;���!߾���]S6ꘀ���bԎV-�s��ch���"�Chdf� Cm��7�3!�ݐ�}f4{O�( �6��	m�F��;�;��ɹʝ�NTs�8V�"J��#�/Ȳ�ܤ��?����h"'|]V��n�һ1}-(I�3Ε�@#y�*�#\��7�u�qb`����=a����Q>��
&f{oI5�ZL"�=�h?��C�S�C�YB?b����F���U��j�`�1����)�d�9��I"tю�3�z҆�m"����s�k��yRX����8�@��]��T.\�I<�|.�N�8!)�u��e�r۠{���+%F.�.���-w�Vq+t�.c3;ۘ�P��O3J��%��d�|	p��Q���=j�ٶ���|;�$V�l&�}xm���0�Hr�c���,��� `h^�G�Q!����� �tk Tc�VU0ى��A��׬�#2nl���<Q�g����l�=�ISfyq��*x�����^\m��>�#�5���l���ќ��Uc@U(��qK<z�F��f�������-��dT��UB�ϔH����R���>Z���J����#})���x̵���P~��"4��2Z��%�t�#��y&��[0���H��u�=B:=n�9�~���@F9|R�b�Ro��c�"�#�$���[:�M��l�o�"�mJmCvJI��3>΃�S(����m(�����xL=<��:w���6t<����u�����x��țM��ʕu�->[�]"BL��p��An��}��o�)K���nJW6{k"�Qk',�)焾DW�Z��'EW=��r��8o9#N�8��b�!
��f��Mް@����Ί_%���o�>�m8"�)��D������b{h���Rh��W��[0�YB�����S�e1�Ѣŷ�d&���
���!?X���s�¾��B5���b�4�|M[M�'���;N`J2]��/��:���%p�g;A�-�U�-���_�d����K�D��p��>]�d�%�f4袚�,)#m��
�\��4��?���Z6X�)�FthmrF��mӐp;�w�o�LAu�����|���I:�����	���H�OY��E�V��2����c|�y�%���8��q��l �G����/�.�R�=��f��������	��IC��T	ȑXmO?B ��UZ�����N���I"đ���+3�ݮ��[�Zd6�0�M��~��e����6��k*�'��Mu��0�k{sڝ%4)"	n�|�Ͷ}��i)y�M�&���R[z��k��@u��D��#@|�7��g�iUDhcj^uKHR�>A_�cn�Q�"P^���x�z�dw;=�F�\���Xߝ㕶��-ȩ
���h~%ӥ�$M;��qf��ݹ�-�ٰQ�q�6₲ŧ2��0���pGXc[9��D�ۧcV"��R�1��{�鴪nɺ���uE��<�O댘�jn�����,+����d���y�uurS�fI�LM���O�P�u5Y�~Kd3'���	�~��&彐i_���6�ZN���LA��#A�R.XQK�
��n��
r���G�9(�D���s��~�l���Y#?k�wB���	��:Im|n�8��".�6�i����l��ʑ���ә{��G��p�m�2�N�39�5�U�ǩ6^�7��G,8������ a����jv�Ԇ�Ӱl��v5��#kt���"kF���6U
Ywp��[�^7�-���Ϝt���K��fj�Von���Yki�^��v�rMd���Q�4(P7��hDz�X�u�j��Kz��3&��$��ZS��_яIJ���9�Άl� SF$*Qb�Zܘf���)�#��ڳ���L�&R�=9������a��]����� ƮNS鈎��ɩ� ���I�dO�GA$����EK�����m;����U�]����2�-z!���9��o:2WjU�LՆ���K�P�ݺ/q)mGf���ZZ�~̎����AB���2���ŭ�8+%�]�J2�)�,�oϗ�;�<Q�}��b�6�r�5q���Up�k�������,_8oQӬ]r��Ok	0�E~Ó�O;LTKt��7�p� �(�O^����u��i�;�wg��r��:����3Ǫ�lz�OO`�ʡ�/�T_�
��l-*�4ݥ�)�x�P���0qSbB,�����ȇ��G��ض�0\!���� Z %L�  �pD~;b�DQ�rØ���n���^�4�����Ư��Q����V�`��{�0=�N���`ȳ�5wϰ���l7�2/3�%F?q�C
_i�ە����j|A2�o�} �pDrV���H��Ү�S]p�
�����L���Ͷ3�?a���(z^̢A荵iЅ�h,��U�'�h���H�i����j{־�K�Y�+]��X����{�'������2Y�	ڍt"c㜅�<�i^��!E�]W-��M��5V���<��ߐ��g,(K9���s(0���y���Bk���@�;e���x�{�����6�0׌����yU��P-+�)|�#��C�K\�JG��#���l�𘹎�咵���H�]���qR���"��|!�6'=�$���sv�Zځd��1O�:�BݦD	p��~k�|£����j���������.d(���3�6ߠڭ���~vHJ�Ǩt/a� 3� �A�TK������K�{p�kX����0}� vC�1��&~~�����B���Eñ�k��Q�v]�B�$w|�#b�Ib`��!��gA�tỊ�#Ҥ�I�K,x��K}��h.�p� �k�)��J؃W;g�y�0���M������G�q�Mw�,B�"=e[p����S�2k��2;�l|�������c=*O�)���:+�f*Z�w��������S�Q�k|���Ɓ7����C��r��
�buY��x��E*�f�1鯎�	_4Z����gcy���0��aT�ؠ ��ګ13����!G�A�}��,#��8$�;�ؕvx�\Ŭ�!`��B��Z��]�؄�S�-��<�[��$o�����Nq��g���Il�Ċ�2�9 L���d���y��l�h$qL,@��E������:��߮�IW��ب��^z�=��`�ќ�i�5z�Q��oWW�:H�[#:h��}�W-0�:v	P�OB���1M��Kuh5����9�!��E��q���k�,�KQI+�	��B/G��ҁ4O�]޼G��v�F�,_#c���sqٯ����ڭ�PJ������o6����R_./Ƕ)h YN3����m��tGR�����Ǖ����/�!!C2d.G�g�`�T���r4�pgK��J��)�8y�Qq����@�����d�+�4�I�2ʭ`�^�oI�Ae��ׁ�q��Wy.;�:]<K1 ��-�1��J���=!j���]4��z�� 
�܃�I	�����֮�B�I��{�c�Oc�+����-���+]q�ڜ*'�����4�K:�s�c���Q�� dWH��1Ϳ�g'~¼JٳeX��Q�z���0a�3΀e��sC+2��d�<K�M'f���k� 0a��eСH��O<dj	X��8Y��CL#���gb�0�����I���ܰ:�҃���y~�v�T� �Xݜ�O�.�z�D�� �a��H#U����u���n����`�ʥ���P1ì+=p�J�*4�
_&�Ÿ���^�Qr	`����2Lp�/K��EI��>���Ů�I�A���\��OO3X���Xe���2��r/"Z�̖w���M���$�zN��!�D/n5�TR�G'��.�&�U}1�&F�/8�RU�
��՚X�P�(5(��Jslw��cin�N�Im.�a|[�d���1SPWge��r�ʧ����~Li�	�Ù��hL��s%���xr�<12c���4�g/H}�4��O��t�#��Sߤ����6G� �w��m���2Vy���6Ҋ���b&ΫA��FV����8�҂�v�U��*w�I�<��T�[J>�6b/��5NA��8��X���Y�"b[�k/�,T1įb�D�`aZDG�V�ZW�t���y�Tsj�q���2Q�D�^�a���4�3N?��?Q�}���o?�q(�������a�kݕ�r��n�홊��u�E=[��t��n��ںV��4���T���R�SJ/�7�!,NxE�%��.��%��7�rT�?ۖ'��K[	t����=AiE��x&֚	���#z"�^s/�Rb�ݚ����k�M�wj�H	��ஂ�d]�#ݦ�p6S��+,֒�8,�W��g�m�Z��w��C���V��X�*�I��a�$vEO���ʒ'i4#��W,�[��L�^?5h���_������L�kDy���g7�Ԉ��k� P:K.B��5�t��Ռ$�C2�Ujj3	o����v̵��(xM'��geHz��&Ox�Ip����:p?���1q�zK�
Za���j	5|NN٢	M94 �vFG�����iĖ;�� \C�ۖ����K/�Z�����0�gzy��#������r� ����x����:��m�9���&��W`�m�馣k���B˄%�H����dQ`( ���c��V��U=�<� ^B!�ԚiC�l)�ʹN	��8���$"�7 �{��ȧ]e(hw�å ���(B"�z� ��G(�ڐ:A�T��O{U^?�D,��鹳T��|�T{������O@���G��шz���Ȳ���K�]�g	TC���L����VDG�����V���,�lڢ�8�NB����L�s����TTNZ���a�G���Q�|Ea
p�Hy�E9�f0b�@������PXך��~�.���"��[;5j,���4�';��Z�l�iY��LRz-w-��R��B57?v3�>"����B5�W��*GKOUk9�xK 7�L��&���Ǹ���a}��oue�pv0O�Zɧ>hϝ�XE��ٓ���i�>�̰�x�I����`@��6���ָiJ����B�ר��/e�r<K��i�u�]��a�^	�ې�\�U�|Z���`���an�F-`�۽�c9�
�>9RA_�ȤO��Bl�&{y]��Zf�_pZ�
�)��r��m.�ĈA�����m�|����E��=����=��P5C�h�g�h,�wq �?z� ��S9��v�R��ǒ����A��+��">F��^G��Xm�^�{z�7�Y�W��vo5������rSZ搘Z��FBx��̙��ݽ8`�%��m�k��BP��[�ۚYuj�_�u�T����`9Ҥ;�?�[��H��{����%�b]����Q���5�<����"�<� UC��Zj�gn����J��'�h����������^��Vp0s��KI@8�}-/k4���2�Mg��7�@��uБ���4u���<����_�l�F�y�QAF���t��� G��G"Pi�_M��6�^�K��)��x���Ӄ.��:s�τ�Nx?^���Ygh�9�� z�k�G,����6�ߪ��VO-[���2=xU9����_�� �����V��w� ��Cd����`b��&�]f�����kZC��-�fD}�n�;|s����QDS�5��"�.`�O��,R9�§�������~?��Abdܘ�o�� ,6��q��*c�D+U�O9Ulc���r�I�&�p��ԇsZ���b�c][,��
[0��T�[A��ȿ���g��&���L��n�pq��C��3�	��r� �ꅀ0�/I�+^��`N�Zw��i9k�m��#��y!"(��0͂/Gw�N �M*3�˅lP�M <*���Ԛc�.;�T��.0��0=IHl�S���Z<7�I8���%�K�K���� $����r����Nh��p�(�h�ߕ眔���H��dR<������}�N=^ֳ���u�M)�2�d1�szJ���x��iv�U0�n���}:�r,Q��iE�U7	+4�4�?��|�"�k���w�.2���߹h<���8+�}tm���x5�-Hy� �6���^�ሑ(�����;�N���St�T����^~�w�>��� ���O�5���17*��ˉDZ��A�E�Xx�J����P�|0!���q*�C*)A�9K��@O��m� @��G�ןP�OԱ��gҐc}j�eᄃ�t�h�7?����Z*藤���p�Uӡ��'`�;b�����3�:n�s
{s�B4�	��;B�����>��g�~��߷w�(�Y������q	]G��o7cȏ܊���o �lT���߂������p�+1�[��͝S��u�C���\qE�}�pe�tMD���G��:�)sG�.�E����CO4X����������T��~�k>6\I�ԉ޶W�����잮ML�"&ޟϽ93�v�����}qS���"���Gu��ߡ��l }l+��</��~8�Q)���_��/����m���4�8.^��"DF�c瓟�!L�m�W^`H"wX�3�K��	f��A�}��{Ldڎ�;�;�;'�y�bȆ��n2���p��>�O��-/��JRT���&7]/�����BF*>��^Zc� ^z�/���W��9]=쓊��xf'h��FP��<�1�ւ&��V��<�dᤞ���V�ZCx!{h��Q��[���5�iw�`�29��$s)d�������5˺�Tc�^�B�����;���{�&�o�h`�8�I,��$�~��I%ڿ
�X�FyC5���f�;� ��ƈ�h��Dܼ!�*���5966@8�8����}�Q	���*>�*2�.�!�[�/�*x����n:H���<��:y5�1�_i<_�<IV��S]�S��U�v�Ec��i��#�@�@6(��̆)�(��~�e���`���S)j�����y�;f�=��k�	rU@��{��k��m�����(oQ�döM�!h�sf�S�Be�H6Px�Dm�NayD���(�Rs���;s{�^THϖ��*�}_�*�9���E�k�y�ZL ����F�
B�A%������>4g����?
vU� n�e�i�3'
��`h⹢�<XR	"�f7.Ą�U���ٛ
�g�� ��7Zm4����7J1k�� P��.��u`L��`$�A�bϩ�cz����*_��U<�b���Hu�W�H��ɥ7r`�^/w,'���W�UC����N�P����zS��\��h����a�U�۷%4tk�QE4�[�־�AW����RG���P�7tf�D��>b�)��<�c�4��]yˈ�8���Rf絶���0�꒷*�����䵫Vϧ�C����Ђ )H�!R�yW��o��I������܆է�ׇ{�/�r���7�ϣ}r������<�خ���.���͋2ksܔ���CV���@r�]��9ew�<MĈ��b��)qMRBA�Hg ;Xs��c�Jn�s���n��*:����I��D7]��k�{$_?>L��`����/G��<�4�x%뭓�*�R�4�Xh`ӥǔZ3t�~#K-�HA#�T�9�G}==h���Yɮ��xr�xև(���f�,Q`$^�Qo����ؾp@f���q��7����	l��;;��'K��~]�%7n(�ֲJ>.An��>����Q���GJ����`��M�ݟ��!6L�1�T-��a�	"��٨���U���yv#��X�|��i�C4�L?2�ME% ��	�Raa��F[ {����W�P34��<8�$[����[�jC�;%T�,^>�'e �ԁc�V����p�>�`e6="��>OY