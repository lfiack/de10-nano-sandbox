��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG�V������ܴV�������`��m<��1��M�Io�|��`�#{w]��7�^�����D�����)�VY,E��*Ǳ��C�L(5�`����N�����W��h�2_�(�::w���{��4L�����z1��#ڪ,׫"m�M3b�[�[+����e,y=q����M�K��&w�9�=�l����z���m7�S@�??�+�����~�R5{�2����P���e�K�73��;�f`���-)ޣ;����)Hj�̅]��p��bO�O���q����QL�ا�R���u����~6�8Υ�<Ue�>���l1d�(�c/�<�QP*����c5dI�}�rb�z��gI��#
�}��*��p4���	��9��9%mǇ��=�r��+�LY�Ve�(I<��QqUヰLA�0G*Py���zNGzgp�*�R���;J��9`��"����T]��	_�)�uv�Y��KQmM��	�,�H�*<^�@yt��\"\��x~B�
�%�^L��������SK�:��6ӴP��\�c��	���V.L�2�S�w.^
�5Z�XP�u������n���d2=��A�Z(�N$1PC��}�:�Y���W���h��K��N[��k����Aǭ1um1�D�R��^}�?z��4�;�R���vcr��lZhP�3	y{Z�&��Y�%s�V�Ck���Qr&����R�GhL��8��337���J�Q|v|LQ�>�� �[� rd���<T�={���ˠ���<�����?Ӗ��d��/#�4>��o�JĎR"�d�Nh�x��}J4��H��q�D���	u���AJ��J�,���wL�* ���/��v��1��]��3�Ƽ�X��;�xIZ���>�d@pf�N�d��0I��2!��=�{eވ�3Γ����P�@46���T��<<��+*w;�sLq�i�Q�ơs8���󄋯e�soN䮔��)q�)8;�e�FV�ז}J��X���vQ���ᛈ����&�����t�ն1�aR�2M�PU��0/����=��ϪMK��^�]8�r���|K)p�}R�v���Jq3�W{!.�~�R&q'H�f���	o�{�$������q��^�׋L���.���_�ލx���lƑ>sL�L$?8	��4��_��2=ۭnR$Ѕ�����$v��������?(�!*��۲�8�{��8͎&qʕL�)���������e��A��_M��Z&��:=�mh��xJ�v��ؤ��Z�f����v�)��S����B��
ބ%buZ3�����B���n�f���mѼ�S�, �52���<���c;�֙��q���o�������EH���^l#J@x��S��KkP��Db��Qjm��J��R������G����{U_P2��:����N' KZ,3O�U��<|���&��s/F
Ϗ�䆣�6�@q��"��sJ{ɀ����N�Ð�V�|=�#���^��ϸ�w^K���h8:ȇ�`�I畍͹���έ�̌�o��t�+�
2#�z���>�2V9?�[�Q���ڍ������Nx�/bb<��w%W�Н����w>���W�)yB����ޕ����#�?a�x��j����Q�Q�g��cW>���������=�
>��Ǻ3��
�D��9/�
"t���k� �X:~������|�!��K��y����N�h�vJa���n��8ik)����)���Mf�94V�n�C\�eR~B���q���Us�$��@s��S(W3qr�L�-�g{��'��ɳ���9��螞Q�8`:�x�XS��sUJ��R�#�c|A�z�H$��P��3����W-�S	r{ۉ)��R4F�^�'s�3Ⱥ�0��mt���ds�U�nC+@��q+����h:oíR������5 �\]V`9Ik��
��7i�Z�6�\�im��]��8��\443��_-���^��I�;����Pn�^�� �&6bO158;zNt��?Z��X����݅5Œ�0�\�I�%!}A4�NT	k}���%��oV�x��&�H��Qw�=	��Ķ����ȜE�覹���XH~:@k�1��k3��?��'���y(��j_	����;���a8���u#�f���0,3K,�g2R���S�����^:i%��\��̽�$��b���Z*�r�:/����p���$rA؁K���'6E�b����._�ގ���l�6��cH��2�L(:���?�3��̀�6j7��K5L"Ȣ�gפ���w�^����	6����Kw��m�e����B�(0�=��k?��� i�a����*��kw.�~��kt{òI�5�n��WAK���N�$V�LT(wQ����%�TՈv�<�vp&�8l}ص��g��