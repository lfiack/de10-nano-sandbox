
module nios0_ip (
	clk_clk,
	reset_reset_n,
	leds_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	leds_export;
endmodule
