��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG��_ �9FL�����h=B���|��s�O<���/_2�� ��h��S����xr3���]i�_��2���13Qӫ�2|W����]Ł��p�q�H��4J��p��;������2ȱ`�|ߖ�4�$c����f���f���G�a�����\�(Ҙ's�q�й�	�	T+p���Ö�2$4���9��IUN����s[6Au��)ڥ~i �,4a\󺺈 �ytfţY�Rb����1����l���ڡ���y
�%��N�2��.��~	&� HO�L�i����8�F1U=��qF�:P]`�6�c	вwy����3�O>�,��/E�^�j�c� �n���׶�㘉�������x^p<��4���
u_載��/0\�bw����+xy�pK0.��@L7�$��G9�2�ʕ=��Aôgt����\i�Af=�a=>9�����&|Q�D�p� 
xho���6����fQ�&r[��S3|�g��f��/����L�[x7� n�R�0����O�<��x%���K���펵��A�K4�R���dK���M�a���N�T�$�̾��}��A��ڝPn���mB��ލ<ES��fI�VV<�(c�$3. /U����qh�)�Z��zN�)���o��S&�6p#*�xMS�9k�rh?����?鿠D��䥤��4�aо�X�� d~�	��x�h�@H5nJ7p�}�H\����w�WF��I[l�΃�a��-;R؂Wf�'���Cb�1v���_�|y[B�=�@�]V���DĖ�v�N��O��^/|�/���
��_6�RK��Z �@5�yi4@S�(WI����LSg5����OS#���R���Dr�UqC���M*.�x���W��J�	�	�Q�=�Q2�7��x:�����	��h@�9c*U�T*����Q�Èm�kf镀�4�}�*X'��l{A~���P:�ѨYݨ|5t�k�r������~,��/_��y�"���{%�к^V�����Ж�{�؃�d0�rE,��'`�O���>׈���}�cF�z���eo������^_rW����V2`�$l$$ ���2�Q��n�������/�]h+�s�H�sů�F2�.]�����4�jM}��Sv�~C�muX���rm��H�ܡ����Q�g����;4�T�d�D�rR750%�Mi)x��+��#��/�p�13�%���֟#���"�%F��wW}� /�^�j��}�6� /?�@���%�>(XJtQ�t� �r62�[����w�aYh��_4�$��j�Td�	�������R����:��Y7����(�.�b�G�N �]�I���SUj�daz�g��Λdgs��Wګ��P���u@��\�3�]��J�o�R��e��-j�� rzK�T�~��b�N��	D���5L�qy��L�F$@�n-����cOU�zb��o %�u�[�
�9u��j"x�;O���R�m�GW���}Ul�+s�p���Zn�K1�s��hyP�r�e2כ}����Y�b�m���L��Ot�wf�#E��i�n���ء����as>���j��:�諔
�
M|�w�_�q�_�VE��g�*�O=A�w��q/�U^Yy�::��R��f��Ezn��8�$i'2p�1���}���R���~=�q5H�����^M�:`��U
�����I�]b4��:�.u^�}�ۭ|�[l}y!Jv�se?s'\hx����Z�J�e�����#b͊zA�� F�0(��wfa���f�Y�h�Q�#�Sy�r9<\��,	�
	�=Φ4�ԱVy�[���˒i�*��+�������fߪ9W�r���,��z�L��=G9c���P��d@�m��|��B�<���QYBH������c�C���;��s�f������]�'K<|l�n!��A�[:ixt�d���0>���5�{>c.e�|D��H�='�)rd����-{l�O��%�}1�к�s������+�fh:�/`a����2E�0r�{q�f�)��hއ�W}����:}U�^=���''a.�	cP ��]��CC	��ԥ���w��i��.�����[臒�c�1(T㗌�=�䄽:�$��~2F��ѫ;m�ΗF\*q�O��|���/.�"�����3�J(;\��KJ)Lp�w��L^�ҹ_�#�R��K:%arg�-^yl��_�4� z����j�S�}?�#�����{�3���@�_�P"�;����E���H�O,[
P�[�!W�[���]�,G��{^����>쵐�LP�3h�MO���bjI� �u<��{1գ{ھ�xv>�$���Z�I��F��í$�*�D�-`�\�`&��-
��w�tk�Y�+�.-�bl ;x��`	A,��^�H�{�jL�H�#=L,��!���<O��DZ3&����V��]L;��!�-�)x�\9?t�'������߄Zx="�n|��6[g�#����NR��T�?p{Sp6Ǔ3C�?�RM`z� /Z�K���~�t5E�'��S�E~M�bbPP�"
m��lt�SU�2�a^����!8����%mѯ�e�IY������)��"Aӯ���y ��$���T��f�t}It��3ƚN���bu��:����[j���^��-]k���_���:/�u1��@��O���j�aIt\s92�ƍz'�)ڗ���lֽ]{#(�z�6%/�U���إp�����EwM)�}���r��蠔P�΋�K�O�ԙ�H�x1��A-�5������#��>�-V��zVK�6@��I�S
V+[�	qi�r�<�cU�0�s�AL(j�y�ek�����=�x�b>>g���/�TMd�dk��(S�8bի�<�6q�&� �XT&Y��D"��k����o݉�l�M���i��!���}���̀��
Ǭ��gذ�ߜ�
��߅D�	h��Ԅ{����D�x�Y|�s>K!���7��L���������ٖtN Ѿ�����0��>���l�"Ĩ�g�L(bd�u��~#Ψ{i� ��<z:0  N�Pi����Ӯ��e�_�ͤ$��o�V+������I{��&�b���kӈVc=G��K&�AP0��te����5Ȓ�~�S$U���:HOR�=� �2�ٞ��e����]��x�T.��g���b�J��?W���`֖1�+���F����� Bb��;��j�p��e,�Fѧإ�i����Ӷ?T��tTtO��X�.�.�%&ۥ���� ���	���dK�p��&�s
}���e���͹���f�"�E���,ET�_�����}��U��R�ȺiC�T�DC踧��^���_��Y7��j��)$��e�R�W+���)�k��F�)���@��ĩ��~�4hlϧ�x�x6�\Y���nO���?��5C}���ۗ�n�l�>�V˷�l�);-݆�"�N͸d�(�,�.���-�X�?!M�RX!�|�7q�pQ3=��BR��d٠���p7<����G�O����G���H�60}�ޭ��u��
e�e��ҼUmJ"�zЖ���:�;�l���.�DC��Q�65��?2zrs]�@��y	9� ?�G��[�IՕi��HKz%��hwd�&��r�^J��?k����p���7༫Z�V�[ƽ'�0�5��V���{�>�{�F�،�E;�f��A�eL�����$�-�*~�^H��k8[���$W˿����6�"1�"z��_�D"��?��}F"��,����=����+c��x��&���������b�� ��'�%�?��ˣ'�E��w7e(���
�D02�������?d��өݵO�RbM<5j����cՐ�k��v�J�zc�bd�R�AY Tp��=~�S� ���F$w�����4��<J�8t�����9�݈�k�,�t7��p�ɟ�-5�mA}�ԍ\0l������N���c7$[eiFQhX8�?ɵ��Gŏ* ���o�0�h�����Xd�8gu����,bm��j�#Ϙ@��x�;��W�2��ؐ��L�˞jJm�j9x�P��>ͨS�w��ǒ��Z�D��b7��}"�8�i�!_�j���@�'Pzj��/
���S�F��"6�r���|����`?_p�l�O���������9^�2Ǯ@<i7��ް�is�_\q/��db�$XLޏC)C�ܫ��WőrE�%g ��tK����0�[��_L��I Ƒf���(Ȕ��7��o�vPbbf��(��)��o��Ѷ��Q)�k��l�����)�o#�LL�9��F�{�d�1x0YK�� -��Q+�g���Da�>.�	�,B ����8a��,�z���
�L��r֦J�{���(����:�p��8b������]T1X�(v��;ʦ�8@�cȯ+��Qr@���8M��ҋx,�躳�cr#t������Le����g���u�v�$0,����R�ٙ)n�Im�����sS���#c��ͤ:�_=9�3p:�y
q�%녅nA����f��ֆ�@1��0�T��i�^�@�6��Ȏ����4l�����p:n��2%��2�m����>��f��@g��<�!ϊ37 1|���	�*�[��Ң��yoU��{��?�F�>�U6= �{�¢'i��^r����m�j�k�D={Jh�U�L�0ƁޮnZ�s7�z�<���ߎ5tJ��n~�C��<�������|w�~���?��޼	��%bL<=U1(+�>�&�jrvDM�?��u��	!)�%#H�A.L�������2��4��m��/�?iG�/����1��`�&�Le���%IK�}�$'�%��j�}�W4�,��Y.�'�+��L&�1�2n84`̲�$))I�^ z�츊��7=D�T>�)��f
PIΣ��5 �9���� !W����a�.��!�%��c�q���Y($�l`J��w
�g��@8+U��}��9$��f���S������̓�B������O��x�~�7"�F ������]J�f��Ea��*q�
���b��O]P������B(�:'�Z��-r	�D?TS�(���JzgK���mS�!��E<{=DW�/�=>���E&$�T�픋h�a�sU�w�]s�B)�>=�������}�1�l �����^�Ux���K��>W���4�;l��猒`�=���_��?L:p��_@_�1n������
�>2(C�Lǂ|��.������l�̈q��7�X0�#�|��=A��µ!���������t���
X�mYQ(ϲ�����<�p.�Y�O����T-yT�~%)�ː�~�'�ޥ�%��a�N�O���CIE�6�j7ՆV�(�..�O�bk%J�#�|l��)��X���j��X��@y<�� ��ax��SÖ���m��5��P�a8�n��Ґ���khȦL��[���ykV�b���x�h�DnOm�'L�Zp3ć뇞���qfJ�M��O*r+�H,>�ݸB����b�7��&T
�E�{�� <��e��{%����>�pɵ��1�jg��ya���D@ y��}� #��KD��6�bGpD\!����R