��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�A 晶�}Sn%�yS��O�VO}�����;��G��Y��#ݓ�Cp�n��m�*� k�7�S��t ���`K�j�E���W��(*�o�ql�b�n$�%���J�S���_L�Ï'VG]�7���$�4S��I,������_]�z4�U�/~tC�l��aI���u�|�6i|��mor�N=�O��'�3t║]�3[��bOFG��M�f/$(���ͅ ^
p�gy���Hv!�6�7�ᇼ���~H,ɳ�U-�v�0��c=�e���7CP��H<�����S�I,�/Q�@�aO��3��2;H4b0k\��7i+8x~��ۢnEwlћ+���,eK�NM[MM�h����yk��5�4��q0��HqPT28g��2#�9dj���?�į
>�m���i�(,e=i��EV��L��|g�T�^�`
�6D��G�#�W\(1��Mέt5�Vaɨ�cH��W>�#�N����yh�r������瘃8C[.e�#I�LI��aD,�#sQ�͑�̗�<N*8	�N���&�7����ts����V�I�^��kK��#u�z��DӠ���(�Ҵ�G�7��ZLDi\���)WG�2m�����DH�NƲo]��[�˃\P�
�\�H���P���A8�lK|2��|�N/m��p�XۥnP���x#�4)�"����s��tn��q�p%w4k���,��-_�������wb��$�ĕ5{�
'��V��C4 ����<_tQ2;2e�����n�D�#����s��d)�ص{�U�N��c-#�O���{K}�}U�Z��od{>8h@������'�Gf�A����"ig$�����+��҆�t^��E���z��{�h����5{��0s�A�ڰ���97�)�b҃1*/D7T F\ED��!����_�j����q˟ �|���"��- �",�Ó�#�N��Mט=�~yeg�ē����X�0����O$.ڭ`C�c\�11J�'�6���������9Bֳ���*S��/ �	b��B=R�*=��� (L��u�G^\�5���&l�u� �f�B����?����#��fz�u�(�$���Sh&�4��!#���F"���=X;y@
o�ᇨ��,J�;�r�K-B��d�Z���������^B���vS�XIkkyf��r���F-v�Pt9�@W��C�GMy������Z�p�]p�y�k&� �\h<�3!��ե�Z��y��|M��R:�rX���e)�9I(��;qr)�f^J�wY_��u��6Fέ��[��9�����VyT	̠�r�D�>X��iUI�z�+ߠ�t-��W%7�3�ZH��$B�=ڵ���n�g�Cu��@���M�D���X��G���קZ���V�3��h!JjK%d\��8@r�k΃q���XE<��t��|���(LM���ϒ�J��@��rmu}d�%��<��mb]��>ċ3�ɱS�V�g��%�n��%�.pp�X������~���-�M��{��R���n"%%��S�f�wV�56��Ͼ���.M_��]c���-NlDR�d��q��(y͆�yFk�q0'�<$S�Ұlk�jM���z��w��s�8ΌgV��P�~���a�>-X;�r��B���0��FVN�t֚�T���$0Gt��E-�>�1d꿴b�a�C:�dFLN�s�7&��o�ᱩ�	 ��U�[�;�1�x�u�{"P�G��z�ԇ|��`\�2����cŗB`���&0��:GB|�'��$�����9������/���{�B�Q,�%cdh�VS��;���I,��8�{�b�d2�`���2��XO���^�T�bM2�dH:)	�1zݲ��1h����`у蠧����N뺢A3�$=��}��%����SF̰K�`���U���!3�廀P�����H������ބ`l�]q���i��vy��/	�-^���)��šɅGaS����9�$qm�]Q׵��Fn�!�ܢ)ٻ� 3�
�6	~�!�c��?���i�C�ٕ1Q�?�[���E�
)B�U�����g�~㥉,�����M�����뙛�hɷ"���yY��R�ϢGRsK�"+�,��qJ�R�5�Q���븛�m0��?�$<em��c�ht��m�p�˗��C��Tff�n���E��}v*q���+�P�T�Oqe�=��ԇ��x跾Bv������䗜u�����r�4�6�t�$�NJs��i+;���J�n� 6������E�x���d	`��� �����`ԑ@������uXtv�S+��������/��`�֔ZD�s����j� at]�C�]�V,H�a����L���{��+=�]��@.�#�R
'�~�M��#��:r��$Q���)�}W���0�Zp�	0�Ɔ!���y[���$�<�$�ۃ��E(��_�S2��6/�iRAȾڀi+��>nJ�oG5j{�\�]*'�b�?36���FY�\��M"J�%�[яw�sкu���]*׌fD^����o���p{ٻأ�$�_���������63�v���Bd�S�B����=�Đ�_�F3�_٣9Dٹ�=�X��:!�������̛$�;���h���{�U�7l}Oq�Ե��1�V�2�6:PJr���h���m�`���~��e���/Ho5���=�5�L�Hɦ;گ[���P�!�/0o2�5���b���?��S���癘� ��̝�G�c*E���z�Z�f�#�Ȇ+2��������&#PH�]����F�7-(�Z�����bO,@��P��2����j)3Y��/:GЊ/��@*�k��J�H�����uFŭ+��q�Z��MyV�^�T��뤒6���h}�p(�k]�a(�P������b\��Y�-���#��h���qXs�4<E:b��<̡���vJ� �".�*�3�='��9�����q;���Zp*�U�ĝfl�t���p-�@�x��7�jEpl�,�����f��$��c�"�0����Fل�Id2�kr��n� ˒%���y~dg�v�U��4��~�}�%�+g/����MJ`�����ۇ�K�k�ec:�JD&�{lp ~���;x8{E-[d6)R�Z$f6��1"�H�`����`L�
k��������趩�� N����]�k��@(�!љ:�!S�:O�4\�������`a��>ugc���d�a��
Y���4D,�B�E��q�o�lS����N��j����ΕZ���;(G9�u��*�qt�	��~g��R!@s���G���Z�`fC.�ӥ�n��͏���b�%���;�;+����M:d�G* �n��wj�뚴A�|��I�$>�fɍ�/��[���,����}/a&�ta��g�i"p�bn���P�HVzP� }��S����A�N�D�T�lqh���ǦWKf��-ok�&��Ƕ�"��? �tS�O�&���b���A۔�%�h�E�*g��a���(�Ʋ�Ŏ���n��xE�oҟ�,�%G�].�[D�c���vb��D�W^��;ȑ��p�1�3.m�S���Ue<�a�>��,�IO��'���1����I��R�A8��\�eg��E9Wk�@>P��l����?8$!�1br'7UC�S�zUb\��dd=��L��`�vg8���Ke�u"[�ӈn!��R�(��3������d�6祭7�Ap	Q'*�0�P�FNj-��7��e����Ao�7�<��M[߄W4!n'v���ؼ�YHZ/�ޥ��1�A`��q,L��&���0�fЄ$3*.���c̮�~[`�ϙ��a774ƞl|����&�4`Et�V0���e�9Q��n ���E�~�4�W����,�Y���������c��洓ܑ��ͷ��.��Gv�����$7�CKi�d6�2X#�r�>�	v��;�Z���E������\>[�ے{��d�Xin|�6�O�Ķ�6��B>ϩ�QQ�uT�wxo\zu-�Iյ��M
Q�ԏq�7quKs)V9%:9J]�Ў�[�B�;��	��ெ�F4���t��N�?!aͭ�kXݽ�
Ʋ}$�����B�A�AD{�i�(�^�7`�j���q�I��qy��H���v~m��G��'$�pR��l���)��	�<~o�oF\B!��XU��w��]���CO���*�H��EU.����L#��+=���9��C��H_Fs��*����f7DA����\Ǝ삁��� *{�82�ݛ�W��m%n��E׆J��Ւnhg�����;��� 1��}�4���5�s�l��x�m�ޏw̉VO�de���-A�!ײ��.l�:O){�bg?�^��S �����V�F��㹠ON� ���~�zPR ��e��ğ8�g����A����Nz���/�R���[!@�������m*PT`�f8�qN�hc�J�
�\��T��e.	�	eK���_	�j6���n6�;���1$����k��{v��#���NR�`��c��I��l&�X�$b�
���_x���oot��a�Wb�ɜ�	�h^���2~	,�p��p��'8'j��'Y�f�T��ߊ�5B�B��7o�����pfޏa>��,�X�Sl_�`��k��� �覵j�^�ΔG,N��XP���D<�e&������{��������h�����fs�j*N�ᕜu����. ���I1I$�~���z���<w�-u"W�i�Wt��}�8�Mcr����*���JNB� X�έ�j�:�:�'�ms(��:��[֍�ߌ�:�$7�|;��e�m�`�;'X�^7$�9����L��;��N[/�y̖����_Xt��Z+���`WR�`-����)�������5���/�O�7��AJ�5�ùd����ɤ���*�56�d�� 6b���{Xs��l�an��D	���ڲ@���T�)ၧ�{mC�Km�D`�8K
�O�n�Q~M�Й۔�]��1��D ��I$�,�����1P=�c��l��Z����z�s�lߢ5_i�l���,�����,�^"�&��6q���a� �63��|�*������ʆ�� O�L~|k�}t��`�ӈd��-�MI�`R�:C���<�e��1�o�|��c"�wPG�:�f��8���IaؽH�-��g���N�x�X��T�VБ�$���z
���2�2�+#Z�UB�snq�#H���:�� �i�B�C�	�8�������8�����U>�]�%�KQ2�l�T�t�g�3w@r��%�K�Է�I�L,��
��:�2��#G�ѥ��!��}SD�� � ���`ӳ��K*Jla�;ę�"y�e�'�j�:rK��
�S�"���}� U�kF@�2���s�������׆S��ܳ�`����
[;��G 
s;�qGQb��_&<TE��4k!��#�9m	�o����֡����BOg�[��L���v5��Oj8�N��</W���UP�sS����,�t,��p�g`Ki�U�ȗ�e�G��{������3��2.(�*W々���{�_�Q���2jA�`a�'�x�}Y1���C[�e���f��a6-��'��(��t�������St��']]xj��+:��(��t����N":�~Y%2�a��<�@� ��X��Xۄ� =���ibH�4O���Z�2���uM�O�=�\$@_�=�N��[����h��Iغ������qC�|g2Mva�*�L2�Ue�"A�lD;�֛��l�)9�T�]�,O�%�c��B1��R�0�L-9����W�_���Ux��k�P��-�qU��
�z��*_z��p�ב=D�O+�;^6�s>����6`	���ј�"����D1H�:�!�r��Ů�ڢQ�����s�/C���YLY�=?	�K_���e�O'�[�� ̎M� ��~�L����-��^������r�����LaJ�Q��=G�Q�d�a���^�M�-��-��Zٓ�l�X�Ϧ��f��J��~N����v�Z24�P��kii�x���c�@{�n�,&Z�����rS��HPq�G�_�������o���+؁��֑ޠhR�S�k��� � �.3W��n"�a`�ɰ�'NH����,��|��(�Q4�R9�/������>	�+�����&����pҚ�D,Rw�YZl��*�#{c��ehY(���x�g�/��\�A����H���g�k���/0�K-�}��+���jO1�qJ�@�Y�?��~48���2�/sJ��@۵��Z��#�x��ո���5�qX�ԅ��$���Cp4�o�&�{"߹ͻ��c���đZ����mL�>}�^s��ni[���vcz�<�P��4����>`���&ִ���_C��\le�$�ؚ�e�5������ �{��Ԫgh�q���i�Gӭ(ux�]L)5i`Q+��xH������[E/�� �Kp�t
˲�a'��,��X��]�l���"�8/n�o	�cy8�j_����!�vQ�b��o� ]m����%[Dy�X����h �]W3ږ8�RW?i�h�R������OEjT���
c1�!��̥��^3�*�(}��YJv�'l`�,���r��Oxw��Ī�0R5�َ?�3`����g���C��ip6���(�7.����=.߭!�����)^#6�$B9��`�D�E;�6�I�O�i��v-b=�N��bhd��wj�bM������Dr����ʎ����93]�a꟤ں�a���,5��Z>ޗ%a�
���Y�xTl2��2��G5B�u�Ey֢���- ߪY�e�1��8PZ�^�,K}6�[^q��j�r�-�O�߽����8��wt�E�gް0�:�#/z�y�\Ӌ�3�p�jꃛ ի�Y�b�)�l�2\��3Q�/��PY+*s�Z���P���@��ħ�W�����K�]��7�oR/x)����En�c�Vl��(F�����>čo۝�5�U�1j��bVǔ��}ò�G!� m���7���G�U����"�Z���HP��ݩ$�Lm� H�E=�xe����AG����E�&ݒމ��+=��<a(�ث�r�����O�
Ad�Ka(dZ���d�8E@e�z�P���>��p�{i�ޘ���!\�ʜm���!�c�b#Q	
�,�?MR��
��]�L��C��UL���e>�U�oH�R�7��P��G @�Rʆ�7�����@�M2�3O{.�֌⵴�<Ia��q�#WJ��4�@��j�5�4f����3nʤ嵖�}��Jx���==����}S�aa���F72�\�P�%9?k�_x1%YȜ�9ս+�oo�� �b���]�?V x._T�>r8̝_
/�X�s��������	�3��Q�l��_�'�4�`T�m�r[�k%կ3����*�]�����2&0�@�H��[���R��SѠ����X����*���B>�QF�PI���A����H1�OI���\���>x�(�5ˬ���� �qq����]�GAU�	���h�q�-躔�7|���UGցǓj�w��WU�4�MC}�9��Pؤ�ځgu:�6_�0Х1�d��܋P��^�����{¹g�M<s��17O�E���ݥ�,��5�Ƞ|+/�o
��%� ��yՔ��3�ĄX�+P�내y���H���擅��r�� �y�®��/
�ݻ~<&{Q�Z-��<�Oq:��[5��vC���P���ü�)�0)��ߍ��4Aē��K�	��3�8��T��F�= �،�c�.<P�D^�XWr���x�CX��$%�F���6�Y�tI��U�db<���*�<�(����5g�����A.������!Z��3#��)��a�G���RR�T9����a.�iW]]g�J�ղ�R���@���T��:������W��o��\��cCC؀�֎�t��E:gTܫ����l<%h~�e�Ș-:��v�e�WKm)�q ���Fx���(�"}ˏQ:��n�"��j�}.�}\����4-ܓ�p�ն��}+��B2��ςؓidE�^�̞�s��Jx�g�g7&���z�Z�|T�5i(���u��ˆɱ(O"��dX�G6  �25���c��t�@��J�m�Љ[D�����N�8H�4�h�s��W=��W�њ����[v	+��%�4^`�eW�o�>Ӭ��.����c��a,.M�^߸���DxV	1�+�n��i%�mQ'}���֝5�U�M�kB�(��&嶡��jߗ�ک?[Z��6��{{t�M�As_>��A�2k����U��0ak_����?��(��J��z�z	uL������9���{sA·Y�$��k���71�+���t�VϪ,7Ɯ,'�}�z�k̂��2���H�cM�x������i������5$%_�a~7��mv���n�c���,�-��:� T�'����聋.��f������E�������v�AD�`?l�C��=hsQ���2gQ�_㽇_�>�ɅWłe5�ծ������
I�۞Z޸��dYQ����êg�E�D,[�'�w]���%��`�a�|�s��D0��p�]͇n/9�7�J�y1�2J)"���ߺ�f�kR�l�Z<��/�]b�ؑ!�?BUNuռ���y�H�L!)~u�� m�R6C�(�W	�/�(wz�7G|C}^���p���H]V����k��T��J(-~��{�|�a_�8���H(�[/�0������E�l=�c��hbq{�.�(��G~ᘃ��%��#��y�z��*��d�s�S��D.��T>��楢��J���+�Ĉ1�m{��1b,_��[n����"T�X��l�3:���4�� |�r;�e܁�E��C�ݱ����cB���/`,�}0ZJ�Z��������$&5�?��BPp䑤6��r��*�)7�Q:��A:�v6����S�Y���#il<���{����e��8ns9�ϼ��G�3��тC!��?Ͱ�r�n�@�%���� ���I�>�"�?Fh�"q.	J�c���K�k�2� p���D|Y��+���&I'�K).;�fR0,ۚ+�H��vj\u��1mE�6ʀ���2�O>�_�J��T�?�4�䕊�?»S��<.I'*lh�ߒ�\�a̔�j�����wsk�R�wd%�0�R�h��@7!i����n�"��a���;U�\��3�~Ĥ�Jv�t���a�qԽ������^�����Ws�?������ڬj$P�+ �Q؛qA�8(�n��@V��d�m�n����T���27`zRW5���õ����h̂��3b0���������qֳ��T��ȏnb�k-ǐ�i���{9�5�v� ���Z�����s$��ҳ�CЭ��ec���B����姺2ݰ���5x���;���q��"Jƥxj�0q1Ş�eŗ�Ҿ������H�����*R��E��*�ˮ��ȤjF5���cOD	�L�q�����dN����^Ј���*�SG�*�4L
�g:��k�j����v���c��{��E��>r}ӁPR�Kq}�w]ܜ�E'�hh#�"v(�x��:6�ʂ 7{W���5��Y1��J�9�r"�ٓ��Q��Sc:A�	��Q�B� ���!0c�3h�WF�䖕�J+��[�vA��>P����g�Xg&�W/8
������~��F;�{�Sw^�w�4���@q*P�P]D��FpФ�Cu�y�_��ɐ,m/�@p��K�h�_��Qtt��P�ʖ��r|���/�Y��l<��ʹɬ5!��)x�9Z�C�����QKTr {�����?��$��eߤ���ו��cd4	#*4>�Rɭ���,��HH�m���;T8i��]���u<�W���[_��g�3���t������.�^�H�:��5C2X���!��C��֣Da?��7�j{��Q���	��*���N�YÊ���'?���P���ʹ%J;I �S����)��lᕐ%y%D�	�����~��Y�Hۼ�/��"U��1dz,aL%.'��M�G�)E�(�!��,z�o��:�g�R��~�W�Q�_���s�^�F��Uު��R���w���X�C�I��L�����/��~�U�u�e�Hi��^��QɴyZ��Å�-߰`�hQ�Ӽ��#]��Mt������Pq+���xh�&6ng��[��:ŀU���>
X�p�Ĭ���'��a���V�'���;�$��~yE�	�;�y��Z�0��~=R_:`�{�pC�=����B݅��D��M�>��P?�^^W8j�mQ���L$��Ylce\R����&̚#��,��01���9Z�=g�aO^V{�=��F���ֿ�,P��i�{�S�X�g<揜:Bl����CҾO��y�G�zLa��P��Y��P��7rP�����uC-��E����D�zd�$
Fz �B�~xi���M�Ϲ��G�V'(c��:������STW&딉@����蕒D��b�a�s3�ٖ���$�F�����$ר���6;��ݟUL�꥽�6VP����$��V|�3�̠�)�n�K�KN���f���`�Zv��w�R=�l8��B��,���N��{�H���M�L�M|,o�Ŷ���*�Υ �o_x�v�~X�q@�<�r82yIrSٵ�{���m�KqԒ���ݭ	駯�KqNňh�.���=�X��B��,\�Wj8%H�����.�y�[e����3E@~7�j�&tHB�0���kt�)����:�l���`%��VZ�t>��	��VMk�n�����Ss�Y���w�@:�T#���������`��8L���=�*g�W��3���|$��t&T_��Ӽ��v���O:I9`����F{��(�|B��)Z�ү��͋��0�Sզ�jd2�6T'�G���{�;G�d�u�����P���aö|��ϷԮHi�5rpO��������g��ԇ>�N$�?N��b�_���+�6���Q:w�	��]z7|�@2gy><i�KO���� �;Ao}Bo����'w��b/����D}G-�BΨY��a�?44�P����c�0Ħ]�n� p(8���8�/N%������ߐG�츫:��x{�ZI`�i�%�e	��N�'�B�%I@S�)/h�)c�&�͚�	�E��z3� �m��@��5J�U���n�.���>u�2;�j�1���}ZY@}w5lӯ��#f�o��@�4��$����zƉj�C�CQ�m:n0��l���3&W�1*t�Tض���±�V�7{� ��LZ��wo	�� a�d�|7��ԉ��1Y�<4�z�*/_���7�:5��)Ѡ��� �`.��?�'��`�#��=�$Gl]��l�W���KQF��k��G�g���[|�gM/�&�B��dh�����H�G��-i�0�aB��Y	L3wKIb1ʟ�ۆ`��9fO�%c�Y��O=��j�DY��t��}}�(��B}�qn?��wU�_�B����ż�BwѰ�E��	B�t�괖D$x��]V�$�3�!�5���p��bk���W��R�k��8���mƍ1_�+$"�c�s�����Y	�Z�ؗ$��
�\�	m�5Q��$u
"�E�[��0Lk~��2��T x*n�:�8}�͓
�؎Rt���gY��x;��}�����(W?ԟ�gaU���~�U�x��������<x$"v����rk~�j�ʁ4\Ej�Ú)2M��-�Q���qJ3�M� �� ���(e�%��?y�
h�}�BY�[*�zn�3�"zY.����������UZE���A9�M��Q��"j�7�U����O G57Q��W�"���E4|��.�G�{L��hDܶ��He�H>� ݰ�_�A�3�va6��^��b� �6$�~�/-��SU��r�[�3n�39�y%�B�lB�Փ{\6�	�Kny�*�a���_Շ��kAc��mӡ	�&t�g��No�XjX�ʊ�l~X���)�z��^���fc��k�5��kHz}C���D�����ع�k��s��k=�'%�I�k�AM�����ޠ*
�Ց���!���x	6���g�Wr���n�!Dz��G}=IWOƹ�$�U�R���x9�,1����?��T�v���EӜ�A�̂J%���ӊgĘ���Ծ���.�k�܅��x���T�y��UKĬ�9�3�d���ޭK�S������\�)����HH/x3�@���[�N��� K
�� ba��\�:Ț��r�@�^��Go�n�G��ɥX�;"�t��%��X�=�¶3r`J�E�M�P�� $��g�J��VJ[B޵��F��d#&M�]�c_�Hů�� M��
�>)�Rpr����;�~����3�B�D�<�!�,iT�k=�gI������qw��T�U?�V�)���1��'�æ�[o�O ��`�2z��U�b�Ԝ,%M*1�x�i�#j���v��1��-gڸtDq�c{�����:�}�(��h@��  s�o�۟�}��t�==2�����M˖U<�b����:ܙ}�����;�B&+��O�l/��N
���;~��C��ق��m�HW �'%�I{�ל��oZ{���X\3�I	F������rEf{W�p��?c�!.
�_b��ݟ���8���}&`�YFRhHCդJ�<B�.ŀ�(��% I����x~QyS��C�Fo!a��i8�'�m�"��"�p���R�j鯐.�#�@Z��U �+3�4�vT��n������a�m���9�����q΋�T#��%���1�`�@
�5�}�	��1��q@��6�H�+���d���v�_�΃�������qMތ�z��J�J�#������R������-pp\��r(�o,���]�Jq�nCC�p�?Н!��A&�Q���I�s�T�>��;*�R�c�}�n������bH���~�����ě$�-��b.>B:��C�
f��*j�������'��|�����*Pm�� ���մ �H<&u�Pv�^&Ke��P�Ƞ$?dJ;���?�hf��K�/s�ƸNih׀�7��L���ka���3_K����Nq#c)|�Y]�Oi��,'y�@`3wj)�{_�LA� �J�:�"���y�8X?�pn]R����"��q��z跴"���ؿ��PQ�������7ݓ�)$��wW�*�"���@�d�"��?��;-X:2mS\?� =����I�7���>R-'3u!���8m5^��Q�{����^_�T���2"���r�Q�����W��&{(�#e��	�	