��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E��,�׮ـ�-�(,��FQ�MX)8��jY��:��,n!�H��k�Mo������3��9�p2��B�vo��S��E�4��6Gc��'�Sp���kv�ù�����f��p~X�Ź���V��ru�����6�p��>����TC��䨰��v<5&�c'��zYJ/�(�Y�s�X0H�[�s����}o����Wz��/�H�j�Z�|`קw�f$hә�|�o��,��Њ�v�Bǒ���J���=ba�">��3O5��k�(;��e"(2u~��dl	J΄�1+����O7]��ɑ�GI?�1D��	��~^�[ԓ↦}~�5����_�FG����=��C߼����2
''Y8���aƌ�*jt�P���5YB���b9~8�I�b����%�4��Gb��wt�W(�a���X�dwhǦXL�i;R#�O�<Q9SdU�e����zcvk�X&)��cƸm���Į�k���6���#}��0��L8S��H���1y1HU�q�����*�������,��{��kWW��g�$b��bB=-RR_��m����'hwuϕ��e���7��f���c�X_SYT���B���{�f�|�};���bN��3菩�q����o��/h�a�<�-�Da�l��h�� �#k"��\s"��V^���}�}�v'�U�`/|]-�($���`V����v~��Xݍ>d �^x��ƶ���"�cǐÓ5��?J�;Ts�V�O���V���������s ����)�l��S��MN�(x���6|��	�BU�aN�OӔe�v3�n��QT{��z-rW"�_r�M��:�z@0���ˀ�6���t�:��o�]i��*蹯���r�n�� ���wgǄ�p�¤S��Y�9�"r��(��XC4o�N��4��C �8Z�vuS�K6�ݍm��Hcqu�a�Ǵ�-*�n_���tH��C��!��>{��f�Pz?�X���\9�X������s@��j���&Q7��WNƥ8�|_kH���R¹��F�U{K�W��O�7.���,. P{E�$�d]@�I������w�:(��������/��a�-�}�Uؼ���k��~`�����;tv�V	����s�#Q!����3�‹�w��5 ��o�yYP����P�|xSh7�1�jn0y����
,�I���M&�;Tw\���bĒ��g�-l�Ո��@�����Ug����m�6jDr#e��3�� Q����������?t6���,�fA-,�ɋk�Gի]Es�J�bw`K~ǖH4���2��^)#�����i2&b6�8Yq�����UQ��@?�<�[%��7ݪ��#�Hʪ��d�����+)=U�:��zcm�<=p�6%�±�5�G������iy���z��h1�̙cvĭad}�����C�"��4��,.��l���-���jc���=J�8�ŵw;3^����ۆ-_8w�!ɱ�~�/����9s�qP����i�b��1�渤R=�n�2�%���=|:���f��$<p=&�Q1o������qT��G�Yn�aN�W�'Z�8z�0�����4�TJp�O*�Tnϩ�3�
�9�a�^����$��'�����D9��iJp���i�����}x�<} �d�����|�9Fʼ�2��}�椪zx���$]�Ik+_�S/*�={ �	�o�)��=���|@�$	��;4�ǭP��Y�?A��;!���zKД����r�'#�\#x���n�՘�i��ID���;"B�);�t�C�p��pXl��fZ�N>=�\t��w-���w?���xB[CxZd\���qT=�G�ʸ2^����E8�i��t��l�ژz��xrVxt�<�"K�o����Q �l例�^�M��{�jcG��9#���w}h0ō�= �tV4����m���[�)I�j��R�t�Q��`'Ʃ�o�/6��ۺj0�3�"n���%%�z�m-r��@�[�x���c�o!��=O�����ٛ�$�Ǌmk��*���Q��rJ�V��#iٗ��\��������U�޾nQ��[�H&��L���Q3� P�J-!��F[��T�L��W����"�J�$e�鋏g�x�<�rHL�k�Ң���QЕ�ժ����IVk�:�B��� �f�}��(�yq>���q�+9�GL{�*�nR~6�W���Iܵ�E����˚i����O̬���(|C��+�T����e����pD��Icd�Hi�|K��al�[�>"	 �@� e|kkLˉS�m�~�߁�z�Y�&W�y/ps6�%p$s��a�hh���rj=�(b�Il�Yc���#�.\�0i�w�=����s��X>�{ȴ�Z=�t�Q�&�����^�?*�{��D�C�(1��m���a�S�]٥h>{��I# ��`�,S�t�&���%X�O*l*��|�	N��-&%��UtT��O/�pũ���z��k��TO`G�������V�\Yé�Md�#��ˎ�[Yk��iV�p�٦��I����ÚE+��O5���B��j��0W��}�	�$�oj{(5�T����}�02+�-O�H�Ϸ~�w |��M����I�3�$�
B��*�ʪ��?�V�-�nAm�͏�X B��4@����2$���v�@*���4T>y��q��� �Z� �y�?�V�bw܇���,�ҡ�j����݋�Ua0<�ߋ��$��@���Coz�ڡ���$w����Ƨ��zVE^j� �V�g~��r�EwŢh!��EY��Hۗ�L���E��,�Z��X<���Z���a^�?Ls{�	7v��h�ϣrʊ�x���%�{�ֹ�8V�:��լz�F(��:U��ִ}�El�P�ODc��oY�:�|޿!$}	1�� ��L������������66f�A���ۦ�)Y��f�|8	��������t�+�0f%�lzT���$!��@��c��ȱ�����*��_����Ͱq-_ɪo�!�s�m��)�I��/D3D3�/���TJʫ~�f�H�c�����5�����6�=V��Vv��Q=�kN�a�Hr���Џ�S��i��N㦋q7O轛M�v������S;�U�tp��[�N6fd��wޒ��j��v���Z����0_!k*��͏�x��t��\S�����k����H�E�3v�����7�V\}WS�w�,a�
<�G�Z��o�W��}!*�pϛGr�����O(����\��,��x�L%;L���M�*RJ �s�4"�.Ծ�,����Q�F��mt4=B�qF=�����,)��d�ɉ����lMcJ��0��/=����XH��4-O�D�M��,��ә��w��#���6>s@h�P�x��`3�,'}���XL����o�x�x��tV����]�lK�c;V����~Z�.w��t��}E.4����m��Z��3$F��@o���2�ϻ%�8�7�N��=6&�v�`�dܠټ�ykg=i%Jr���;�z�"�'oW^'����֌�i�g�g2��V2�Z]#l��f/� ���K�����J\����k(�͌�ш������)� [a.��	�z�E.���u�(MA#É��PG~��°~�D�_��gf���<�7�ȓ/	"���x��?7�(s��Q{`!��'z���l��[5|��r]��)Ԛ�e��*%��̪�:���IMRo���5�������J��#�BD4�f �����˹�������m�����H�9���A
1���?`�����SE���d��eֆSe��4U�3f��c$[�/[��<-H���7�m�@�ry��&v�_�2@�=� �,����BBbgH7F��=lDm�A����
k��1����|#�W�#�h�,~oN{?����n�����Ɍ���Sh�Hrz~�n�Q���.�!�����3��]7�و�H�"�W�r�M�>�ȵ@j(���/���>�x6�̜Fr)`�������?���e̫Xu�)���u����+��uɪK�6�"����t�R�e�'u�������c\��<$#T�}�?M{7�zE�ԣ�=9�pU��!ͅ$�N�j��$D^�ʄ��b	*n�'J��>-i�ߟ?`���,��7�_�DlD�?_<�{%��Zm_)7�j�]	���`�ӹ��fV�� I�C]��+h֔�]T8Ѓru�o⠟^I,d
�-x5c�|�q���:�ř䏃��-�m˚J&�핱<�I-�Z�.$us�9�b���b��Us���bgk���B�����a���=�U���/F���C��Ya?��vϡc����M3����ָ��g�A.bJ�m���-��Ƕ�Cm��g�0��j���P�-�%Kk�I���UT����㩄dF�	h�`=s��>U�A��3�� �Ηu�������"���8���J3�1	��3^]"3����+�*s�T{�p8�̸� ������!R"J�6���y<g�<�O���G�V�C�ޣ���#�-�ի��n2Ʋ#�ߜ��g���wA��$���w�Ũ�uS>��#2�7>i���9om��(�2�|�1د�O�����0b��A�D'�*F�pm\ �j��~ eU���� �إ�PjrN��'��}ɂ��C�Z�/�,C���������y}Þ��P�b���D�v�kz,H�(��I�l$3g�%4��2���#��O�i�����R�V��ix�/�@Z��� [����cpJ�J�,ڔnp�Q�Y�}_�
	�5�#iS�a6o��GGM��=�S�9��[
˥��s���ѧh��E<ˬ��j��g�FHcv���!�:o�GC�0376�\�������vN�چXR���F��Q�gp��ۢ삒�����3�쬜̂��7��B%0k����r��%1�18�u�~ό�#Lu��+&ߜm1������k�|l(2E�q�Q��d�x�q��7�Ǎ��k�x���,0!�����pՁ����/�+V�l��Yj
o;aj�m�U��C��%�vA*֡��,R���6��V�m��4�]�[��s+�*���˖H���+�SFa�I�=�!�
���.�{�����@�W��G6�k��g%�XK�!7'7"�\���]^ug ��,�u{iv�;∖;D�� ����֚��K�C�@����5���V.Ԛ����:���j�((ʞ�1��i^�-ȵ�G\�U��b�	S�����,l��z��d�LE�����j��<A��=r0����,����ʞ��H3	�զ�4DĚ�.NLw�.d��K���Whn�{���\ʐ�j���U��g���AQy~�޼}Q���VH����4Cvj�l�T�����a�K%��E*��V���H\�7���ɇY�բ˗M3Ij
�\��؀dk+���' ��<����,B�;� �vg��Z׬�x�d�����`�OP!,(	������|n�j��`(� �\���7rB[�gt˾��9�a�U�s+��~_̽����)[ �K1�e �K����t�τs�1=�1�x\'wG���2����b�x#��������F/�njEh�phwS��q��,zZ��c����9�b^(��� g�����z'+����V�\�+њ�>G�plE[� U��_ۂc^�z��믮uUL"�5�~�W��ȷ��Kf����Ծ�����U���Zf��~��g��c���̉�e���ƘB�$1�a��6Z2�v'�p���o�����P�E[YӚb���e`��cR�,r�}���TM]!oӪ�h�����>�
�}��e���R�l�y�����j���� ����� #fiw���:<�����q�u��X�I�V@��������pdm����+ǿ��`"��`�A��9qyKt^U� �:���G�����6.�~��<X]�a~(E�~���I�7
���s�3�Oj�ޠyu���=�6�!����9��HwY�x
VWQ����s�.9�y�����u���T ��¾']B��eiuin�H@�D���{%f�_R��5H=ȓ�,N�(a �}5�cb����$w��K@���ecσ�l09/��z��V����ִ�j(�.�(%�X��yl�M'Ÿ4j���L�H�=آ_ե:Z�A	_eȖG����O�ę>pM�i~�K����'�hc\*Aj����7�4=o���w�dL%S�i\J/���fdO���}�Ta���65N��e9� �����:�Vi釆�t�8�]��h�Gи5Y���w�5�ޡ��3`j�9�Å�v
�[mS��}4����(��7R�Q!�PBkjr��!�  V������d(�"�DcV먋Ӣ�Kr�C�:a��ۛTi<	��H���<�ӿ߆�ČR�,Nr�	��a���
aӗ)����R�۳�{�g��K ��Zh�OQ.
�߳*Dp��ɖTz����T�-ѰRd�w��f�����%z�?�kw(?�[�J��"�L���}+W��&�"�D#�Q�e�-�
X��ïlrN������{�TR�m
�f�fb����N�㝘�/��*l�W�pX�_7�ZR;�,��d�*u�^p���P�ع�TB9�qM�{�p�̣�\�PY���n����@��8�����}��g0n�ڶ�hH���g��3s@b������\���u�q�B���-����"S#����2mV�X�:r��;�{]dGR���Q5�N ��Y	��DZ"WkD�t�P�"�
	�>��e��uՈ���p	;٭(�o;�dԛ�ϔ^�ʟ�5�=���� #�ӛ�(�7.�J�j��Zi/Kp*4���>�����1��k���s���2oQGA�;_�JhFM�]��:���SSL���w��xm����*�c�#�8������"��=�2ȏ;J���i�Wǵ`���hx�ɢ{[����̽���A_����yv����O���6#�t��c��G�����!Ey���� IO~]
?e��^6�E�R=����6������(�\�:����95YM`��_�[�( ��_�j���k�ۘQ� ���ON���T���bc	k�,�Q��&|՟��!���z�[��?4���d��3����XOU��Bk���AP�n��f腙��"5:wFX�t�1��_����1K��Ŏ]g�T�ǱCɲ1����NS"�u��Β�hˤ�����kΚ�Ty�'�b�C���,��[sc�N��a����z���&s��;/&�֩������s`>��x|-V�*mzJ�4~�'7���U�R��cc�}�P*$��ne�	����LIL��e�!}�ø��&`�8cO8�ή����mp%С�#�5���4Kk��t�%� f$@Pc����#ޣ.�*�n:��66=����W�I{T�s�l^�2�+a/��U�\$X��n��v��k������$+VHj�>!5B3LG0��M�����¡����w&oR��7� l<O���Q���I�4����'�;<��r� �/�Ŀ�s��Ϯ��-U����K�������0��W�r�kq�5���c��ib�x�Kb��O�⪷u���+1��(��&m^~i��Ѫ-�����3�����^�fF�s��ݔ��C�X��m-E�/�N�c%[�� g�� �á\�n"��3�Wӛ
�O��[�t��+;�*&��S��2Z�f����(G���N�5��ŞXܺeQH}Lh,C�d��
���q�z\a@"itk
�p�w�ܺ������n����T�6��M��.T��ֲ]�6�~��9�5M�392P��e�;a���4�%��V�B�{�@�:���\�
����*�@B�x�2[�������Q'.�P[�(�c��:��3�p�;k'Ik�?��/S2<�Ѷ�`��y���\���Ŋ��o�ps���5Sc��1�]T�7��A��'w�P�����D�IF�����Ò���FX64�'vo������H���, ��f%�l��0�`���8�W#Jg�[�V5�3������|0!�Q��S���������s�??�����3���:YL�!�P�¡��6��d8�}���Ꮃ0R���|;2�6#N��Ĝ��l!l���zMԻ�?�^���+_���9�>)�ak���b8ȴ���!��k�3 Nh読�Y�/�>sDS� |V�
	n��V��c��w
0܊�+!*�����퐛�½1N�O>������`��ؓ��-e�1'H����J����{n���� �±u��['������h3j~I�-��g�
l�L�#��1���4&9�OI釡k�Q
��#\�wԽ�v��O���h"wq���H��JT��8	'6p�=����e=`�\�)�Ŝ��tM��"ݜ��9#�޲�����83���I!����y�S�[��D��5[��G�o�Ry>B��"V�)����E��z���茭z|t��vg�}اՐ}|���q}�	�,�To���mR�7m�`bhآ���w]&ۆJ�H�n[����&�J���EL	4���s��k7nJ�l5eP��9�����/����eA�=Z᧤���s�y�ю��n��r�Q�54��"��c'�Xݳ�|�ِ'�xj���M�R�$���c�)n�a�����f�h�#��wcz��.Y����m$K�d6:������U�
���A�/aȝ�������5�U��^�[�����u�M8�� ��5h�E���A�z7���DxRC�Q(x[[e�uDz0��Tp(4���B{=���?Z�B�եS�

	;���؞�v� G�����O>�E���q
��=�!Ⱦ��t a$��F�#+o��t"øۦ�4���_�,0�\����uC���A?`A�]�����d�� tb���ǕE ����k���'.n��}~��_W�⽨u���b�D�ڼ�\G�w{�g��;��:�iÉ l	�eTG0H��]�3A|c�5G�,7��.L|a��8m�^J	/�=�m%S��V���t{�����v�L����B l2;��}GR��:�Yu��S^ �<j��EF�8u�Ǚ�D��g=���ʑ�*HU�;q)���Q�P1�bԶ�z�#��?B��`kMyR۪�C`��g���Uj^-ǋPFd<�:L]h�:��H��m�uj��IӬ��C�c�Nm������Y2�A�E\*�px����*��P0�a��ʹ��Y.��:o5C賷hFю�E�< ��A�B��|�g�EP�K�瑅��NL�Ξa���? B�U~�z��z����0L��=�!���\�]m���Hh���nK�t�f�Nݦ� �<��:�n!K�S�[������ �5sn�[�%F��ũ���.����G��X���P��Z��)I;b(��G� s<}�hY�8a����� yһQ>���t�0��q��״�s�S|4)(a��,D2� Me'n�Z�{�0c�A$�.���EQ�ت�jB6
��>�Y ^��-
]9F��J��&p���݃s_�{�$��\�t�����"��e�ߜ��WdjJпj+���癪yju� ����A�q�����Z�I�����=����R�t�@�M2�i��j��ح��P�bƺ��vNc&�l��$T-%�S��I�+d\��J�S�L�j�'W�P�7$)w}�h2�o�9�~O$QBA�JV��I)Yh�
���}��a�k�D�~��1��w�ܾ�1ی嚜�}��1���f2�$�;P�c�/���[
n��$Ԝ��m��t��>��1E���\����E�f���5�K\���3��нY$7s���/��#)_��-t%��@=�Ν8�֔�PCĠ2F�W<*��fO���[̂�s쮑�߾�k�9Wa4�z�B �����W�CǺX��Z��c�v��0  ��Y0b�:\��Q���ȹ{}�XEZ0$��B��__����U�X�����ak'��C��</��VDEz�a� &b��6_�RQku��rQ�H�Q+�s@��y�Wzۦz�.�Ň�a�f3�S��=d*��2q<����M��B��j�N����%�>"04�:*�[c�O}�ZV�L3/�y��i�,�'}� *�U�k��l^� �v��cǭ������� 5�$\���$��Q��`��͂>�CD�l��>~�� ���p�0�I�CT*�#z{�xw�K��@�Eh0�%�rA�;����5�>�y8�@&��ϕ2���6x$0�ᡠ��Iߨ�^䍘^:��p����v���5z��b����,������SBE�J��d/P�����f���Γ�P�Å"86I�z3�%#��h��NCjI� <>x��8 "bl�lS�ʗ���BWްE�Z�r��?Ǳ��^]�2���Zh@d��o�>�_����W�ߟ��6F��n�1*�J�~��J��
h2��e���T�_� [P��X�Pᄸ*CW/������Umwn���{+�c���w�5&�\��(���~,D{�#ѝ�P���s��E��qJ�ln٤�[=JL*'P��㾗�S�72�Qw���-:���
��۴"ZM�p����Ɯ� �o���(�f(��:|)X^R!��v�xZ�28	2b
��]UP��[$��H�o��u�e"Ue�BV��
6��>P���<z۞�^Uُ�!�ɷ���_������/�Gro�n]G�O��.�%=p�Y�m���5�	
W��7 �n �B��\�9E�3��4M�m.��,��>i��������zP�(/_ϗTjO����lOJ{M�/RxC6ӵ-^��ISyyGz����U�L]r��l����1�fk�����7Y���xx޺����$���93n�>�;V���P�	6\'�G�Iĕ���rQ&����(���0��Z7�\�=o^�k|�:n7�&�W����![�5	�[�G:G~4밮��W(�@�(��4.�acy�?1��%��Iq��q��m;�J:��7^ N�}o�gom���V�K�D�m�u��NO�}*�¥^}^H��ah]@J�/ۧ���p1��7�#��T=Lr[���J^-J�ј\���A�=���X�p�44u��4���ʚGo�aS�1U�D� ����$��?P}Iu��Wx1D)�����v���7��|���:&�f���I�Iy�+`ko�q�"���MqqѭuR�խ;�k�DR��iۿ�p�$���12gZ�M�I���}��@6Q˘�a�k5g����ت",TY��~��q���/��H���;z�lõ(�Z T �e�hW�tbu�d����b�B�|�`B{Zq���J�9a��`F���>&�Y�n"+,��6�4�H7�Z��8G��ԔA��
Ciyn�f_���>���І7�NӴ]�S�g@��;�ry/���;׹�r*��i���������%)�k�l+H�7�kH��_z�&�/@JK�sfvm�����mnd�#h�|MцA�i�n.�K����3��˘