��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_]�Y��qu�CZ;S3�h4"��p���= ՛���g��j�� �{��v%FɅޅ�C���o2�)/ �~���-_'�1,8���M��1���O&�������P�ۭ�M!�m,h�X2���k�
*���<�Ϗ�]��F'�v�
�CJd�d��6�@�d����QUK��2)ҁYP(�>��2q�J������!�=h��
bz�ΌIY�(����]N�
�U�	�����b(��Q�1 b%W-�5%+/����k	�/E���+=���E�_"�S ���8:���]��Q�[W4ɋ�GO�S���a+����V�K^�U�z9���C���x���j#~�,�<d˶F�·�.�LL�[����3����4�w�V�D�x<=������V
$LЊ�u�͓�Wl+��p���goUi�S(gi
S���Hr�A_��&����[R�e�����hCe����d��֗owS5�Ǒ�a�#�v�i�P9+�:��P��&�JS�yi6��7��㽑�DԪ��$�y�@��4�j`~�[�X�Th�؀�
4%0�н�ێ:�\u�D3L�_{+�=���ET�h��\�N���#�?����p����%S/���L��8�����kZ#�~>
�4v��zZ�'�yu��tk?sS�P�Eu��{�t.�+����9�8gf�"�0�Zm�~����R8��a?��Uh��˓#�*�o'=>�dp��.vPSmv�Yɚ�k_7o	9o�Dh��dʋE.�(9��'�	#��]���v�:�G���)�>w����6�7��kXۂ��/�Vf���p\� �~+�JnY_�^��[ )={ ��#��kS�v1�蚜V���#���듗ܩ�q,+��4I
<�=;��\�	r�_�˟�B`Y��$��D2*T4������7l(�\�n�Z��7+�6&}��Qc$�w�-�`l��N�R+YҢ�Ѳ�͟�e͡��$M ��@$��$�kx��}b�\A�m���<�{��+�X7�t����6��h��34��������Q)L'��4��~����8���J���0#�e���t��=%v�f�_�NI(VL]Vυ�^�Ʀ�,r�&�u4��'����"��痢)Ѡ�+�Y5�ʐ�V� �TZ����a�4C֚��֩6
�oO���7���ob��\�b�(�,�C�HJs�{¨�Ƞ�N�ˁ诇Z�p#�`��:�z!���w��_���v9X�$���]��48:�a��X���3kG�����D���l��qpI�Q�$xX9a����,����!X��W�d&߻Vr#�E��� ����d��%��2��܇pV�)�����J+߃ieE���Jdxd�`�Fzڊe^1I�� !#��!DM�T�*�?at��;��?�=�h��[��BO�	1����Mf�`.��S�L� �2�[�U���u������؞��� ������z:�$2��u� 11����J|�*W���Q� �>�d�>WZ��Q�[z�� <[25%�q�K��I/Ə�9XA���"[�RUE�/B 4U���O
xeF�Ӳ�D�x���{����ۡ�`���Eӱ�'�~�����'�����s�<~���GS��{a���y�0��! k���`«p���2<�W��rKl��?`U�A��=�L,�Z����tlJ� WИc���Qv��V���vs�z.֡�SvX�k�4��N��$��I<iOa���Z-�u �}{N�,��E���@ݢer{��Mᔥ���+��X:��F��ф}����
��?0�J����n!;�>�gKQgy+���䏦U���מ{y���}�32 �3$M7F<4k�VӚf)>=q[p�[�X��ڧ��_|�tK��j�U)�����C�7��h O;�����ď�MΑ�3��x���)������:��A�����15���q�~,����|��g���Ï���B�9:^��%E�E���R�1�iI��4��zY�U�&`����������t&q}�f��	fU�bP}Y�pә�X���i{O�;u��==�����c����V|�z��MDD�S98�Z�2��	T��5����AѺ_P��B2�93��^Y�mׯd�'|�nR���vv޴V��sg"V�Yf��-�~8��.�3����+rF�mk5� �E�Y��
KV���ě��ׄ���*˯2��9��A�g7�j��y_����k�9����*1QH.0R!N�3���N}�������g��:���g`��rf�fN��Nn�v��W޳y�UR���C�2J�Y���J�Q^%���P�#�F<�f`8t�I��M7~�ޯ�t$�]]n�i�}0�Ĳ:W���kďav����a'��3�W�0��L�f��CXo%��
��:���J�!�Z��8�6Q��r
Z@F��*[�����Ƣ ea�n;ܥ�G�cܻb��ۄ652�����Ф��4����?	��@���A� c~��!���~����x#�u0�Y��������TV�ñg\ø�y�֝Fm�g�s�)��OL%E����F-Q��/?�������RL��H��a��~�'Ƀ+��̹&f��KE���o�v��\�A�����㫮�Z��8�eoh�U:a�s�~j��[�o�Wל/��"�%��{͑��\�?��	�ZcB�Y7L^܁>"#�Z|��>ut'w$�o�^��@�n3j����1���i��e]�U�����ݗ����Sf�!����+�N�mݷ<�f�B`�����>X}5����:�ʁ$���*e83~v���Y�I~�H]���րF[=a1�1["ĝ�!`�@�62C	�<3��}�|�;��y
��Ӽ��`r4r'e�r0���e�b�dӋ|���w�o% R9L�d�؇�>3��]�ӱx[�؆[�ͨLO�G�O��1O�%h� ��!�FӦ�O���T4��Y@��9l�~{�UZ������ĲH�2��vy���FY�}Uh�_
fSI,��/k{�C�5�c6i?ՙ�?��9
*	l*�K݅�qy�ww�m����A�2��q�/	Ί����q��� |Ծ[��wW���/|n�P=o�;~5�
	�.����Q
 �CL�j�Q2�U���ڕRT�
�:�5����[��e�I�A݁g��O$��:��T�1>��t��|������t��б!��H�fu���Z#z{X��Y��q�<�X����1���d�!��@8�ܐz��![PD*T��WœW9iB��d�"�Y�ҙa?Ǣj	�#&K�b6�ձ
�։Ol޵ۖ���a�ʣE9�H�W��-\�F5gT��@��x;����[�|y��lL�Պ4m�X�����Ý����I����;Q���y�:��7y����ד�j]�?�p�Ψ��|�e��t�FbB'rXSP��t$�MH�w+;�}2�yY�	Pr���3���i�`���G�f��w��A��e��u_���~�S��zX�M����;���|T��&�5H\߇�NjXpR��.'�}v!p����}tp|��l�-`�<='6&65�)8��"��2�-��S���m'�\9�pK�,k�-W����&úI~ �M�
;�"���kfBVWk���,'	�b�Os�Tv^���B�*���@|��+5I���Eh���^�V`#�P:��;�vf���7&�����+[ ���}kVf��n�o�����YPf&�;���G��)w�M�>\!��I������^,� ��{!e��]T�y��3W�-ߦ8QN+d--�l��0��f���4�D#	��#�`�li�HK���.ڿTM^��M�Yxl�I^�s�Q��P}Ñ��$���/�f�1���M.cC]������z��r9Z�v��~�ik�����y�ؿ�M���,
�0<:~��'${�i��Q���[����P�  ]sz]�L��!�� �?�RQ��q��ѨL��T�����(�]:}�F�'�p��ݍ��/�m�d�\��&j#a�2���Qt��Qf���r�$a�C��"��f���f>��q�SfX��K�giN��lB��� M�8�P#<ڋu����?����]�"�[�'.!l�Zƚ�;]mfe����*2��k��
u_��à�~V�㜦�W.|��9A �g[4�88'y�WJgbR��5����Z��cĦ �����m�J,��2D������S&���ɣbe�h�N�fS�cHu���{�|zRp׷��D�3���8J��7��y�U<B�6s�ʊ���:&6���ȉ�Rm]4�w�
$����v�F���P�\��i-�^e�[pӀB�WO�]��������7�� ��Roy��ĨHlaF.�d>"FIcӅ+Эcpf�a��N�_��l��{�*b�c�gv�4��}JN�6�e���~Or�J��A__%r4�P�+�L���lv;B�L��;"˝u2�Wؓ�͙�a�g�\bbh��K�?�Q�
� 7ӕl��_0c�?St��za5.�8 �~�ԍ�;V�Ɏn�(=�Y� U�i�nȢ7�h
ъ����M���A��t�ֿ��A��r��W�/fY!*P��X2;n$	K�e9w�����zҵy����ng�V��8%*�T���̮j�w��u.bY$$#�>��~͙f�٭��6Z!F2�š��9����E?�G�4�r�M��i0F�ݼNEM[�5m ��S�'��-E¦�2?��217�[�4�1�h�a4d�L�+O������FZ���9u6�w���[<o!^�6B�sI��>��*�@�al�������ض[��Axu�P�N+�e�&	 O�����=�4A�^�� �4�J��]#xHh��z���*�zl�T�ll���y�/�^���,}��{��yD�\r�'�n�-��v����ϻp�V6���o=O�ɑ�ᛷ�`=��vY��C�FR��8�.>%w��a���mVV�bI�j�x'o(���&���Mh� ����e���4)u���̮��u^H*�,���K��������1�t�9��K�*X$䁐:�"J%n>\�D��U?*��"4��;��-�d���@	�G����qL�z~��)A|Ҙ�4�2������'�F�֢��i��� }�r�.O7�A߹!���]3�h�����	��?��Ѐ����;5��N�����݋�m�6N�'�׌�G4�S}ܹ#pC�ƍ�*�e�Ʉ,g������m]�1^o8��d��ގ;��g�ႆ	^�16i���gUs��t7�׃��N�T1�&	쏣|�ꀧ�>*������\C����Jp|�fr��j��A�4��Z��G�4��PMP��au�u�\@��/bK�+��,����)]D_�1Tʓ���A�J�ܷl��V!���/ ��0�E��
J8�Ec<�&��ⳞI�``WF����z0ȍ��ܑe�/�*9Kt!��ݨ}� �t��a�h�����Ҿ�����.�����<'e�MS�M�x�ۗ�J)��EI�nL^y�bϗ)���榯��/)u�]-|`�[�}ad��:F,R�T�����!�j���ˑz�W�Xf���F�c/K����ߴ����G��x����P�W}zq3�j0�����W�p�����^���x�wA�Xv�r�*�cM��9����7
��R�uZ�@��9�Õ� %ͅi{�������DCseo!KLKS=�}.���P���\$Ӆsf�lP.�~.:�q�9iL�4� ��mȅ�,G-髱9�����t���~�K�`6@aE�	�nA��aT&X����f9�u�uG�Fh\1�q܇h�捌��6��S�!Ջ�u6��-m�˹/0az����?
�I�^�e���,35�]�o�~�9ej�X��ܷPy%�!�e����gܽf�� �A��RX��Js%�����c>�z�?�P��U�os`������%�R��RspIr�P]L�D���+4��}d-K~��$:�Gb�%"�y��A���Z�������)-�o!�T�]˵��¼�G���QY��+�t��pS�ؘPEU��>�-�vy|����aQbp�vX�_|z9J�$�v�#����B���I����`IK4�xG����Z�'D�!t��_:��9*��PR���F��M�](�6�h��箶�If���ʊߣM�)@�@�<�\ځS6=$�W���Ӣ�-��(�c��B$�a}ޝ���
�yX���A{��
p���:s΂��N��8�&Xo��rC:q3uOa�M�Jpj�K�t���p�5�"����Q�n�a�F��W��B�z*���\�o�YLc�Zd�7)�M��fiKV����Z�	��)k�1�C��1"C�f�-c�*�hw�U���mS��*�g����jڽkHU�۷��}^��U�����W;��������j�5��Hg���x\q�y�5������ƭ�Mƶ��F��p�OC�H�M�5�:��?qܔ��y
z�x>�$1�
�¨�U�e������=��}��~��ま�Y!��Bx
��v#��!a�-����7�r��zM��o������	q��޾��13�نGͫ�O�m�8�wf3�~;p�HV"("c������ �J���~��f#*����E])U'j�:��E��Hl�˞vɁ<�ONZn.��j��	�,A8Vr�+�J���C ��"͡vT��΄�?�@��RT�׶���d��"n�l������ZY���p��g����"�hvЌ`�p:�@-�T�C]hV���h���෱W� �|A-��(��L�a�������l�<�0"�a�k�f�!�7#1�t"�kĮ�� ��]���/�"�	
m�u!�qX�+{�yO�꾫�+'�$�wS;�R����J�k�����l�5��A~�ɼpn�+��z��9 (3�%V�l/�������b �S����hP涣3~B�;>�{ҿW�	-Jq����ɠ�$!u�f�7���5�O�:�j�'��ی`3��&P����@�<��fR�����S���N^@TAp0�!i']u�ā:�H��<v+�9j�]m���?dJ\���H'F���9��X�8�,��V0�J�HB�j{[�U���'2�AdU^ш��P&�죥Gʞ��Yj�p�S�����ѹ̇���1ṵ=T܍TŤ5_%�X�G�FTHľ��5B��7i6uzP-ϯP��/�§�#@В�a��a��ӽ
��o}}]/��,�v�K��.�L~��Q
M��8ȓ�=`a1������Ҹ����Ut�䥆��A��0���*$�K#�FeU3�=��*#�:�/��-�S�8�թ6��*7o����;�I����F2���Ã�Mykk'��u@!"�z������JlZ�t�c70�����.I J�גdm���iH�S8��l޶��3��cӾ��Ģf(2b�˘����SKg5��EV(�d��CL�� �I�L����Fvi���aq��B�
�����=�f��gtq�C��XC4�B���1��û
XHR����&�h�]%��W�`�#���h}9�v ��BZK�δ8:5L�w��llG��桦~(�7����$Z��(IY���j��	�p��˅-n�0QQ���^�ϔ8�<T�����R���r3
/�GcB2�M	HCb�>\�EH�#�և�+����GN4?\E3L]	�7D��_���lϙUҸ�X�qt��)�6qR ����6���ʴ��V�Zr�Wut���jI���$ץoAU,\)dp���=�t�4�@��� ����<��M����kb��V��[_8C�x=!��?��|��ֲ{�>�/�S�و<G�a"�)��r{`�.�C7�:���B�V~Ӱ��L
�(�S� ���
�o�~t��<�,k�ł:�_m=�{jr�Q��o����5�R����c�,L�<�/��|��u��oN5��XS9��)��!a�� �N?��ya���2�7	'2m��S���^TqkU������XHP��t!y�_��Q�ն���<�+�S�J����ǭ�Bm���1��ދ��x�ݵ*MTG�[ � tr�Εz�`8-��a1h�*&2S��/�Wu�)�#ϼ��{D��h����QL�����; x;�4W�7D�����#w{8L�F.92rE�P(���/�W$1���.�S=�"LO�u��GX��s���}���q�A�Ahi��v�ūm�J��	Sr�+�Պ��GC
n�@��B}������������S j����!�b:��wEx\� }�AZ��Q�ڗ<��tq�"��ȑ}%a{s���5l
�ol��� G����Ĭ? J���g>$>^KY�/���[�+EJ}�9���+�[���쬗�_unGPŶ|۷g��G�>�),�f�3��m?Y.��xӗ%!�g�胻*Em-�5C�E�i�"��xU���tf�����%��/
������k]�44ҹ)oT��ހ
8V���T��.���>D���w���d��i2w�VC��ft�Fz�V��k\�/g���'���0����o��K߁9
�:�Q�e���'/�hI4���`�X���4�1�Xb����\�,͘��p�~�D*q��'{!HP�\�V$Y@��fM'jc^ep=U��(tU
}�e�\�H������4����![�ǵ��g�;�����,�Ӌ
 ���/�t)_�]g_��d��=Cǁ4a�53�m�����S'�Q.�/��;N5�5r7�D�+d��P���9`G(��0!)���l��еބ�!�����yy89�3,c��fɉ��k��O�t{Ձ���� �GNs!O_�S[�`�7�uA~�* gs�K����-m��{!p��t�F�SXv���$2h�O�B��
ɇ����'){]S�qo�3���)���`�ʯ�M��Q�+�>X�_S%£q/��!V;�[@�Im'�J�¢7�J�`��O�/��^���;!i��ʪ���ň~�v\L�	��}ބz�|�.��1�I˥]����&h�C���M=�f'��Ȑ�����Vl�!�:"6qM �m�������x�a�^����SE��� �z�5:6O�b����y	`wTk�F��>!QO���[���V�]�b�]T�1�����|1F��G����Y)�ˮQ��U�Xk8�킁�V��Mw��*
�qj#�M[�K�(Q�i���H��&�A�g����I��Yc:�`'�#k3�u�>�wPe<!F"�)P�3-qW�B(�<;s$Q�Yk@�Jh*�d����cP�Q���`���#�{���I�
��ޱv�|�H)����;�{�1�1�6ދ8�]�6��y¡0�j�զ�[1)N��?f��h�³�F�M�Ҥ#<t2H����.`N���q8��Z6��
���	�z�+��v�#S[#*Mwn���(�&�ծ*o9_����+3J��͋V�?�,��7�tF��WAk�V��l���Uf�k�O8B���0շQ�z�f��umW��a)�)_��#��`G: �L �w�iOi�/u�+/��Å������B����=;Z&�~Ѡ��Q�!���Ұ����\�bQ��.�A	PMKӛ��ag�����.�YED�0C���c2;�#�`�]�$��v>��D�u�Q,��`_��Eƅ�Zħh����&Y���*n�iVv�j舲������[m�qf�M,i��$�%���c�ŕ�eH}d�k>s_]<Y;���2��L-��c����ϔm2}�;H�Il�.|:���ɞ�Ŧf����Õ�?��.������T�G�K�ܱ$�7�8!�J��9VWT�ڐh�\����k7�3a�!7�rM �hZa����%�.PX��R�x��EI��L5LŎ���F[ׅ*��X8� ��N�n�=��*ibK:���l�{Sd��×%�ێh��ć�P ��iu�KɰH��|�6��k	'|Ntd.�CZW�bc�i0%yB���L^�($e)/M�e{�Oh��-?;�GB�G�#�A����R��<�e��
.\�*YH�#���Q�� "�>R����k,S�E^zNW��L��GT���x�b	)1���7@A�$�ܗ���B�<�.��k;tƫ��l��&H��`�#H�8ꂩ�h�O)=������c��y��ğe8�=lS��H�Ά����l�G����%D�܁���N�~q|:�X���#Ǻ������3���$lL���)�8���������o�R��m�#�Ӯ�'�����T�x0s�Z��<���9dúA�'��?eH{_~}Y�����)V�Z�?���y8�<��Bـx�X��"%��\U���	������o��V��H��xd�ϔ��m�"�o�'�dB�x��M�""|����bGi4�/I����.M���ޟE��X\���R�?�����Պ>�4���**�I�.�Q2Y����:��r[:���wT���e����k�2�
H:�7�r?b4�JyP$���~'馺�8�c��ތz�5�ڹ�T"nv�k�`�  ��/�E�LS�8A�~�4}���Y��]�X�ٝ@�Y� ��\��ӌ�J��l^��}��͝)��,��[')�+$�6k��XcJ���>E|{3s5��$~u���'���p?p��Z�g5��aVL�^Sa(t���+�]C�a��� ,�ՍH��^�N
y�=0,kC�~x�b�"K&�SD��w��X�j�R��3E\頧h�ѩ���Y�c�D�0��>�w!��h���o���4h'Ǣh�C VM��������woF�n�
�_Q:�\M8�0CX�t�F�%��[�R�}��?��ZY�a�u'OΞ��w^#8e/�趸�G�d���D:�&��t*� h��I���ur���Ƭ�퍴�X�l�m��ku,z3֏���r�{�Ȍu6|_��u�@C�������~����,�̜=!�[�gs�(����Ü��Z&(^�ӷ}gbQG)M�n�^�ߣ�Q���Qx�R0�8=)����xx
�s�J�[U��H�MxFT�h��P��r���;�'�.���=^��� �rr��8�ļ��:�D�z��Q����K��C�
�
Rf��~eU��~��m�����`��f^��s>Π�߯�C"�ծ98���=	{����#*��la��7V,�L����ѥ�VX}��7-<40�hu�lI�>)��*���-����h#=�sS�2��4�/� �2b&�je�#�F.��q��PB��?d�����n�S��̈́Ĵ�޿�����z��Ϟb'N7V�)Ɛ���@����6�����vz� ��X�l�?)�Y�k��_����:R�z$y�;Ω�)�ڠcůp��/�|op@���J\6�Nx�&�N[�tKRgn/f��=����Y@����5'3�D�Gq�$��#��ǀ��J3�Ṓ�M�[ȣML�bNg��]��"f�\�)v��o݊�XBx����W��&�b���et~����+%���z{��-�]nd�y�;X������L�_'��q̵�9�*�#5��O�=6��r�3��Um�`	�� Tmw�|�R������T���գne�ߟ?bBp(��%eFԀ�0��B��6>@��=�����fA�GOƺu���x����aYc9Ei'W&NY��m�1��w϶�\��/�"<����ir�����o��y���-�a�Nz ���u?��u~?kc��q�?�
�e��C%Q6�͟�Q-��^�H'��-�������Zn-�rKv�߉�/�ّ�(�4u��o�b���U��3�e��Y��7M"gnu�{q�ep% }�x��pk=z���c��ŋ�b�DJm�%���{�{���U�a��0��0�D�I�>�wI�r��%q�ɾM��e�E-r�I��f�	��e��k)����I�������=5Q���
�=�%ݢ.��@��U5y���)N_�G��W��>��z��(������QBMO�]�8��H1|`��r+�j�E��O���c�^���C���ZZC�!X��`Ņ�2RG���!����Z��,9&�8g�o�s�5܉L(W<Z 6~�
שF�O��u��,�N��K�U�[�Lck��=dхLVA!mt$F�6Z4�0_�j�}�h��,�Ē��{����,�k�H�ە�8#OgmQL��1��J��{q,س�i��>0xU.)�e�ɥ&�q��s��*;�Z<��B�~0c���?��
s&���&aa��*6�r	�E��%�/��ݰ��� s�JE�ÄG|��"̆�8~D��2-֩�Pw�ѹ��+����H�,d�v1�� ��J����N�#�"��D����P�\�1��4�S�ܽ&f��5�� ��s��	<G��Vg�vÕmp��e��dJ1.�y+�m�l�Ol6��l���u���$G�'��L����J@	�9X����U��	�c�:,��H4�S5��ׁ��.�.h��0�BIh;
�5�t�7��un� �v��i��V"�8Fpt�s-\���3��\��q��Ӆ��ٌu� �m�(8kr�.۰�1ԊG�C�;{t-��H5� �b�Y{p��:�B���Oo���c2���/X�t͂<G6�-��QG|K
��KR���o��N���LM9���u.j^�G��U���J�;_a38J�R�Uw
�?U�e3�,PP��H�նHA�Xx�$z�򄍙<	F�9T霕P�rA������	��"DJ=�T����*:0i��<`��^�ә��q�~uG�E����JS~΂� ��SC��9�	��⯌!���K(N��bmST�8�[���$.���c������<z���.����� ��wx�%���9:*�%�� ��Ѧ�Y�v�dϴ�wm�nǘ���]-c�8�n�a��յ�g�����ڀ�Z���R	�9H�`V<w:���W�=y��2 ����Ў�]��!�p(]�1C��6vE	I��W���8�V������A��a�n|Ř�0RSŪ�wct�`R)��2$>M�y�K�xβ���6�S>�H����@��Qֹ��a���x~�����+*�yA���Z1�[d��v�[�Oe����M4�O/�H�uFTZ�Xc�����ƻ�*��R.����n�ɵ3��x������E}�/ƌL���2Z�+�G���5i�^ �r�����4������V�%�S,!�<�W@�ZA�"���.�������;)>�ʸ������$s��}��1N%g�
��-�q(ʅNf�˸���e1t����6s0�ܹOۓy2�%��oR��������'�}YU��7�̜c�큌��3�Ɣ����&'=�NPGqm�N�9C*���yTR������UpE�;�oK�Ap���b� �[7�Ս�[0� �vS�����v+ ��Z���]�oj���/EF�1�?���,w@?7K�w�Uiu@J��(��?qj3[�a�7�ݹ�����u5=]�$�*�#���AK``
��;v9�g��6�Ә;a��;R�g�oN'��d��%ª ����p�])�s�¯l�Jj���9!]^j��ī����웣;�f�Í�:�{j�	�|ϖV��S�Eι\��څ�Ѭ)�'5���{��T�7�������%��o�A�[���v�}%�}˄���Ĭ����\���.��ܖ�9B�'y�����(�{��Ϊ�ۋ��
kX+�X��a�9�(������Y�"�~�b�9Z� @z����J�'�E�vzu?h�~�B��k��
�%)����XD�3�T
�vR2�(lv��I�#ًЮ���ٖ�B�$��R��q��KN\�n}H�J�W*�٧�pp�F�<iX�}3iZ	��
�z	h��d�&�Qt�ˬU֏����f�Sk0X"g��7	�_��k`
U_�qˊd�#��Ǻ|�)�⹝�A=�gA@N2z$q1�M(cEhy?0l�����7PF��](�BQ���W!l�p��*�*��N��k�Z�mX43��1R�p�@�����ds�o���3vW���]�*_-�f׹�JL��&����m�����W����>���!*���d�˽p���'+�]ӨZ�fĠ�Yw���vH�y'�'�ʓӧ����m	�|��ԫ��F�S��Ǥsq?�q��{{RϿ�*�����
���#����َ��X�cm��
��l4 kN������Sc�O�,DȬ�I"��x�a�[I�בd�3#�h,�����`�H���=c<S�cE�s�b�i�<m��np�Le��E.���\���2>�49�$�C�F��K��A�d���xAǖ8�,kw{,w�� ��/=�Oe���
R������a�
*h
�5���]ucߔ&j�Z�-�c��2?��b����1U��"���CG@S<�����}l���76zÈ_5v���BՀ�^M�޷RT����UZ�=6�@"H�#�*�U�C���������� ��pY}� ����,M����V.�N��UH� �w���Ճ��E�1�n?7@�1�yD->�M�D��@*ŭ�k1�x!co����^ŶP�8h1�F/�U�ٞrP��܁��Y9�����gXm�4�:�e�vB����H�Q�iw"�N�uU%70�>��#�yh�o6Ք(�x$���*�(��N�M�� ��oy{�+����m%4z8��ݹ*�� Nǹ^'/zurX\�(�$Z�F��Ts�<
�O*���	�G�7���~w�ԛe��܎kx�Y)Z�Y��y*M�����Ivr�����U��{�T�����w�r0 �M�F/f]p� ���0M�YߖP�8:u�Ț�ВM��R�t����e}{<��/� ��Ycݶ��)p���@8������WPER\�� �&��{d��i���}��K˞����ß�QӲš������Ɍ@q7'�c	�1�=�{��~U;�i�I���ʝ2�Y�����a��-�\?���FI��p��L���S�}�DQ���.�e�Y�b�X�g��Cz���P�t�b�h�#C��GZ�,���4C�����Jr�`���%��H}� sZ��	��͹paZ~*�WYƉS�����*Q��1�S0��=FY�x�w?�� ����|Ρ�����9o�~*��u����o����>�O+�yF��ո��@�W�C���:�A|fΜ�3ݽX��f�!H��x���>���0]6td�1�k�b��鵝�N�ɉg��1��$ 󖌙V�I��a�~�e��itZY�i�@��3�w�Ik>��2|L�i�����5�bp^�b��AA�ƎQtC�4�;2���},ڤ�&�ˣ+|�m2���%�߸8]�&&��P�B�7]�V�D�ٸ��e����D�Q(s�m6@�*�˃>� ���^`z
�C���k'�F�����C/퍒��-ZD��d�n��'E5r'������}�E�b\W|�e�T]����j��31��S�� �# ����#e�X�N�cJ�M��Q���V��@s���l�়����vw�,�z�?��.]ǂ�7�O��8/��E�_gs��@(��lv���>x{j��O ;y'��6����9V6#Xke����v�[�Lq�n�%m��bm	!�gYM�;Tٔm�>z59��k����\�+�����3��'�<�d��E���N�x���H�q������K�ܲ!��v�D6�`~��Po����7B���a��{~��z+�W����3k��	R�'wy�̦�6�������69��(��=d�gĝx�#�x"��E���*=�T��Q1C	s����}�A���ƌ��46�$����q���'3�esx���m�
A�氯=����Uq�(��p�ɀ�����S8d9
�\�0��:�F<M�&�MYnc:�M�kKɪ�b�������{��iE6K���$� �VGڕK��=�S��>T#<�6���K��-B�G���*H�O)��m��W���F�SwJ�(�r"�6*+��
�#�����B�-/��R�����i3�V�����ɨWNÎD�ScEt��ӃA�aXO�6x�(�B�1�-�� 
?����3�����hnɴj��:�E���A��V:��(��6���3M�T�bV��fC��`F��eZ�k�W�+�#�"���X@A0b�T�� �}�(}J���b,Ǭs��� y�+W�\֟@�mtA�4�=e�I�}5{�K@��ɧ���*����ʧ�AVik��Z1"���I��=և�:�q"����UU��P}Ƅ�8��s\�,u�����$̛�]h��aJ����Oa��6 ��?����.���!#��Ȣ��T��^�Ynb6u���7�1u	�9v�	���ld�2�Cz=ۤ6òN�)�(b����ـ�瑠����؊q��@�	̤�+���Q��B�A���� 70����0�0����(���at�؂6�u=�`�`7��B���,�xQU�6�r��=�Py9�0jEӡ.U�5��W��Qr";*�;�V�����8�a��H�p���9��o3�s���b�C��nZFXi�M�F[ɓ]� 	T��mƸ����p�9�BF!߿�Є�uD�S_�9��f��r�Ȩ>�qʟ�:�C'MEH�q(0�&���Av!O�$'",r�)���V@�}��v�B`�Fq��LPv�	Br��g�#�)_����
��P��$�	rf\6�E�'��lr��&�6U:���΅�iN�S2��!8��;�����ӁK	M��c�O��1�rj�N���pf3�&+�����7�$�ϧb�`�T"=G�$}��a��n��q�'J��被$}/��%�<�Z���Xu�2�7�����7� ���΋��B���O-[��I��.���-���,�CGgq���c�8힦A�^O�|�#�fۘa>n�>0\��
ڽ-���+]틕F��<\,ޅ�4���`fRx�M&4��_5ڟ���$��L��	�K	@�V�v(:�2�Z���u��'����c>�6�uJY��8�%���L�u��"m�j
��,
*�?+�Q���p�%�^ �)Xv�(f���`r����g���>��7�$Z9��mgn2K^(��C�p�mv7�*e�MK�)���{8�5>�F@f�x���g����������� @ ����W�Z�k�K뛇\Q���$1|�5�jEhu3�IЃcT*�?�]������#�����f�'%>����p/1A��%��e@����B�2�\"?��c2E��J�EW��4!MA%�6y��9��	}��P	
R�_ʪ�r���x]�!�����v:�{OP��_k�u�aX�g�ǅ�@� ��?�(��4/��И����!��,>�3��݂g��)��g!�9m��q�D���~�ȏ~�i���%J��D�%�`����+}{�b��c׫�r����eȍ8��&�p��X*�^�����y*w��G޼�����1 1��vNw��9q�N!����gN��e��V�6y@ɖ�)%G�f�К(��tK���"�֪4&��?�$����d�@�"��ix��C��j�NiZ~�c����{�$R`a�� �ut}<�@��� � �^$>h�"�5cT�� �~xFz���Y���0��Q�j�� ~?g{���)�4�C�ߢώ�� #n3@��s����pw|+�#t U�z���*����ď���%���@��z\u�J�K/�=<�8+��Wv����׀)ĠVB���(gw&�@!0x0�'n�F�W���q��%�.ƛ��I^��J�)f�C���U�6�iHqr���6�?A�R�L\��GHT�ݞ�.]���hƝ���67gdJwb1ɃX1����L-ޤ9Y���7��\&�d��\U�{o�����_s⨓#��e���ħΎ�J�n����K0�˾���O=a҉NL�䆫%�q�J�s��RAq�-����H���}�Fu����\�������HoGi��*m���~�s���v�Z��~GK8�v�W3���v���;�jșu$ю̎,C�أ�yd
���<�z�~Җ�`|)Y�8-�g (�BFЗ�d��l��x~��PT0�o�;�.p����r���2� ρ���;��T���k��I��sRp�*�l�hOK��x3�8P�G�ZV��ܙ�-yL��p�������Ɯ߰](�<H.Y7��<��o���ó@�=�M��Ch�9�d=n��v�ޱ�W4� ��3Q�]bC1� �?���-��~����x��g�K�k�љkjl�����s��x�?�~�!CB> ��Ѫʐ{��W~� 2��2��M��ɮJ���c_.&�w7��c�wI#���"��k/�W����<
�~�+j��f僄��^�,�+�tw'�.Z��yp9 �[- �˖���� �ځ�i��j��v�&cS������a�x���u�����9�����j�ћᎬ9�g��G�4���n73���ʯ�0��#(U�BϪ I'��"�����2�]������4�T9I����" �x�+��H��v˶vLKّ4�?�/������dR0#Uǭږ������\`k�����4�.^/�`�u6zv�uΚlw텒��	�8�C'&�&�	�*�FI�N�[�i�R���#����R( by�j��zS��2�5F4�������fPv��'k�Y�YD�/�A��S�y�����eS.a���6��$��f�ҏa'��Ƀ+�����n�"b�'	Yvd��F䢃5!/r�R�����ܭ/9��Z�H���m�/�G�iF~�+b�-�*��k0�V�P&D�a�� Y�ާG�� {��ۢ�����1�*6WJ,�Q\Q ���7�(��}?����;�pr����W�b@���+IZ�����+a(� ������'�J2G���U���)�ν�� �^����K��k��s}�?O�o=Tv4�k�ɵS���j���e�2�rƣi���@����[���d���}kH��R��%�dt��� ��	�TQO���ΪB�x@��w-R�z4]vX8�4P�1�9?���U@�f�@�tx���ax੾�h�]��O{��L.��G,U':���m�N/{��T��p�9���{��	�d^���1 WYA]�J\=�0�)�!V�J��}LQI�o�#mΨx�		�����.�Yq����xA��7��O�/zH��_��?�@�a/���w����:�E9� +�)9�q)X}�V�0'����K��%�9����AK0��c謠,��H����S�Dп�;��-ɳ��M~Ъ��7�<h�𐈙��޲��){��>�/ק\�Q�,a��!��i��"jb���l��Q燇�Q�{�NP�Ϝ�a9�!E"eT�����U&�L0>~K*�Gn���.�Q��#ɣ�-���q�eRQ��	�s!��R?�1D�7��:�`#��ݮն���A��}�JŔ����_�Z�����ƛf�s&���kQ;\N>h�~��-;�7��r��|����6B-��ԡ9��Z�F��������w(��6v�*4NP؄����b���7�L"���Hz��������������8�8��1�[
�b�AX$4��զy �#��3���@[��y���gQQ�	����,�"fw�bW��B��]�J�JQ!]��@�X���H�pXiP�@�� !�ݛ#+�#|5��a�Z���b���V�s�><������������>�h�φ�:��.~Z���8�cb�	�)-���XZE�Dx�|�S0��-�@�ҳ�ϩ�(:��G�����ѽ M{����+�X�O��":3���<<���Ӛ4����AɤB��s�y�a�-�����uenmwg%/bM�֫��zƃ)�b��F�|��K�KB�"Y��&wc._�>V4�T��m��K�U��C/�%s�e���}�I�~*�]�8��6�Z�Ⱥ������ʔRmk�h�x������v�Jw�\�����c�߯mߦ�z\>˖+�F7h�s
����;��p+{&-���.��1+����5��� ��͙!�>n�q���&��4�ԝ|ޏC@h��-�=�c��=��ײ��Ó��X%`W!����.}�$��&�ۗ�v0{ְ�l�je�]�4�]��~8m�(]�=�7b՟��X☲���&8����F���yD�st���ҽ�Vp�]"��>�'>���Qއ�����O��bpUQ��4��FERv��^�M,�����r��JM�_O�5H�3��Ԇ>�{߾!��Y�7x�S��t��d�i�����Vb�Ì��r�$[�Y�2W�E>���C�܉��?���8B��X�="�|=x�;v�x70s�(��)�&�U��K��W\a���+7Ê�qf��f��m�+�k)�DU����M�a�l�J�����p�b�/�6=ﬆ�L�ء�[(��ܮ�����SX�|�'>�z��C�1�ߜ��3G#�E<D�dW��G�� ���"y&,���e<wS���-����}.��v�^k7���K��۝�����Jx!�A{vT`��C���H1�SF�w9!*+2]�~Cp<2�VHNW�ߟF���|���9N^��`Z��O������Zp^��)�i����_��U���ٲ�� )�����ŭ�2�i�}�d�$|�c0�
�c��Q㒸'��Q\~}>�,4��j�.� h�2(�i�U��*?�8�&�6�Ɨ�R ��Rm0un)YOV�����hN'�m�,	ݛ>� rW�K�E��@6��2�����#�8ѳ�sG8c�=���#���<8��Z.�8~p*5�QF�7���̜�m���(�^'�]�>�4�Fd�Q; ��3��6��Ȏ�*�g~�SM<��`�ᮁd��,��Fݝ1��o����jZmI���4D��џ{ }oIo�V���7A�� ��¹�i�zVa�cm򽽅��C1?����m<��%Bz�w�W/�L��fr`�G�b��&}F�gI���cF�!��B�B[͉Oh)<ƴ�u�W~W�l7�Z��o�ڠ�AgY?i,o^I�,��.p�Ȍ�c4��-����g���(L�
�Z����Zk(��iG��(i��!���P�xo�s1��=�g�����Gb�%�I2��bD�CX�@z|mUȱVd��sI,;ìN���O�����5�i�t?��Z�K9���V�ַU{ ������ApO��i��U�fu��~��w���s1��N��t���^��^�
<�x�=�7Dx!I7�v�`q�t{{�G;{�5��.���/�*��BCP��0�au�yK�=���^,��|�my%�7������0���%|�=�M�ݕ:^����]wbFѪG�I��Z�%��.��{ruv��K��f�;�ji`��5�3�KWcaa	>$���U���,m��`�'Ĉ�`���)q~2\D�m���\l��<�A<��ԞF3����T�5��F�7ܧ��5��l;�p�	��E�\7�}��q%k|'���6��@��NK�*�u����>½ӄ�(��]�=�Z	���|����Dh���%G�����!'�r�s���@`M�_����ڜO𗌜"�jY�P�1�Vh{��H�}}B^:�~��ѓO`��Q��K���~!�0�@���)��zz[�,ف��%�{�-=YH<��������a��z�6�����)�u"��i���J裝!�Ǳb_T��ӟv&�{Q�iW�I�]��Y����Lđ)_)��]�7O�vY9)�F	r�����i�cQ&�b�D���I�N�T�fr*���Ci�w���G�}d��3��<'.�TY~S׺,ns(q1�M��.��=��F�⥘|����ͧ�d1�T���iƱV7~�l�W�ӑ��&V�>���J�}D�X?Y��H1�r6@.P��%2��2�Xc(P�<6O ��y�9����o�hR�7�l��'�k:�6���u�znꪾy.���4����É-K}�@�Sю�ُ�n��V�^�^���k�>��[���Y��y\(��!�m�.#a���D����!`@�>�U�md��@��a�:�Z�z�XB+4�����I��'��#X������`k5{��=,��!��?S�󌩖y�oӱ;��������'H���=��ev(����!@�?�4<f�?�(��L&��Ĥ���D��B�ۧ�CP>Z]��c��7�[��^�p�L9}_�E������e�}9!��
hyn��F^�)�xS�)S�d78�=�.��X�����o�ԇ��Zt,eg��A][4��p����E7�})8I?�(\K?(�X:�>VZR���[��|�ú�*�5}����R�Nm�Ao>�j[' ��P\$�4�����hP��)Ds����^-͑�߻Z��D����Њ_.���i@�����\�ĐPO㫲*��CȄN�1RC/"�F�j���l@
0�ƌ�QW�sPf_ ���M�l�UV�^�ԡ�'���ɬ�����>-�љZ�uP)IlS>hB�O��C�Hr�Q�.���� h�v[k���" 	"�HQ(P$�AHv�xi����_)!�X����n����������$�?�mk������r���YȢ!ʩm�=6��a9 �X$�f�ۉ�5#�������:i��"��j�o+�&�:R#'2�c~Ǟ@��,����p)� �^�t$���Q�3��,��H �ui�Ȋ��oс�tK�}����,0ͳ����L��F����/{Ь�tV��'��2h(iwX���Q_�q8Wg�@g?��Bi�>O椑�����0I/XF��ҹ�o���L��s�@]s�@��(�7w�E2ɳ������#�>��� ,�#�ώ9=�����ݧ����ۀ�r���M� *R�<$F�q-�G(�`5ϒj��QF����쓎��pU]�H�Z��E�9�L7�x�
��N{�Σ`YUe�.b4�X�@�1�:����f �T��o�����L�?��*ֆ9���il�d�J�9Mz��
�f�9_��1ݣ������`�a<��+0P��;c�N=���.HR�����m�h-�Oo�*��-�� �u:�%�����jfpib�|����=���r۪F!����be���d�Y �`L
�Ap�]�Y?[(�/zIH<S��cb��@A	�C�!����=��_�jGM�}�9ድ"SQ��l�/L��M�򚙵L��<�� ���Z���?N�B<�`��_]W�*XU��΀�64�o��R�2 �p[�#d���W��l���S����,B?�c��'��x�h�#����?�ZnS?E��Gq4)���+��;���q_8�BF��q��ڧ�77��a�;��hؤ@��19���4^�e2�S�~�3F���mQRe�o�r�������"�!H�w�_��l����k'��7�c�@Z`	�?pH��z<�r{]啶VM��V��o������y�9�3/fe����看#�W��X�_gIa�YC��h)���1Gs���6-��,P�lm���
�:8 �4Fd�c��á/Ӗ:L8��� ����p�U���p��;�g���ģȣQ8u�7O����O{�^�R�C��9r������I����tq���D�ʶ�}}p�%��5�X�i8��DX�Mph���K�
+*��IV��I��L�=�����|h�������zO���v�mިۗ�'��E�cx�C�(}v=���lW[R�Z�PgV��!_�>d�p��qYT�3��QW�=�t,K�iqZ��u�{@��բ�ѩ��&�Dֽ�"b��Kj�j��!δ�O��1I�������*����hw���`(&��4����¡�@��n�[��^��X^��`.��t	d����w�04����<=��]���!�h8ަ$���.v(:�Q3����2�\���Q�y�]�]*��d��ί�*���ۋ I��Z�4#��T�]y��"yD���H���__H����B����Yp'�e�(#!o�*N��E���_z�ZyO���z��q4�
�aec��Jg'0c��9��:�b�����%j1i��r�^k"^{���1����x˞�E1Xsh�`�g�iuŷd xR#3�L�:����[E�S��"s�"�;�?�2�ze�nC��]-/����������;�BZ��/��X�-��ׂG��,��f�пo'��J���N���ᱟ?^! ���4�y~w��mȅ�q�E䜑s�gP5��8m�`�@BS��[����9y� 0��r$��v���U�0��b�;�%u$A���K
�Q��p�b�S�]�LmD�s܌ DP�]jv���D>����ir׮�T���Ҳt	���Q�zm͈�iώ"ff����_S<�]��zi΍b^�,�Yb9�����} 7���Z�s��<���Rv;��]�A�`��zT��Ey6G��i���t89�4��2~�PW�����>��h�h�
���҅�o%ҧ��:�6�F��1/8HC>p�4F�W�-x��Z�� C7[8�$�q)wQ{Pb�I��W_��%�Z�x�F7�kF�ct�9�pu,��.m�G �������VZ��*��lu�M��eA��k�jcM/����=6���\bjiQ&�s���?^��M7���Q|S�4u�m�p��rFm R��;��K��	�H��l-���2��KU�k�T���L�1?3��5����Y{�$�T$�9ԉ�-S�鄩8q���b��R���Po*��\i7\\2::,8�
�v�q5 ���ڏ廎5aU�~�n>�9������_�`S�SX5A�w3�-�9��W"Y22[xm���$?{��Lܠx.��Q(�4W&ř�ߙ"�����롔Ez�)������Ё�w�Ǜ|J�j�w�C�#�=���-2���XƄU�Ճ�SE@�+9k���\d-P�d�w�N��D�H�[�W�a��/V�wt�5Nv�Xf�=�%�$���ǧ�Y��'�ѝ�[�d�S�<�x8j�n����˗C*P�F�Ϭ(��_�84Q��Ev�\�a0����˩[����J��_�ɼ1㟠~��0�θ7��g��$�5�܍opX�S�՝�t�Kq�^�O`�@B�9J�|Ah¢���:	���}!j#���&W�lѝn�^����g�^��~&������ x�)ڲ"Jb� f��)�
��z߇�Dq��Q0d�]��'��L��AvU���FQv��1�ݦj����n=�޸�m܌.����,�y����k<�T\�Z^�4n)E���}��=S��
���M������t���l��"\ͨ�5��7� �e��2� ⣝���k�����e��۹k�76K�h���8���K4����E�J(Mb���燌
	S��D�=�%v��ۍ�Js�w�.��Tv��k�t#��`��u2n��mg��cSxN}Ey� -�8j�
Ԕ�"�zM�ӧ�ޜ 8ù,e�U৮s�xnz@D8��"�Ɵ?��X-C1u�%mS�[W�j���UQ��/��\� mU�K��aP��H��r�Q���r}p��huIp��;ߐ��I��݇N��M�Q<�,I!�ٹa�C5:�Mg�R^Ыd�ˏP2@�9������D�\���\S%	Z,�&���n�!�7ޞ-s^ o�C
J=���zsT7a}�/�����
�TuSvἺ����w�'##S_H@�'3#���Kv�yqD�b�v�{x%�����n�Y�_��M~�>Z�6!��\����q�@�Yx��a��OJ�g���	�9,\����^�{�1�p"��%����oUO�Z��b/���0�7��%�նHo#�9��r�ҕ�OކxW�2ZO }}ƌ��b�#�8)���V�e�]��%E=�\�Xz6���	Sl��sH��)8r���U�zl�gE �h��w�h�����)'�̾�!y�Ib��a +�m)ysn���M�����Vl�����(�&�/��������Κ���F����B�ϊ@ꁈ��9�N�R�J����C�P?r9V�'��<T0��d*���"�Z�� :�U����hV҂�RW���]�<js��Z����L$g��R8��CT��񦿠`�m�8r�Α�Bʺ�,��^��M#<�'>YM00Ji���C.��CL����[a. �]�t 	'��� ��U��	�U�13��èqX�r
����;O�F�:�y����=���N��X�����vô�FL�A�\��mt �+�-� ��B�S�*�,#r�+cqN�V�����g�N�e�Țn��q�|�p�a��#�Q�$$��l��ؔHz����ߝj���ׂL�A�� ߁�ܪ��pj������Ӝ�b^�ݙ'�h�&�K�"|uNT��
m��(Qqo�X����:���=̬Z�;�k[��C�hz_}����Y��}4��
Q���N��Is	"�?�c1�`4��5�yچ�`�ʀQ0�aZ�AC�3��}�c���qع=+x���X�{+4Q�F��@���U�g-뀝��e�c��Rؑ�vk���$�4\A4+��Bd1�Gk��Ű-J�I���^��dwk������@�a�s���(ZĽ�}�ꎅz��9��ybɌ��p�o�c2�ϝ=a����
��"?<��*\ǈ�t8���q1��Oo�������f����\�V�@ }�	�U�����Vv�'��x��S�5M��ҥ9М̚��������5Ɏ<�`̀9SV]�0qLxmR�	l���'�o*~��R���ʲ�4>���7K8a3�,�����A�����<h�]��"�����9ۀYE���A����J34M�`�H�l����2l*1�3�{	�����p�$HIdcv7�V�;'��#�Og䖢m����3GP,c�|3� g�@���2�a_}L�=oz��xA�D#�{�������װ��d�
7H�H��6���kBw��cF�K-3S��i)�[2�V�k�	!�8zEƅ�0�R��uP�e'�$w���I��,�AA;.<�'1j���K
߂ß7H�O�����v�!�C�	�+��������n垇���w��w�k�tP`	��P"K���\�����e�����3����r^ٵ����k=4�>�_�K��d��I�������$�m5;=g�e"Y��N��E�|`���\��(�������]�/��%AƏn�;=w�ި�Mt:���� ���e�F�bv���^�O��]������߽D	O�$��c��4��9���kf�sPВ��+��X���KD`���u�;H��Prw���܏����PE��"h�<֣Z�P�gc��j�b�V$I':�!��"���?#��z!W�����cI�S�� ���}%C;���Zl����l@FÛQĵ^]�ג�֖`�(�-?H����D��5ǂ�<����L�H'��kސ�&�'��'�',���'w۵�i�#�Ҝ��v�;Q�G�l����!Q�m�?~�߱X������ڌȗ����ۂM1g�EƚU!��p5HM6~��$F�� S�!��lt�����Ջ%>�DJW�>�W�t�"��Աi����u�F�$v����Ud��~��"|R>�v��4{f�`����C��Sb=�"�O�����b�r�o��c4����e�� �T;����<�%O@�D�|������J(�l��	�0t�LO��*(.o��}7c~bӳ�´Y�b�J�!��>?T�65(�Z�P� ��Y�S%-T��A��j��Ew(�J�S{�Oh�9И����;HV���Z\͖����������s�
�i ��?�Dj��U�����Q������s�.n�j�zh���»,�;�%RY��B��=�u<�hkP"����O5�JA��ݜ��y,|��Ta/��ڴTGIK��	vl��x�:sz�_��A=ni���y6Lx��RK�Gb��t�<ϵf@%�
�������on)��g�맥]�<���S�$�<`ĔN�+{�/�DݶĐ�v�����Zd��%�x)/����k���R�Rܐ��� 7����6B�Ġb`Ld�J<��Ȣ�r��l�ch�i��C���?|�c\88�#u�X��:_<h�������G�!���w��K-3`Q��m��n�)'#c�R��5�R�,��t�1H�q1�:,�Yj	T~��H�)ͨ���1ΓǄ��� D���̡F�� dwAr\�Ơd�'*���V�}yB�8��и��l���,�h�ä��@� ;Bdu���q�^�ƭ�_�L��F�qf��R���8����B^I�� ���yF�+	Q�V{i1�?{��A5���us��i �)}B��eݍ]�A����]!<"����M
���,,��%����u,]��ط�#�焜a3z��W�*��Je�_�ekB����"���Ȗ\��V�)���l�K�2C�IȝiqSs3 ����zx���,<8ʤ�M���$���.��剗F*������s��0�Z1o��D�>�_ۄ���i\����D�:�m,ѻv�d�}�{�[t��R}���	9w�^�A��$��<IH��cO��c��UuY*�r�};�s�h�ɐzo&�֌���a�Vu����V�W;��g�&-B������}��=� odq�|p��k^T`{-O�xi'rl˶���˩���Z�1�d�QKBɘ�ɵ��
Ӗ}��9I8T��w9G�W���V����	b!�9�<����c:��7��a����8��֕�]��o�	|��wW���}�>O���@Co �0%%r	��!���$��Y&^�×ݫ9ɀ|º���,���%�B@gg�"�jc�/Ow�%���*B7T:Ǖ���r�cґO�4�5��&���~�|�nJ����ȃ�`Dѵ!�Sz��I���������p�R��O������L��.��B#{���⾯�Y�m�p7�{��?��nr>#�w��=��Y�����'s
�x8+�j>����g�P<�Iٜ�]I�sU*��������Y�Lf}
gBlN�����A'�˒Ł��(��[�)��{e�(���y��K͋\Rc�J��0� ��c�o�%jX�]�Y�Y�����)Ӗ�G5�j�%'�t��.hb��9��<�� M]�^"]C�U3�W��9�*V�����Q<���^�jT���&��Y.�ܡ�4��9���{V��y��*�V+�2#j�$�*�#��Yxؓa�J�Q̋�7w�9;5��"�\3�z~{/q"1ա�}�f���v�t	'z����R�Y0b��p�/��e����NΟ F��� ���G��P�������3�C������2�(�d"&��oWv�u��
�n�͝d(�;�3J�5�	�S�-����7q�W_rH�����y��Y�0=5��0Ӌ��?������'�܋��n��?�7%����:t�L��doY�����Z�"�[�$�	sJ��45F�q� e��Ed+A3��JN�m��O�x���p��G���lΉå����aR7F<�Î\���g�z�X5���Ű�^������]�W���i@]
���D��_a2�e�V��a���q�ڷu	o�}�T�|��F5�'4�w��y��Y��h�A�'qݜ��mX�jW����p4k"V�qF��_+���e�I�OH1\�˱>���e��G�Zt �_�X�K56Y4�F���>��x��>'"�0ûͶ !?,�����\�6�m?��:˳q(�D��4pq�I����}�X�\�#5�U�%ݮyȕ��M]�_M��Յ@ȍ'c���'Y'p� ��_�#=Z8��\u��{� NK�D�]o�C�z��gz+`uː��T�_w��D�L��ߖ6VP��ֳQr���k$x�ְ�t��@9b'�Y��q��i�ϑ�7�YW^�#k���ZK�2p���^�$Z6�|<M4��ӭ҂����3ǖ�!�!�N�Ԩ�=%�J�I���i��Bƹ��MlX�1��A��3�`�,�M~�I���n�4�1#����G��z9e+�8��!B쓐h�>群�TE�t	V�<PX���d�s#��N���^�U���ϰ�3��˔(?��ۨ�J P� Yױ����R�qݗ��L��%�s�j/�(\���残��J ^� �_�X�����0)�no@h������[���F J�q��@y�'�=o���!�T��(E������\���]� �/43nG>Ԃ>Ք�����ONc�k(�ɞ���fY���02��Um�`Q�}~��m������؏ы���V+�/m=�Y�Y���*<�����|?�%dM�}�0 �9�/Q����&��Z+܀��B��"X-��G�C��[��dv��fs�v�y᠁��,�y����-�jV7��� ������"��1j4\$�E���c3{���b�Nl�"`¤>fӲ���*P������y��F����%��	�N��TP� i�<!�#��.��kn�>h���Q�uf1���#�C��Z�:�����z"�/��ڳ%��d1�7�)M�8<(y#�{��� ?�D���׻�&X�PM�(j��s;����Ӓ��f�J��ß�N�aڋ]K�a��K�w<��(�S=sW����cG� �����4k�đG��3;}#wz���	A<u�c��G��q���p�c���WCϖ}��@5��u"|y����j��B����c�;��K�o<Q���s�Z�wϒ���\enGs?H�_�[!�����#�m��Lv����"�$g������;��\w�>,cGb�Y��N-��Mf��*��,�gEBP�O�4��@?Ld�a�����E�F�����	����;��%��ܧItS���*|�Mi�.b/���2�\�@4���を�o%_�2+������q����J#v�P��Gԫ{V�ܞ6!�[>@�)�x&�9���V���"�ۼ��_��Mt ����	����}Y^���+����C㏌�Q���7��G�$m�A	T��c�d���-L"�5=���K�m���U;��#CƐR��2W Y{�^!��Khĺ�߻d�����Xm�t��t��(������_�Ѓ�/}���:5}%İ!v��g1��A��D
%��������Uz<s�������Ê�<���Oe�L"�ݘ�=usO�kK���J<	f`06�:���-
�7V�������۳��`��#l��)z���x�?�N�9���I7�f[����{��kӹ�6���Hr{���Η�"<���k�w�l�@O,�e����������x���s����Pe4+F�n���I%E�Ts��Q㏧�Cs17$ G������g��[q+s��+�/Z�G� ��^��j	!�T�i�����ӥ��3���˹sK`��·��_�]�l��!a�qN�ǬmQ�*��1���=�"��]�8fp�����2���
��kн��� ۞���������-p}o��Ľ��]�g���Ģ��0����=:�w�ۥ���(����i��hA��̱����5-�)^����6�<F
�ݑ& ��}<%�	���}pP��b �����v`�
Pl~��� ���t��`X�9����N(�c�S��X��M�E�B��x���vKlb>�R�o�O.� ��a\��*���lB��=���6�Rr����P�Lo�R¶���\�f��J�r�G5@�(���5�P~h.X�~b�	����_�{6������ک�/�C���c5�fc����\c=y��Wȟ\�k�@�w����9��B�l4U�ʳ�c�N�[r������ڋ]i�����Z��#QG[���_�f ��w��B�����*%Y�Z��m��=��H0X�
8��wUڨ%��w&�!�`�v�tѸ6�|��zC!������w��L�$�^���U���Ė �g��eE��a�0��m���ء�7���@��1���e����ߌt�e,��Ky`�s�Nԋ,�k	3ދ���@�y�5������ B6jS2�8b�i|�	����dur
�]��#��4q�
� ����0�E�\l�n�F}�@�틀Nw\��u՛3�s�w��K�SHiQo�نz��*(ʭW�+�l}�~�|�[�;�>L����~�]���$�)A���D̳�R���K@Ș$ɑ
yhJ:��EYg���U�iY-��|쟅b+�B׺��������@H@)o~ ��*�����+���L�H�	j=�*�gLȜ&ҩ0W�	m�D�{��Ykɒ�96��$E�~�R�E=���]�j.�o��J>�O=����oE����g���oꪉÎ`t8�qU�>������.2:�6�@xL�b���Sv&m�[�_ $�@
�&Bf���*�C��X�5��˰��D��2���j+�j���O>�����i�NE ��2@,v<pj.��"��/�8�п��nۼ�6X}Z�;�~��|z_�,��{dݴ���0{�!��
��%��I��g��2����?� ٛ;�Fa�e����Y�foU��om<�/#5�KE�CR��M5�����y�Nw����y�R�1���o:*e�����i��0��xp�+���6AH��/#`�֖���4�Pޫ͔�%7�.hϸ�.=ոk�b�m��'!3�-�㱌��t�mJv�0>_ !HE�	f��A&���L���}��o%��&�����1���N��5T���?�߽>�+b�Q���@mx�j��5�B�i:�%�&iz���T˙���6�J��A.Q�3{錾[��(u��`�c��[ |qi��;]���z���z���JG�k��pe s>�ěW���[~���{�A��a��H&���z<N�~�pDi[.���z��Nl�ߪ"�A�xP�R$��[���{��PI;�i��>�<��ժ#�Q(��k�-�m_i�1�-�7r"5�/J=����dO���������S�԰n����i 1�Hg�	V^��64��:�ć�>I����a���e���%~W��ܬ
�+S����r��p+g��m��ѷ��%8� �gV.P�%��E���l����d٦�������[L�3��[<h
h�w^��$4F�����(UV���mPLG�4��iXý�~���_�VsI�8>�d2����2��l�߱�ؤf�V�w�����Na��6�\��;d�=j�h�!:Z
7#5�����&���?�NC@.�^Y�����*��#?�~E�"u�M��G �&^ˆ1���d!k�显.��2�����c#�E���k�cd�غp%{��z�&�Xe�v���$��3S��%����/�79��b)ʡj�p��æIc�z�X�ZOm���3�R�"zq����fꖺq���j��d=
G��q�F���i�=�5�n1W����2�R����k��P�`��D�|1��:#�@��6S����.�K&	�!�^�P�UE{9�"����O =Q��u��D2{��J�j��i�`��i.��!Ad-�A�sL�y�2Z�ٰh��A����6���H�2�t�I�P�؍�G ������{����8_�����Cn���T�uU���N��"��D�j�
#�
d�[�R����
�J�^�g���ց\��� NL^��|��p0M3��|75s]��Z��L`L�A[�v��D�9��d?�"=�����grv�V4��G�M�U WE"�Fi`� ������ؓ�˻�\�u��I��lq��;Pq�w�@"��&�T�lɼȻk��j�x��H��<"�G�l ���J��zs֛'�|�F^T'V�M�1�3�����l��K�ȡ�7�����*;-���>[z������[|�<L�5�X�]�ĳ�������ֱ!
���Z)�OH���i��7Н��r�گ�/+LQOq̥���?��|�)�2�8i4�)��� *{aZ~���O��▧�C߉��c~�=���u�X׆Y}_�����8�U��]�p��8���=�Z A�������]�}�>/h���8j����f����E���&O�qO�&E����]��U����ͯE�=�P��nG�.�_�Whțt�ڃ�����,�E>��{��v_5�B�����P��j>1ٵț��B�-��@B|�k�nZ|4�кV�dv��*&�Y������,©l������T�����^9��J��-qP-�n�h��ˢy5������/2y.I�4�/��mF���\���uR��O_�7Лo�֌+	G$ƶ8�|C��G�b�~�D)u:A�W$;�l ��p����<G�dmCj�`��-t���e���#+!Lr��1���U+�����נ/�Z���%����������﫴NA�<���l��|<�M%�"�+%){�^��xaP�ugȲ�x"���MW���]��d7Q��Ê��d^p��^ذ')������M*�RJٌ�t9��ݏӨ�Z�~�G�?��C�����	��
���#l�&�pe�i)��vH���8���X, �B-n!�St�)�{ey5�h��(�$�b���5_�_6��JǮ��ӳ�v��y�I㚆���A��UJ�W���o��������(��X��������G�E�1�[\�"i����t��`5%�'m?���⇆���3�Z�ߣ0Z���F�v��@�y�>)zn��L��G�Z��t�yܒs��L��?�m�qr��@��m
� k��w\��)�&!�wڲEl[_�T��p�J�����)�B��V���:{�ly�����W�ח̺(�O��m���p�,kp���t�g�Rk��g���L��-�\#���� ����iִ�(��>����Rk�R�ݎ���䤪s�
��񯅏���8;�J�*p��?%�R��^����IW�W%�E��9r�h�T� �:"*([:-���k��%�	y<��
x����V�����$�����<-(Ō�6fz_m5a��6�\.h
�-i��ל	�(-�ݜP7Gy�Ĉѕ����5U⛿�CL�����1rC�a[�P����T_n���+�椫�B�^�{�H���;����NOB��_	|��D5?��R!hխ���~u��ʉ��mP(:�5���҃�2.��<�NU\��$�*�8@ ��l��`eU�h�BO���2��~`�cF��l����@\Og�x+���< �]F�(5��HV����I��>_���:�7�\![�;�BD �r\�������rA�G��R����\V��I��(�U�u?B�Ι���Y���x:�F�AG�����#k
33[�0����-��P(��cp����J�9N����A�C?�v�١npڿ����[�Ut���t>��^tn�CIГ�(0���� z� ���3������'����4�+�g��"�'$c�����o�K@��}���ڒҟ�h��ݲ����+�P0S�J������'A@K E���£��GB�
��^�!��L��v����R�|�����w-�>]VI��U��-�<��I�&����ȫ~-%՟0l����V��(In�q謷����
�k��"�rÓ�s��&r-�J�r)W��,�Riᬻ[���"D�����3l�X%���(���W
��D���y�������w��&(2	V?p\d��6��Ǥ؟ҩ��A<=$SL/ųF�WL*m��%���B���Z{�R7��9�wa��a��|�bJ��酿J8V=��@n���z먫����f�4�{	�@s|V����`�Hъ��n����r�ݴ�GQ�rq��RD���f�e2$1�'�ل|ISN����0�nj�F����A_C�BE-�]��3I�+��+D$�y��R=��������7��:��rz�<��Dz��o��i8�5ʟ��:�`r�5|<�V�گ�9�d��٤Uɒf �vz���ک_A�g;��UM�٬)��F�2���G���wp��5�j[n��v�>�&���� �4]����l˒��K~�M������f_O�dv��)�2��~�?�*��8q���਺O��\�˩@�iA����?�y�
�&�F������"r���E�Ǫp.0��>ԳP��khmzt��hK#wޏ��)Z�x>�(�Yh�j$�%Y�R2b� ���r������k?�<r�2�|'��������x���o���?�>R�R��05����t�	�w�RtP�:�`�L2!�h�y��]�����^�*2⦓�L�y��n�zA��=-v�\��� ق�7S��*q����t�\��%����#��wsɯUn"�=�TÈ<�&�<�j���WX�Ø�4~?Ui��� ;��$�CH���8?�0$��Y�6��9���z���K,��Mj�L�!��H���m'웖1;!�)����7�����q��W��M�zt��!�j��w��R��a�kp�8��]����9l3��}iר��p��aw����ms�Hq���x�˽�ߓǥ�l�_y�]P�։�Y��O\��6-�q�L��X*�{�m��7�X�r�&��M�-��x��P�f#ٌ�WWRo�� $DD�6��C11�r��w^&,�y3�C������+Y�����e����r��cRb��ݾk��Z<$��ւ����"B�Üd/=4ҙ��8�"zC�����t�I��a�0�e��E4=Ӓ"'J�B��Hw��!��Zub2�e&Ǒ�
����)���f/'U��6Ɣ�m�����'~�!y)tb8s���gY��
��d0��;��\�V.O���*6t�Ά����n�R�tgK��y�j�:U�?��g�������u\/��q�쭼�'�!n ?,�Ρ}3A	��0��M�<3�C�˥
ù��e�8��b�ض��=���]�r/���D>n���9��S�Ӱ7����O�Z'��Ô��irSMA�H��`;ԇ��O�����PX��1���w���q����V�Ţ���zvi�Y�.7�g,N �{y.#��ruF��J�c��F�+F�]7�Hq�����^P��e�U�|b�����Q���R\#��1��KJ���W�8�\x=�h�/QW��{o�]ek��$&���E�<�7�p۠A���c��\�v_���v,`N���槀���\�v5n7�՜��ڶ���ܖ� 'g�BQ�hSY�P�H[s^9�+�8Nc	��+����̖��ZУ� �N�'*L�n��Bw.��^N�z"����8�>�'����P��9��=�۰h���Ʉ��5g�qP��r�m�bc�Em*�>�،������N���竍�&1m���i�f��0�����cy�7�]֭��0�i��_#i3$kl�I�y?�_��	��2Ok~�b5{�1�8p1Q!?,-� �����}�q�G<;c�p��v�6v��@g1ؑ�#ߥ�HҨ+�C0x��,o�>S�E�<���%~A~�.6炌�ۈB�~J�Xqܣ��+��)��~s�N�%�=�!����cTUۚ���|�鴽E��W��5�cy�٭�O�װ�b���Y�)��XAM��2_�G����3��z�h�թ&Z2���-���[����������������u;��8���n6/J	�K���C�_��R,�4p{�K
����P� {���V�e�o>�X6ş
ӏ}F�xzV�]�����Q�߬G���aE�n��3�D6�7E=8C�ġ^z���#[mD�������_ҹ�K�c$&����&��:�)%�`�p ��Fd�ʺ��}d�gk=���E3�*�E��7��yg�"e�=��Wl�Oa�"����8��������oXlʙ�	(�Q����yG��s�go\��k��y�(�>�  ��ܑ0��_�w�tl���>u�?��f	�������k��X������^k��r���7��ӻ�⦦E�p��#�6�����-HteH�}�������3���9%�cg��~nv�kU��	T�~s�l�����.7Fƪ*�$���P;�8Sw���yȄ�1��Qg;�Gو�ƲB�%��\��/����SV"��5)�@Q63����� ��CC���
޵�������wv��N)N��E��$�����}����۴G_�_j���Rչ�71y��} ���p��e���4�]�HGtcq^rUĐ��{�@Z}J�m�**x�E`#v*Zw���2?�j-�e�B¬]�>��Kd�g�_"l��+6��Y��(H��$ØQ�z�c`��vM�}CeZ��������4��Q͝�/1em��,��-	Q;-�w]��~У
!-	��8^��VuD��1�e��X����1s�$7�©#�$B�������8��N9s�ͭy���D�y����<��Ĩ�a��p����}+���}b?�t�z��+6��$9��Q� �|�v��ĩ��I��4F*�kCT�Vx���Ɖ��Px���=C�ڱ�h<7�8��UP����ŗYr�/>��+���4Z��x����-sU����u��侶$ųz��Ξ�VO��Ԡ �٭�o�T��������t����>�▽+�ܑ�^ծF��^�ȟ�������I��1�����'��0V���^<$͐�R�,j¯�t;p����)�ɋ����K�9ި�~�Q����AөZ���,b�������5���[h6�g��^{m!a����_�G�q�h$!�Ps[�4�$���
�xR͐�-�3��H1�:���|ׯ��ӣ�R�)���ִ�}��^ 3{�5���M/<���6ʯ�5��hi(�(�8Q���~SՉo� �Z���zS%�I5d�0x�l��`^�%AN���BK��L�����hnj=7��)0���p=e��	v�i�o�~"���E�b-��t�|���m�A�$:H�S�z�h��H8�8�K酪9��z�b/���}Q���-o2��s�|�����F�C;\=����+��^c�=m1�]�[v��� M��l
� ?��)��G�;�f���S�`��k5�J�f��ǩ��� ߾ت0 ���eߥ�r�����/�%��=��N����.#%��<�I� T&P�!���3u�����g�( ���8��A���!`��G��HZ6Y9���&�"|���Ych/��;n [�59�����Ha���>��|Prp��Lx/�h��1=�)a�̻b ����@�C��h{��o ��% ����swH2Z��6�2n$�b�'Nh��#�c�9�5����U���8d$(���9O�	��4T|Jt7�ry�ol�2��̀�/	�,0�4����v�*��ly�O�6ѽcsiz�Qb��/T���J`P�	:r\��)�n��W�ѱ�O��XX�9�_�sx�=�ziz�����`8a2R��#=�]l0�^��Ke��Ky�;K�� -_��v����݇B/1��
��2 !���9MM�2ek���-h�0r)��k���x������4�������u��n�ހ:Ɠꘉ_w�Uת^��{����)�0���*��� T�d����jzk���9���E@~6�Μ?^������8�&[)*�ƻ��<����v��~�a�c�!�2T�v�`f \_#o+a�n؎��FIvۍZ��3��_�WS�)ڒ)����m�_�S��;���2�bT�?	�x���Z<ӈ�2����RKGr�M�$SG�I��6.=��@�)[2�D�g����X�)�����_Uw��N}Ǹ��ύ���vE��֚�79�}F
C��T����e�_W��Lê	���݃��A%/�SL��ҝ���	��+����/H���5��!߂.ޣ��r�n�A甍F��)���~&.��o��Y��Y�z#"�s����u�y��~�m�������rTM�4���a��b�H�:��8������֧>d��3�U��;4�w�$�s �ɽ�	�_�$ܫi	�}�6��t�������b���n�����'�)�3�K��˚'�$Qc�m�2����(�ʪ���:>��uy�U�}��X�*MI�M]lR�"w��F�pD)9��C��yS}�~YN��ۭ[�y0"���&C$����3�M9��ǰ�i�/'4�[L�	ٳ��	��a���x!�(�S�@|���
 �1�eaغz�oS� �Si�+��7��F3nL�-T�0�/áo��9=Iq@R��	�Ɨ�y��[��v6���oQ���d5 �r9P�;C6Y)$��lM�����W���������-��6j"b�&�P�?pK��7�)C�J�sP3��V@�ɶ��;q��b<^��x�I��Ve0 �祻ޅ�p�Wty��ϵ���j<��x�\�9��d�pjZtrꮭ[�5�-�n�#c��,l�l����5L>[(���Fb��2��+���#���n�.o�"Oڻ�����q-V�r^��}�(7x,�|�`�� �&C����� �y�,���(%��G������M�;Z��{�4s��&N�����%�E��/�s�L2�f:ˉ@�3�~H���%�ۊSc��t��qG�2�c1���+�7WrgZE���+R,�8�L�hʒs��x�]����N1��1B���%0���
��R��"���?!)��Ԏ(�,Z�	8k|��;/c eJG����\��:���<�Lb0����&����)k��S(¤ޱH���>NI�*H�$Z�	Ew�<��$�Ђ[��V�6i�t>�a���޺�.��ј�k�:L��d�H�+�D����&��[��B]��O��:��g�՜�=$p�ꝋ��'�����C�{�q�X�e����� ��pB��O�ku���V�.�p�Cj~T�)������n�� �9. (��D` ���]6�̎�I+ڗ�
�3u?��@D�v1����T�s�Qo��&��c8�t�6s_�B3�)+���e�:�;0��$6�I�z}�_�k�,C���Eb�Т�Tne���5��C;��
�W��L$D6�wE�0�.�+;
������ұb}_��T��g"�j�b���.o�n~. J�?1�w����-"֫��1����`EJ(K�i���H��K���J�2E�{���	[���cu#��kȍ���]ŗ���{�R��1��i�Rׅ	ۍT]����I��v��>0%�;�^vgf5�^�ٕ����@f
%A�)����$^M@��Z��FA�k�����Z&���CM{۽ҩa�J�F	�W�>&Df��(d{��[�iV�O���.`�@?@��<B�q�'gJ�D��Y׆�%�=�����;���5�d͚�j�د�
ı�|����z؅�䰃+-ת��I�J(�~k9L���F_��M��DIR��<��Z!-��U�]���I{�+V���d�My0�#��H�}VW�B�0�Â�B�}�[S�rA�T+K�c=:M��RiP���
Y�:�[�l�����zK�w"�Xv²�q�u5TQ 9	E����"�p�?�X-4�� S�k�U�a>md��Ja��<3� Ok�o��.ԥa����}��^����V�:�y0�v�R�_��Kr�[E���ZW�A���Ĺ�˹W7{��ǧa85��q��m�/rr:<%9�s��{q�p�b-�@7�N��b��?�Y>����葱��\�L��$\�-Q0(*Z�*�J�џ�^Ht���`�ׄ��7)��I6J!��������!kL0���R������/�1H_u1A�&C��Z!�,���+zÓ3�k�	>A��̃�R�uc����5z���-��0PxcI�X���@�)�	z��)��2l�8^��_��cd�ᢠ����`�4�ȍC�"h�K2�G���M{�9ҰQΕQ�sHG^a�h�6�˽��)��R{4BGj��a�@xy�n��e��.��QƝ�V�u��ׇ���}q���L�{��_��B^���K1b�w�F�8&m��I��ɞc�������B��_��N����5L#6̚]
}�`".A@"��/�,�}
'Hǫ�^}�JAd�[@�*���([��RCYŏe^«�
V,��v�q 2��� �Z]$o>���\0,�\��_ib����2wŌK�S���ڷ`S��أ�f7yٷ�`&Ȅ���[� D�0���]lc���{���\�g��'�����Z�ׇ�Iˍ�m۽�sƁ�A�LN�n��t�^-����)\o��vӨ���t׎'��Z�Z9q����ܔF֜[ܳ�m[&5
Ƈ#����Yu�� LQ�wƯD���-�7��\�02��b�w�'�/��=���{��f�U:5/&a����{3J�?Z\�lj��x>���D	�w���@ˡ'1Dy1�cHo�ᦢ���>�NN�AFh�q����uWtW[�� �a֒q�Qr.q,�m������()��,z��̠�ygy�8/)~�{өԢ�y�k��F�-���Pf�
qL\���h�ʔ;'�(�5v���Q�:,�\�����ܖ��GuY��+�\��]M0����TW��<��<�WWҫ��5&ޒ{+�>t�md�RA9������@,HN{��b�|fx!��乆j��Z�@���q�=hxN��"�ث��o6�ҝŽY�%S޳�{��D%i�O�Y��fM��ĔY�;uǁ�ȏ���|��ޱ*n5�����^�K�Lt	�������V?el^�9i^E�V�9�@�v�td���� }W� ��;E���M\h�|�FM�. C�b�;1a�Z\�n���DD��i�q1����;>$Oµ!�}���+=m1������񘡜��*�?�Bӑ�u��Y���*��i���d�F/M�-.�x�3�O7��F��}�`��rL���\����h-�8�f]c����z�� ��n������e�,�H�aA*�D�bts��@���s�[DV��V*H�i���ѷY�_�_�/Q�2�޴f�Mx�z�f��>����T�`����	�N}Z��1�1i�0g�9^�qoJ�;�!?i�I_��a����d�N� �UwE)ϱ�kFER1��]��u������y��R[��@������n>�z��[;I� �$3���R͏���J��y�%�A��j�>C~��~l.���S��� ��A҆�Sl��z:W�Y@l�����v�SX����Y�W���L�BB��O��0�A�eW?����xG��+���ZZ�?�|[�qS�<s1b�.K8-)m�)�\�n{~z&N^��q�wރ>H�F&H�_G����������b����xꭤ�(��d�����{�c�59'Zh��-A�~�,�w�h�{ZɆ���x�D�xc���>!0�y��]rC;%� 7�=wޖC���C������f^�F����Ě�~�,����m������2�r���>��Y&�W�y����9tL�n�*��&`&p�-=���#�hF�\�Q?b���qG��(�D׷o�:_զ}�4b{��FQ@�Ax:6�a��:�4�ߪ��x�qԾ�������[j��G?��_���C5������7�X��p�h��M����_�;�gw�6�&�)�f!?�9���^`�܋���;��YzP�֯�б�6s{�9`�Iq��~�B���Fy>P�dH2��P�F;��$DiVuL|a�V��.A0��%���3��ڻKk�m-�t�ڃ�\�d�ڬ��Q�UeV�OE1o�ɝ��Cݣ�>�����Da,�~��t��tZ�����X!�r�b��?Nӧ�d�ֿ��]	P3�QJ����9����࿆t,;@�;@m� �""wϹ��5����� D�fC�E�dF�'���p��֯�;�ޑ�=D�w��t<����Ӫ94
�3`򨟯Q�.\�����?��ĳ0_�/��8L��T��Im�n��-�f�-�/�d��`@�|�fPwm�D�JaH`y�_lMDA�	(� ^�.����H��团<�ky>�mӋ�	�F1�8"ht�xó�$G{�������^@�5��l=�|ˆ3��$a�]L]��h�G����~�DM��:�A���w��� ��W��A͞�HWe���#��F��M]$T�����bZ\�.$�8�/4�)�5����,��©����$�*��pkVS8"*���5�q<�UY��4QQ"A֛d�ϡ\�Ң�&R{}F	+���}�^���)f�=MCQ^�(�|@DCS`^�C�FĤ�~�b}&���,}]�z]#�ſm�\�1� D5�5\�-���'����N�B��+=�\ϼ�/��.�Tֆ.��֛�݉k��v\1!�����E)�/���}�DB�6��_0~���N�xȔ8��m"�/z�~�=���(G�l�d�*q2�R��v4��!��ٚ���ϯ�?����ӱ�ؖ�I�����5���OY͎D�{:��Z���0����R"��� `�{��ZU<�K6���Ț�ѩ�ց�I1���_�K��#RR*`�a�,��!+_��Wy>����UN�9�	��{%ki�F4�ipԫ�&ه��3؟|a���Pq8�����%y�'��a$K����E�J!ea�F�1�-#������Ʉ��GX�c>����QX+���@L�7aԦ�'c���@Hx�䮵���vw"\n��K/A��G`�y�)R�ē��[N��ò;�T���f��ЈZ� �=)��`�/h�V�?z��F&�u��m7�z�:��fX�i��ݣB�EJ�7ལ�Af����b�����$��r��2��Db2 ���Q�&F���DM��!%�|���
?z���S��	�Ao	��������x�y�	9E$-���7o�⃭u��:�׳����:[�t����ǣ���c�Y��F+�pS���[��Ca��"�M�r�V#8��r��'�?�+:3 ��t2S�sY��[����q�iG�So�����全
��R��9�yu�H�*$�v^{ ������1t����#V!����+�|��=��{��aL� ׎����g{���&ڠ	�����z?`ء7Zڥ/�J�a�W�8�;<�[��A�&����~�[j�;����?���F�k��:�#-c�������@̴ao�(g]����� g۫ԏ}�֨{�}z�U��Â�Erє��mFV���Xii���Da��+�?�D �����f�(St1[!��O����$�;����� evљI&Fu��LȂ-��$(���|6��I��ʔ�m����C����������Y]H��n�.�<J�����?>Mz�=��T��Ӕ�vU6x�AH��xD-�S@�YL]|��*y�?p~�
���p��p���}��Iuj�(b�Ծj/i<�л��924�Ԛ�+f�do��$��1pda0��փ~&�]~�X4�������(��H�J�sv:��EbP��s��/�D
K,�q�@q��D�sPÝcn��	)�ީ�7�\�|��q�+T'����|ھ�7A�:�T%�>!�4x=$��4���X�R��걌O=�ۧW�hw�5�}�qz��'Ĭ�~G>Y�R�����)�܄C�D���+2N��R@"ьE}�~"�c�(�s��C?��?w�VXlTHU]�p�9��4�V`HNkvW����:D�Շ�ϕs{��!.8LH tB���ُ�Y����m�/I�zO�M$u���x�T_�D��SUOM|�srI �-D>tr��l�\��ؒ���Y
���1��}�(���!
߿���4�Щ���3���~��U@�[�>OMfu�W�!��Ŷ:ݭ�Ht?H�,� #`�#5�?Qhi;>�lZ�!ؗ=�����j��G�&F�vs/-?�?�Ń�~i6=5�`]�#��OF�"�u�]7���\�k3s��E
��(��6�����4a��횇v8���s�������O7�tt�MB<��_NpZEJ����sI�L��� '�Pmw�ԎU��euS��>��Nr_WEV+<:�&B��t�R���H9�3�'�-B?gS��ʫ�Q-%��4����(����u5�`K�?����)`�O��jЂ�@�|�RE�����z!��{"��)������#�:�h�.����ʐ�����Â*���#��g<[���h=�^�"W��WV	�d���*�n��AA�;�6�6m�a�6�x$A��IWz�&��1���;K�m]-�I��ȖC�Ṁk��$��k�v]8�1�!�ܔ`J]�؛E�/'B@I&���ܚD�H�hz�>�6�c���4��O�YxUY�ChtȎ9��6�Ei�Z��J|-^���w�Ǟ)�z�L(�8Rr� �P�&��t�h��$!<��^����`z���pY��$ :k�P�����Xy1�-S^Ò��R�������|�)oV���Yv�qH��}vC���A-4�$�DZ'Xˎu�%��0��D������6iݢ�P���K��p�H�M��教���Ǿ6L�K��MN�� ��P>qi9>`MK1C_���{���.m����Ϊ��» �A���4t1�K[�R��޳��}�Ј��� 1�4��#�:�O!4 ��\>�9w�:K�dî��V�W��2mS��)�W���b Nyb��{��@�]3�����B�E{ �{��{$U"��ڨ�b[�c��,�^B#�u�� �gW���'i,ø�C�� Nnz`gc�cpF�Vy�p!"�D U:�:����x��P�2L��,c�(�f�@��RD9C�⋤dw堼q�3]�
��p�vH4}�Mvc��`sq'� 5X�+�a����k�{GtӖ��ɡ�'zĸ����U�n����=k��	�5η^F������~����AƦ���;{�ѱCS��23� � BF������K���hZ\I��3�� ����.�"��������;W.L2���1r�c�#{'�(�$�l��R5-��#ւAK�tA%6v};i�
��4/D����7�7�H׍^�"���[&I�*]���G
&q�3��j��4�Σ�6?[��QY�G���Ƶ؉(5��.,��8���R\�"����cK�l�Pp͋0
�sR	�~e��΁�_��_�I,�n[ c8m�	8�qv58&������`�cd.�<�	��:���B�#�W7k�1�ɤ���l��hs�R��(L���C�#L)�F7�S�l��j<G������%&�L�'�=)�^pߑ�Ω�z�h��9tgCO�cM~˨��'rx� Vp�R��~�sp�8<$�c�ǧꍨ�J2t�r���S���{�
w3`{J8��IH@�<0ݞ}բ7(T1$��T_��[��j<�eSh�6�<R7��#5�	�Yu���zFOP,xK?�.���b5�/L9���؋���:�s�,h�Ք��Ny&*�����U�v���3-�����_�/c��jp���M<�&��vz�5ƌ{�E�}�����xy�$D�Vi��H�+<�I��'8bEAB�$��O"K��nd8>k��*�E-�JjyhC�M��7zͶA��n��v4�V<Bz
�
ڮ2��:	�wB���w׸&����c|�-<~n�`6h��E��
l�t��A/#g������j��a�gyK����� ��)��*f�W_�Г,?��<��-��h[A�1kUY����U�:2�zYoz� q�bs0���9(����c�,��e�r���]��6�?>�-hR���]$�݂uWt7������chjx��uf���J�������#f��a�����[�mq<�~�DsҮEY�]S-�	d'���(0�:���t�2@V/�r.=K���$V�
�2��kb|xp��S��d�`���6��T�񥽴bny�Z{W�a9|0����ftg�G��s����qc�J#P1���VZz8�ә���gƜ�f	�I?����#N��=9,a�t�{0��7�v�&��7 ���i�C=�b ��i�=��M�\�]�l}�ji���9U�J���� 6r�mc���{��ys6Ef*a�a�Ӛ�1��Y0���k�����1���g���W�Qq��eM���N����"OAR��u��W��-�T}�m73�~�g����`0��B�V����s| H��l�@�~�j�6��=#������
�E.&j�Y��#�:�Z�WM�=O!���i�7�����(���/��&��;y��WdR�-8�-I[��x'�4��ԋ���]�Np̬@�TLH�6%�������θ�-�5��La�&?Wz�����0�T���6$��%�P���b�� M�	���n�_*b��/��
�)���B�����e%���@<�]�q2�}����M������ 9�/�w"���ܩI$b� A�7���f�.	���"���Q�5���Ż/�#.��5�n��@'Y��I��P�{cK��G1��Dd�o�݅��%�8���֟|�N�����Ŵ�IZ�#�2Gjs��%�>�H�Y��:�i�	DY�
��^3 �D3]DD���ch�"��@���^X����T�����n���T}�s���=uzM�!M�t<�]`x~�s�^,�,p�KCB��.�_�h�`W_�A��z@���>�r����.��oЮT]%1�6�X�0�[B��۵�"Ǿe`'���[`�1gO�i�Zk1*��q���?`��sxU^T� D���C�G@ͽj��d\�2U��N�$d�,
��$jVi9���˘o[^�u�o�T.�"� �X �TGkwC�t���d�����3���(�[f��g_h�	��F��Rѷ�>��B"|��?�6�[�k?�A��|'W�АJ?� -��cF�L�Į�]�����1�?���q1�/�x���d�3�V+E�����5���M z��g|ql�)>&�MF?X�?W�W�eS~��6��B���ruf;4h��h�R�z��˘�ȭ��gfN���K)�QS*��$![�9mnGG |H�J��
i�^`g1�\�=��L>��6���+��p*_Cj�c��x̟s}�A�ZPT�,͌-��jY�G�czs+�D�%mz�3Q!�hj�#��S��B��t.@2���7S�뱆��Ԗ&���Ifb��iԐa7���0Q͵_\)䇖_Y��M�R\�3�e��rDۂ�}��8{�Xf��OB)�æ̎oY)�~�;�\�	�<��z L�g�n��?�q_xItcK�Lt�oG����Y��� �Z��N+���2�졣��4��+�Kb�?
��eY��\Y1lA���	�9��֋�ggȽCE���}�ʷ�]p� E��TcC$��b��F�M�Msіg�R�rC�DP��R�G�E��P�n��G
�GC6�rL�ه6@'�����8���㢡z{U q��9�a���y�g���O'��0 �P3�gGUգW�$EZ�>�g�:3�����Q!l j�.9^� ��=�Ќ� +v�u��k�[�f$��\Y��J��o���'�b��T���߶ܦ�:H����[$b9GӜ��%���T��3R0��?�.�wC�l���=z*=�J@fi�p�� Kj�3!��-%����k#TR�́k��嗿s�lF�B������>5g`́vлK4YHl&��VN#­�
��,��͢>_�2�$�����!�?���'�6�Q�C�Nl��A�J3{'�p��$�fg&�_��~�Gn羷�Cۿ��E.q�>�<O�b�TE6�O�&5�c
�qWe���3ۜ���b�(�HfS�Aɠn6�6<��Y}V��������ʡK<EU���-�Ru��eW�
Q{�R��C�qb�n0��;t�Yߜ5w���bY��k��'l|�o��WN�7k&a��3q{`� �n4O�ͺ�
2Ƞ�D�%ҫ+!�z������란�1�:iX���F�F�a&����m �>�%���[?�|����1������kY�]�KHl�>S��SYۿ�6�QY�w���$[tK_G�*���A����o�0��N���h���o�<?j[(L����I!��e��C�CO���l�C�X�g�C(�br�C	b-���}�[M���s�!9dg�K�	oE���z��d���q-s��Vd{�9�=h|�d��lpbʠF�l�z���ɡ�taɟ��R+� L��Up =]B��W���LKj҈�����(:i�ˣ���4Pf_�U��"}.���ϐ��W⡖�)]< Q�/�F�@��yG�	�¶���G�R� �0%�:+N�Z�kQ2�p��	~�ó)�o�����R���P�>S��tc}3�;�zMq�G|�mG+��i\K���˵����]@u�	�y[�Gw~(u�f8�j���%#�)t�c�R��/�5/C�O�r���b����K.m�3�b���!�/�7��ɉ�U�i�죘��N�G��Bt�c�-	q���.��ˁ��	O����` �g�I�����sB��7\�S��Ծ�����DL�\f�ޑ�f�怑�%M�w�"}��$8�i`#��]^E��וf�@�p�;PC�M�����ı��Hr�@,v
:�'�DђU�1+���ML��?V��!���\��;����Ke���Ձ)����;��`��l�G��yh�`�\��=���㫽1��.�/:2 �[[�^�cQ��Z���
��%3��
�A�ӥ�g��ۡ�ߡ\I���=zV�A�h��BZ6$DX����>`gtU�	v*�T�����6^q���ۄ?�2�V�F�;����S��j�A_�eOl�0g~v�6�F ryq�'���D�']j��eV�7�2|�� TAH���=M�����P�����&~��e6��Z�'��&�y�b3��>�9j�]KF7��f��g��^w��k<t]��6�*Y��N�!w��9nI��բsˍ�@����c���6���N�m�|�^]�
��I�p�k�p
��Sȣw����$�>Md����)�w����`f��/�c-�i*�˕�JANǕU��2�z�oQ�S����2�.�-wf1yV�8�%���Y���k�he/O"5 � h*,�y$�t,�Yb3��,�G�E��Y��k(AN��B�����������ݘ�-��}	�Gy���f��}4�ô,�3b���>-���t��9M,I�r|\R4��-`ؽf�ƃP�w=�,%X qq�ڸtK^,%���i�tV/[X�b��w�ܥӖ���͎r��73ƅ�:���	�c
���*�����������[$[���(���)A��	iU#�u�xJ���������d���p���I�9��>g� Fp��K�J]^� 3.$�Kw�$����;�֯U�����X�c$��Nz�����|K���`j�s���U����F�ѿ+�g�SzQɠ���0ӕ�O؍���lN�9I��mOג�J�"��5�����8[�~$���,�6{l
�yNM�5":��4�k?��L��� Q���6p٪T����R��t�	�Z��Y���
S��%�ތ]���������փo�Y�Q_m6��/�7� 
�d���~٬�{���O9�؛�j�l�����ڳ�EC��t%!g���P�	�C�4� ���J*Ш�%�S�wg��u����0�P�>]�D;����re�x�$<B�>��.�<�����������.8�</2K�GXt���;{�27"��^��fء>�L������?��~z�^�b"���Y|�Q���`$��&�e�I����!
�JXZ�k2%i0���hD�'����v������ha|�}[�e��
�A��y�Z�&�	�73�|�+�N�~z ��C=����U�[�<g����� {�?���W�:�������.=�M��k�42���~w�w�">L�1�9�J5�7Ţ�y����x��u�Q����#��!џ99��Z(�j�V�C���5�;`(��O�ZW�;e�U$Լ���ٺ���^��J{0ϙ��5���~�d%�uHF�P�2�g�����[�XkH��?evz�d2
oȪb���D��TZw�#p����Z�f�T�d0��,݉��}����\\ܭ<,���7���j� ��$�Ud�(�^�9�=�J��i�;̺�>8���s�������=�)ɵg���6���o��Qp�`ѥ�I�m�An����_8y�X�#W�����uN����������!���lʣ�6����<B��
�۲Aod�74�0��+D�]J	#��a�_���@)Xy�'�k)����B��oBh���0�$V��[b���7�̳�����}s��e.���qwF������B����ȍh���l��m��7-s� ����v�]���_��:�gEǇ�S�S�I�.U��y� �N�����}��:�����W�9J���L�w�Wf)IJ�� d���fȉ�v`M�&�,�������G�C��S��Yj�=J�B��4�m<�20|4!m^ ������'��y�ݔ�}h�a�ȭ�Q����u=��"�l�U�T{,��#��s9B�<�J��lb�7,�o<v���W��w4�kޘ�?�!��8��#�S�V��;��y����1"��>7��v�،m����E��Z7� )�փ����Sb���;����+�Z�yf�	�L�2��Ecf
E�(����LΪq#�Xk[d���.����o��F�y��'-�o�V�&W�z�����2����^|�6@���O���L����"�5kN��j����`�q��o�[�Ǻ9�8��'��v�~*�Y��f���U`I�4��Їu;��z�����`�5~���G�F#�Q��EJ�V�膲�Y��4O���CIQ<���o@e�~��^!\�ǩ���)���r�3����v�&ɛ¡zJ��-á���h�<��ǻ6�G��u�`'�Ny����~�ղ�a�}a���pΆ:�����q��S:����C]9������}/��%�<1��tS�'3����4��I���[% G��M�����[ϲ���;�1�p�Ծo��޶��@C(��-�F�Ү(f���>!^�9Շ�_��RY���v�2^G\���\�G[D�h�å��Z��6�,I��T�l�|0�f����	�ȮA�p���w�
	-��\!��kGjk��ϖ���Gw���J���1�e��[� Z�+�IV0���'��s�j���B[�A|����]iȥ��"Cٲ�����q�4϶D❄�dţ[�r��T�Zp�*��rin�C��m���?N�h��h�q��?���:w�I�J~�q~��&a,��P�p���[�IN*�I���+Ƭ�a*Ա�� ��n�Q=�.V�ͭ���Yr�hU-�x��rS!�˻f����ҋbv�~���+Q��D}�l;�;ُdɼ�׎r��b��+ѳ��l�Mv��D�^;7���C������I,�:}������+��F���l���B�����H��ը�7���ȴ�^���ͱ\ԕ������=@���(J�՟�L��gώ�fs��#��[��T�!LńGJvґV'=�N�P����<ER&G(к�A!L�x�z�7ʙ4`�I	K��>������`rU�v��������f����ܪ�M~f�"fal��D��L��D�ύr�R����'p�@�AM~D����0�b@�=H0Ļ���/�!��1��:�Kd"A��)�~?����y�\���7^�b�d�~���ʚ��F.�A��W��;�	rH��y�{W㬖��Г�X��迍�
�W8��Ō�6���R	��=����B��vvz,@mX�^F��cqVM��V����&;v0$v"���G�s6in��u�R1��Ϝ�"jg2GQ���;�B����0�3�H�l��!�P.�r���\�)\I$�rB�ѪMG������|�N������t�)L�wi�@�"�P<�l�ٛ=막p����8F�(%B��β9���<M8!��;��ͱ�*-����X/��%l�q^
i%1qr��T�����>CɞJ��xO��C�=kBQ�v"i�b�Ƒ��@a%
��Cɓ \
	�r���ƹV��=�3��4x���[��)�q��$�q�ª%�s�1��R�h�M@���:������v���~u�\���?u��ŀ[@7�!7Jl��o�K���RY�*GI��}�^�}V���PSɸI�]c|�D�'n����n7�9!�Qe���>�e�/��^`����˱��"ט���/�r����I�Oɪ�X�T�۔:���t]B�4~%s�a be�"y5�z���C��o�1A.�\ą]Q�ux4�3*�������$ChmTjE&82��ä���[�X�ϔ2��I<��kɁ�E�vn��Ҁ@���h_�ӹJ��
����m�A�\����mT�{g��h�=t�����,���O�sQs�r�yX�eO? � `�dp*��Y ����^'�JiN�&�HF`��-�R|`B�O��<R�S�R�3��E=�^�p���I8g;��6Ѐs���3.'6k��Pb�3(�K5]�2�+�a��T��q�P�hVv�~�@�Im�9I���q�S��L��=��³�D�x���Y�8�0�"�`�v`'��2�\%S���,�{�9�7�a��Y�~�/n	���,�/~<<?)�oڿ:����龦j6KCpmCM�s��v�x��{���W�ů�8K�����>��d�8�;/6ƭ�10�F$H<� -SQ�pI^���c%$[��Lu�P���I3�a�~A�d�]���`�0Z[�%'�TNaL4��
	P�YP������E�TU�c��;w���t�/
#;�p1�{��t���o�����P�� y$��h�սe+DB���1�%]�z�C�"�&�#�8�^�F����tZ��F[ހ<�g�a�R�xX�"�7U
LH�PJh����W�1�\�����_�r�/���C��/k"�8��X�wO�(���E]`��YYO��3�6�	 [E���\{^�v��ɚ����d6�#\nbM���'C:�S!����5��A�M��s_�heI��a�(j������HN�V�1�ǡ�r�i~8�q�_{"9�Xb]�v���&���c�Kw�ϩ
	��I���J���}F~1;���r��r����	(�п��9OO��s�"6D��D�<e\�lO
�|:��6B��rXmvK6-�����"�Q]⬭���eqQ��m���//W�m���W�Ɋ�֞	�	������?.}��.�LQ��L�n�1I�T�\����ϧ	M�R
s��iV[�S�2��{��@Uh�|	¸���OB}|bx���}"��OU��t����'�m�@Sy�'Q	�p~��M�85��w���-/0`���K��W�s��0@����z�գ�Ǆ,�a��.�� hG1 e�N{�	�
�C1`}6��C�~��zGsI>&R	�QTt��&h���M֙Y�72� K�U�v�
&&�a�c��C��춟�}d]�8d���N>E	��5I�
1�v�wA-�,I�f�%p�}�nl�a_�'�x�VjR�y���T+G8V�uA���K1}�~�,�s,S���ЧX ȇ���3 r��
�(�CF�2c�b˟��RG���Bh«�3�}ma���V���Պ#A�5$����(L�������n 9�QK�k�<�A-�c%�?��_���6�ع3���#o�������I�/�mr��+�+��R��ɴ�p�[���:��$ZV��C�*�|�2��
����A�S�VA{��'3����e'G�� D�O/����U2�<*rLHh��]���#�"0!ގ:��T���6����S�L �����_�߃y�' &��R�>�֥�D�����f"K��n!�_��j ������産�[ ��#\��	�4tA �R�"(Ο�6iB"�$3¦[anꝰ���po)�'�$;>��r�k7иi�J��{ǟ}�-⬛a�-b�Г��8 %N�¥��¤�6&����	TWС�[���,W}.K�Q܅�|N�R\ƽUĵ��6��v�1�,����k-�3(��W��t�����w}�'��:�>ɉ�[�|�5���j��E������)׶�e?+b�=�1%�(T�_No�l����Q�<�C�t���k�kb^�BjW����L�֬�I�H��؂e�v2�����c.�5���p��J��@p��Njw� ;�*����5 (A�ś~��x���M��'L�{�ƩwL"?d	�q�h�29 1s�PP��W>.ي�#�JGU�-*���g%�'Z�BX�ţ;X�%��F9P�Nj�H���`]�"��C�U��qw�W�me�_i�d�Sw��:�"H0+id���|�R�eD��N-I'����\
�Q��9�J. "�T�+Ŝ��x�����;z'�p��Q�G���ʓ�Fr��C��#�����J*�s*ڍ�Z������&j�%K�+�j�ϭ�כ�5C�P�s�}�$�i��:�ؓ�����f�!���
�g��`������2���@��X�a�\e�6�k{t	�0�p'6��}2��ʘ��j��9M �'���h�XBq�zX�U|�xZe��\e6e���AoIwJ5�c0��YYFր�����YǷ�Lܩ�ڵ�����̎�RY[R7M�;�W��L:x�R7�Q'q[�"����׊F��S�%-�-�\>��8��׍\����l��	C�x�H>���F��6�o��4}PoE�Q�/{-��3q��s��<M�ȖҷQ����]!"��gO�E��C:�՝UN�>)x4�y���#�{A�֝��>&Bɭs9F���]i�����J:BVM�d�ۿO4����5m[RpQ�ț4��x�{F��⦙�bkp���h�@9yS3��DrRΐ����Q�������(��R�X�^_�R�q���("���`l��� f���'g�������O1�m�
:0��8�P�%G��mWH���I��2,�FSqr���!(N�}$� ��|�)K�5ǁ�@y�V��"�$ډ��Ԣf�ٕ��b��GZ
>��b���L�����CD�P}K!A�����zV�y9�`��%#3����Ys
�n�Uծ��͋nX�FZ!��x����s*��p��ɮ~Yc�f�P�גk$���
�T�j�V�1�8n�g�v#����<?��Kӗ��#�R~^���<��� ����_������+���X�� J}��j$���*�߆�L��%�����6fk�i�nA ��1q9��/P�,� ��4ٛ��*�"a����	1ﮜ�'�� �2�F�q��ë�bg7�C<�.�â��^��&\X9�dN�%'{��� �"[Y��9�[��#�# ���B�t�Ԯ�,�eK/`"�%�oa���;JR\ԕq�<䴕	:5��y0z0>�C.�~����f��a�C�4�J<���?,�	�TidW��n~��6�>�s�a�A)�0��F�19���6/�����b��{nqAq�����A���1��g���5����`��s'�k`�U5���nh&�O�ݮ���R3��3�;�P���������G���$��,����^��9�'6X�x9^�o&�#��#Z����t��.'���2���٠�n�E-�Lge�d�9[x?y{��_�'@[y,z	�C�&K/�A�$Q=z��`���6"�;mӎ
�Dt@Ce�&�����-ūXU����:ܩ�J���M魺���N:L(��������B5jm�?�'����@���"�?���,�/�3�&��)R��ٛ�_��=R�s���3ʀ� �bֽ�&e�ae(G&�C��yKLo���E�(6<�\`B����C5)oL��@+���ɤ�j����4���/I�we�l�2{v���c��n�a�	 �7���E�'�§�6�$x�d�C�h%?���J��e"Јt|TD���K�
�&�5���C%J�����[�ԥ
P������΅D	"THЬ\KO�=�\ok���g����*Ng����L	?�F�ۢ��R��><Ҏ)&=?�� ��-6���xi��O��[j�M
����7Yv����gj��k$5�_)~Ϛލ��}\����f5&7(J���Rjĥ��R���$��䀄��F�� �S#�Y�L\P�n£af�����C���:@���p�G��`.}qٲӻ�Go��C��|�>�9��c
2�IF�{�b�`z��s���,�	�+E�,��vZ�$#��WzQ(���/�IXH�pI�b���,�[��rG_N�?��h�k�ŀ���2�h�s��'��l�oT��]߬Y`�{Y�|o��8�G�}>ve)�
vS�NKO��F���뺓EA�嚈1cJ�����䞲j%��8Cڵ'|I4��Ʒ�k��*��>ZA�U<�m�P�Rry��Z��R��1�Vj�^!��T� ��$/��M�I���a@D=u]v�V���8���C��7�N�e�V�b@�V0�Ӷg���T�U��������Fu|h4�	zg!;𫡲��������kb/������q�SE��,3KZ�´|vr�o�����;~��R�>f�w�B�o�>ꇷc�Ivs	jA�FBS+�1V�ZҊZC#g��.e�4�ˎ�^޳%�ۘ��^�Xܢ9�G~��q��d��xYg�f�i�n:g��x@���3�D@��Qv��O��g�o	��b ���G�p�(�?Z�"�_�vT�#�
�W(�*���Ybnˀ:���f�Ҟzc��S,���CT8��� �=-m޵�ra�`�] a�3�kU~��A6V�KHv�w�����E�9�5Ys�v Y���N:7K��ZG�/�F�
1���F4��~�ͨ1b0���H@�N�Fd�N�����RC`"gdC�=^���y�Q<�I5T�5�~W�".�>�T��/1�a�z�M՝��B�rP+���B�5 ��5o#"(�WD<d��Neg\�4*�9���b� �:r{����8��Y��Zx4���&wĐ�����4z�FaǏ)K�v�*�*��_�_p�mCE�����$����C�Mp����TƄ,�1��̨&!Nxi��U��R�#��鳅R}������>6��2�
�ߧ+	��	SB�A�Ps_����b��z��~|~�q�Z��uY�y��I�b?jq�����d������S��B�@�&@�~�ҳ���t�=vб�e�
_�ׯ�}�5d��L����*&`c���@�z[�7����kSL�Gm�-c����{�J�~ι��X	��
 ��6N�n)��H��leШ�������ͷB�<92T�|��gSxE}�(�i�2̼Y[1/�>��Lr�P4�~|������~%�u\���D.)q��h�疪�ϔH�#�v�I\��ѥ�<��0WAe�X�m'��Y�w{/�n�3��˸��4^%���őN�G6@�|�}8"�E�
����,���������-V؂=5Wl9?J�8\�]7�n@��F�������t��}#[|�Q��ia����F�&R�ˠ��ꌫKt��<�n%�C�p�<��N��{0��2���s��@�b4�WB?�3ïٶ�(�d;2T�QJ��l�`�uw��'��4�������y y��6\�e 
������5�k�;��KI�:���I�&�K4��+'u`��V>5\S�p�PJ�}`�P/�l����%	�Φ��A�w�5G�W�pu�~��(ё�BL����Z��]�1�������Gt�h🐵�$��G�����g'R�ٜkR�Ԥ���|b/�h;s��T<6�@�*yy��V���[�l�oo��QG �LR"��P�D�ְQ�%��6[��Te������w�C���z���zN�,��
 ��$����۰d��S��X�R�?��G��ʧ�+2�%�}�۰��>������zj�|�� rs��z��f�(�������ӵ&Ƴ���W\�a��*LYUCY�7�F�H��EwW�4܈Cx�z���;9����}�5�N� �6:7�����O(;��!��IN�X]*�����I�������V�^@�4����(�~jN���o�A5���C�@�좬VWQ|Ȓ)m��镨b�ҙ�۱`!��o	�
��j�B���N=n4�m��\8yl����M�~ ���jM:ő�k�����p�B/���ܮ�*$2�ͭ�d�1υ4K�S^��EG�T�٭B}D�y�2�=��p��+���<S�5�Ӝ���aac�=�F��:}�!�����G�AD��+v
1ֿ����~O� l�9�艴-;|㞬_w����~w��J���j���jP�tn��7k�I���AD���x0���k�ރT�9�PSܿ�8�����DU�����a$�i`�KK�V<���?"E��� �q��XW%Sp(�1A�8\ϔ|��i�^���y�s%���]\�e�?�L\�@������G��B�h,��$E������^P�7J�1Z��g�n>�
csP;6��m���$+�Iㄟ|�'��[�93�X���k�6Ì%������Ւ����Q��ˠy\GJD�ϑ���������}�����2����	r=;cKҺ���;����������ڔ
�W��47���g�S8du���$��/��{�g��m	 ��J���&xS��od8/��nfK�8��� ���q��K�@��|e��D/_����!�O�N��و�4�_��vTS��|J$νy�q4�8A��a�8��s:dd�E��;�c��0_:��^�1t�'�CG�����\��\jw�qB�x�H�5���r��5��BgL)W�M�����i_�m�G3t�D�e9�:�� Io��cL$6��OZ_�;�|mx7<㓔�<:����k������df)�@v����'�.� �˶p>n�c��hϸ�ln���=:����RN~Uwo�w�=|_��X��P���}��૞��a1�͓�>�m���*[������I�/w;�|��������&x�o�)ֈn� �/�LI�eb�G�� �?�����RM�<DԱ�UR�?���JI₱�S�9q(i�0�3�#�YO��5��ZAq���( {3N���B=�Y��J�vty�/�B�!`���Zb$��$7����?���*���%*�E�%'[I:|T�o�j�!�;���m������'բ6�[+C�)%vV)�U9��"���XJ>H�n�1 0�J�5ܪ���C(	֌:N{��'�`|�yR=>�Q��i,-�VwO]����A�5�b�3�`�i���/S
��q��	������4����<g����(e�az����S�Җ������N�@"��>x_�7R�1/��/h ���@7ɭܻ���khX�?�馢-(�jB�	 `�S| �=AI��W�T�������Y�z��"v�6�#�7��r�1Y�H��*���'��s���=�F���G�u_h�+��b���:�:!��?�K����u�BO.�w��,�鎈��b/��䫫�l�0�cH�V�3@��ܣǄ�]�N�Y
ڦ1��=c���w��nt����ݸ��n �f��j7jGx��P�P�� ��/�d�֟��	����ǇiQ��Y�i����I��F�;˵��m��I��⯤����\�����5�����H;��7VV{8�#�V���4����&�G�ݧ��l]T�w�.#�^��2�(���և�rH���!o<�y>C�d�T�S�!����T�uʳ���f��iU�N"�S�o{�)Y�*M �)̛I嚓Y0�b�����W�
2 �С��2�GM{0�Ao�7=h)ӳ�M�W_�A�s����J��o�;N�0�����h��u�l�x��}H�@ֻW�*��t��ryԪ\fh�¨�ɼ��T�s����<a��|pj�K�*neb���h]�(����F�M�����v�[�Z�. ߋ��k��^M�o$.9볱�� %��s4.�1���@����hS=�t�?ψ*X��_K=�5}Q����ת}�YR˧���A�D�o�n�d���܎���V=����WV1=�{l9V�Ϳ��R�G�t"]"�͖u�����R��{'
�=&]���ߧ�����K����`{���6��F��0#�*�˙�����C���8�08ԡ�#�z&&��gj+�H^΍�%}�jsc}�mw���Z�U~[L�~)Y!2I�*�\�I���ͮ�J��@]��[���(>�Q,���B��$�@��|=f����1������3n�yצ�� oi����[���y�
�=֐�m�nٿ�'G�y��h���jք�^hOz�9�#Y��x	 ���|�H��� l_�6������V7�^d}X`*mQ0g�_8/�\�k���VW@<�i=:�W��r����XE�c��1c���mm���H�ނ}Y<�)mp��fL�n�Ë)a;LU�Eê�$ٍ�L^t������4Qt~Y��F$m`qq�mN�^L�9�9�z�eB�`ˑfi���HK[:�`u'w��QV�ut�2���9�9��!o4e�݁e�g�����{z3\���כ��W�i7���I;x�`}��W-�IH��&T5P���F,����������_�.-�Io���7]��f�o��6�����^�ݠ�yob�"ǡC]�Xx����]��[6�N���j{[��&���U'��p���������O��w�j?0軸��0�~�܃\�46�� ��[���a����!-��4Jp��TᾑL�AA��/Nt���<u��Ԭ��z�km�WUZ�$ɏ K :��R���߈A����эSfU4��k1�1��O�����V6�"v.�����U�g�!Q}���*C���!"5�x��Y��n���L��
>M�w~Hb�[�'	����^�6X�~��O��7��I}Z��N���L��N�h��_U��O�k��\�p����rw~]�7���*9��Ly�kt8�f?f��g��ǚ���3	������겗�2CT�vv;�s�f�w �([	o�߈���&J�h����������^��q�@��/�嫖*���/�8�a6j�%#�u���x��#s�v��c��aQ�<����R`�EM
�`S�+��f�PϤ���O,�̇^4���xD;��ޖ��N��O���P�đ_cnqӣ��E����rN{�Qh����y<m�+�k�}�fM�dF��\�'���Ԧo�'�30#ˠ��>x�&C�(L��
~mJ+�V�k-�.��x6��dN���=�3[Mr^���������2����^HXl��nV�ǖXo�R̨@	&TJ3_��ԁ��i�2f��w�S��G��;��(��8��&�øﭮ܎�b�P�������׈y���|�"x<�@�y�̯TS:D�Np�R|I��}��٨R��Yn*��&�o�͇)��d��$�� �ٙ��;J"�s���s��0|���V��)l�y��Y=�3�[�R+��k������fb�/f���K�,�]��؏���*pi��@)��r�f����^���v�mat	����^V+�/����a���8\B�L���r�l��(O��cC���ȃ�=0~�NGV���Tc��5+M}���]�>�UFL`	����h�W�'��dR����A(���N��Z�T�+�0�2D��ڳAA�+lpD�=V�@q������o��Utg����WE��[�+7�|eX',O&*�Mn|���f��A1�X[�z+U�2�(�]�W�E�t$[�=)�8>���z�s�T�1�Boq6��b엲�� �4�����s��y�5�����3�i���}�H�)�f��3�IN�cC�)V�۶ L��q�� q9�@��[�%�>�1LoX�Z���@�
(U�� ��� ����1��Z$V�*b���~Ͽ�f'y�9{�����!��ܲ�����#�b�i��@X���mY.���M#�MzhK��뭣�4�����99�ځ�t��b��W�OE�%�����̵&��#ͼ�72_� �E�N�(c���O�s()|.:�U��P+���_ރ�v�S�ٶ!3LI� m�Qp̔I3�7=��A䂪�gi����O�ި�9��D�U�S��G'���e���@w��gk�m�9J.���]+��l����~��Ţ�($�I�r��̳(� ��{f\�af?�ׅ�t`j	k��̠xd!����-�[J�F�~��k�8Y����(�C����KA){����I� ��YM�:�ݮ���9*rg���d���Y�#��(�6��8!0?@�I����M��m�q�a
�7zV%�`ф�Ͱ�`p�@=4��O"٬���
�S��b���/j�?�;�bIL	����s�r�Tۼxe����Ŷ^J�a|C�:�y�I��	7�b����nb����WL��ܤ�m��J�:)5�m*��k,���Ē��J΃��P���%��8�C"���GĢ��Y�j�1�ٰ���LD-��SGz�/�uv1���?���*Ժ����j�I|\e���h0ۻ:x3D����Kb'�� [�o!=Y��n)d��5zs���M�F=?�QQ�_V�`��닜L�0���]``d���l��|ߡ����G:�R|`��g�w�X֥�	�&<����Z�r�M��_ټ��KL����TL�K�e��1�,�0��?>�p���ē"�r/��mn{n�ګ3��|��h 
-��?�e���B��;�R��k�_,P���`�_WE9��K��"��Ċ�VI�g/��R�ף���~� ��k �p""�N1���e���p���i���#����OS"r�/��`���t9�2����-l���8B�8�t��W#�fl#��?�6ڕ�v���a'P���I�^@ޫO��)�k6�bjp<���ftP@�<z�Ò �-)�1���3K�����}m� �5����70RצcO}�������IU�k�%���]�|=7���~�[<�ڈk(��{��U��F��6ĸ�Pu��Ķ�L`_?[k{�;A`����B�b��zw�s��lZ��)�d�-�� ��i�%���_tJ_��fzQ�j��lO7@��b�6�i{)��K^��3�)`��8<�:��sn���acz$�ن.t-�Q(*���'ã�Y<_�M���.s��^'�"�#�TdJT��x��MKy`"�a�9ͼ�ͤ6������k�\$(���˪�t���o��9�"�8��� r�mtU��:�י���N����Z��j��?n�I.d�R�\�hۃ��JOF�CR��ٚ�	�mj2{�q��sr�XYe��0�p�����tj,)>���g��/`fV�u�L3��Q:`6��W�����u\�N�0�ך�d�d��^�6L��W�ϗo�v���Q�B�������|^f�p3�8��F͵M�Bè�SQ���P�Ƣ7'!v���G�P��8�Ik2:?z��$g���5-L�lo<�"FwazS�o��6]dH(s5�f�A�?����b��N�<����<���0?x���N�`B�tTBBID�8��;ΓEo��ʠ(�>�c��Q�j�H{�_%kE!��f.��	"T�Ω�^e�H�U�1��n|߃=�hqz�\���NT��|-6{��E ɩ�M^�m21̳���[�v�k�a�\�%r$Q"H���d1��_�h�y�S!ɿ��:�tU��,b�}�&��q��n>P�t}�{�e�ҹy�5[Z����� ٺ�����ˏ���V�^N�p�ӟ'a�|J��ˏ�j�9��|pzp�v��I�"s��@��{�=ok�r�O���pm\l�$��{�	L����5�k:�cq��$��0L��֩$�(Jc��%��hZ���9G_P6��ő��ƙ6�?���D���d�2��qOc���t��o1a)�1��-����26A�:�BSn�?W�+���n��A���;I���^�?�;R�*#�LS��5���pWdf:��u�O.j��p���E)�y;j�Ժ�IY�§��Dv*��A@Q#�Ά��W7�e)L),h'�+R�<�>� a��JΒ&L+˟�Zxjf��1�d��0�jr�,�n�	��0;�)&�lY!+K���AvR"�Vz�C3��#TkJ=)3ƴ���͟��h?�C�j&qwck�.�1�2�?�Jc��3i|�G�E<j�dN�Eˬ]QK4������'XH{��1:v��]��\j˰��(zϰ��Y�U�hsn�|�u�V����Z� �(s���)���YԶ)��:8�\����O�2�/ Y��h�N�y"p���exj�E��n���y��<k���˸��:0�cYY7ZE�Jy#ş������g�B�y\̔zv๟��=s� �@O����΁c�>���3	��K߷����������Hʐ"�İa;4+$Z�0,���WPe�{34ܸ�U��yB�zdl}�D���^0_#or:& �h����3�6�pz#2��抯D$�x����^3�Mq�f����c�3��-p�D�BWJ]�k���k���q�2T���e<�B\g������t�j�0*�RQ���j�ըC2���WЕ� �
J����VBX$�.
� �r�������^�sQB���HO��A��FrT�SG)�>>��8�pzU@�-A$#f��<S�+\�$OC+�S_�f�ȴ>`s��R�Ň*������vzY�sbü�I7?���ӧ�3h�h�� i3�bzL�9g	�Cs�/*���z-��uZ#��3-9e5ET���y@|E��M����A�)ȝJ��wOɊ��f�Ъ�Ę�C�N�w�ub�IpN	,DJsą\1����$�{��:S�S�����<��/ڍ�:�d�\bRA���3A�0��o#O�!D$exN&&IrW���cIu%����Zg���x\����n�D�ۆC[�þ���9;pK,�H�뤸��7�����8��C���� 2�O��<��&&��A9�4��_����8t���Z���U't.)�-�W0:M�}����'��#|@����:[��	��p��:6ӣN����.D���Sk{������>�\İT��U��� ��R�5����w��J?�w�N�$(�g|��@�؞Be¹9w�-�O�
����*��S@uC?t�4������[I�� � 3[���j��̀56����z7qj�AA]h��Q�A�"�:M���@[7�^�b;�Tp��K)��O������9$ܞ,�� ����#
-�#Q��M��{W�ol�lP��yj f�*����z{���p�}xi: Կ�k������mٛ�r6nj�S��#A(���۶-ö,$G%���`2��`W��Fd\3cJ��i��M��~oA�*�9k����C��~Q���E��C�F��z/�N�����	�O%�,��s���X���dl�x�Ga]���f�@��rdl�B9�E��]�5\{�����[.i{k*�=��BL�b�P(�H�)E�����c�qWsɋ{���Ő���SSn����ד^��ظ!�9��<�
�����2�{)��w�V�]�����M�?A���#PۗE����n�߲��mY��R�]vN�Tx�� ���T��*��R�8��B�W �����:���K��W��{mV=���J<ñ��;̣��{�m:���e'|~�(6����yc�J��|�с����*�,�h����6������>�����d����Z��'�)���֘��5o{ֳ5O�v��d�=(��
lq�#.�I��]�
��%r1�*��.�ɓPS�:�����6b���"%KϱI�}�}�
����qB,��P��Z��jq��'"E�����'U&s`\V�t����o��+����mμo�����/U����.���S���=xB/u�4���f`&�=�9.���V<�}�P5^,^A��e�K��9�$�f[��'ϯ����dqy�~��qՓ����뷬�g9�o>
y�ǂ��d�,�$��vlm��DE��̌\�y	���
_@�g�؋��i��T/t��E�)j��?1W#������t��"�'E���fC/�&-R���_��ªh��߭~Գ�S~� Vy�P� VL4���=�����Zl!m��i~~#��̌Թ�u?�*(a���1�U��5t�s��t(�]�7���=���:e���rƞpIς���|ZF^�����˒�:L��r���)��-��9{I�g}�i�a��(-�NE�!����U���JK�RA�ֶ��bG
�MG7}�~1I=�`*C��Z���^)k�r�L��	ڹϊ#�rQ\��������q��r���X�"C�T?��X�7~����&