��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_��~�og��B-��e�g[���$�Ԃ���#֩�&l��=�̣
����^�����X�#.^�����؜�za���+�rx��TP~��A����v�Z�gs�hyv��"Eb�J/�P�69�-�䑕 ��N��1"�`�����V�v�l>��V]{�2%+�l��s�M�ry.�$�&��P��+��t��V�I�̪�f�,����)&�q�52Q�O!#�׺�Ңe�����B��ڎ��!�����q-��!+lE�(8���t�g��)�]����H�,���<U�)ə�%&���u���S���V"2��A����f7p�n¤=؁(�N�\�x��UY9�4�m����v�/�C=ߣٕ��b�\��e<�B�z�Ksw��-y��I��Mx��mFvRE�`�+��O3~��աU�2�U���gXkDQˡ�`���d��(oܴ(o{��=�8'�N�u���^�:����C�r83�x!��b����ŎqC�?��CZ�jk���)�}K���c�W�|6(N��)�&@#F����͐2v\CM(�K�G�i�C�| �@�烝�z�P����V��8��("�?��0�|�2ynܧ�5���㐙٩�FEApn���l,$������?�F �>�MY�G�����>���q�[{�9˻(�[���hm�'�����T�߸�ɛJs�T�@}�*!x�)� �f����@�Z���{,v�ު�*���F(�r���o�$��i�X�����!���U�r':EHW@��`cS<��>�(kЙ�2	�~��N���p��BzDu��$�x�;�h:��/ni��)j�z6�"��<�I	3���:I5�����&��s��4�@������"
��O��mL�&�k������� l����!��n78���傷@���`J%����B`_ҭB�6@?s����׶���`*<��CzvY��Ja:�9բ9CJ�R�3|���/.[O�����Y9��H.RZ%�^^[��#Bc%����~�¸"�W����8Tai��nT)���fj�q�]׭��<�A��ud��c~23���5U1���6����oI ��;_���iZ	v��q(��T�8+��GR��-Er������е�Pΰi��Ί�]�{
�#,|���6�y3S��dF�ǣ: �h!��2}sD6������2{��BLM�OQ10���=�����m/���O���`{7s�k��%[Q�����y���1��T�6ئ�����n���9��6��� ���`cZ���N+/nr�������:��&V9fA���+���|hb�E1���ad��UҎ-^�k�R��r�k�F����i�n��SDtW�r\L�@`�RR�'�H�p4CdM�'� �M�{��&bc�^�u�P�Jg�(�3�*\��̅܅y-=ž��i�0ix����<���m�^��h�"7ـeEZz��{�~�q�wx�$�+J�l5O�2��ԨOF�f|F�o�z��ɹc��s��<C��<�*֤�!'�w."�bju�c`�<3�?�|�n�&�LH�B�m|綹�P��aȑ��'x M?���&4���,����7�KZ���J�cr�����]n�Fi+Z����}	�1ZԒS(�"����*��cÆ��bc���M�pfrIt}��k��xD��v!��R�&� C��*HH.PóKJ|�^�&�x��	��ʲ�lbD�gj<��ȵm�t�;�G3: Q�t�o�1�'�^�q�9�].K�C�־J5m��������*G�LN�x�|#$����p��@���� �W@����Z��COf�0܆� =�*��޳iߡ��U-׽{p�cЦ��W2�ޕ���e�� E$	�i�����yJ*"������Z0��|Up@Ã�h�����2-���Emm�{ڜ�d����1�10b�֘vG�r�;A��J-W�˔��K��8.���% ��=闳���"3Vܤm�S=��;�^|��xAs$pq���0 |��i}�W�� ���|�(���F<�SK������B�bJ2��2���{��2�����5�E*�:��u����Ɯ��ή�1}�q�TBc���}�S�U}y��r��-u3~_�/6��h�16�J����-�K��0���&M9ِ�7_�!yh4 ���TAϾ���ޭ�3��T�1?��@]� �k��$}@+
K���ku�����v��������oy��i?W���#-4�5�^�._�\�c�>�M���9w@;��X>&�̎gf�n��.+f����:�%��������Bk|l@}ז��i���BV��XlY��8t������ ��a9r��)�$+�ϩj��褨���#˘��������zr��6��y-(�{�I�B1ĺ%�¬"�u<�v������bD9�\��8�y>��}�._*Z��5������
~ɲ3�O����ag=�h�p5��w�.ip|w�4n�DjtQ1[�@/#gģ��w�h�f��t�u� �c��D3ͽK�sk7^j�P��t5D��&�_4
��
����q�l�e1Q��%��@/,Lh��:�˦y3�)V����ߑ��zaW7�R�DR��
�k����/���z\�E�7����y#N����MR���q�E�WK3���ߓY�����AD�v�E��O��D�h��"�P���7�E})�'�׵��k�S�\�<O-���ݒM�3�Kz�y@����${(�3�_}���r���D_s6I
ҍ����`�3R<F�mE�;\�C|������[N������r��$���Ή�6|L PE�Xmn�*��l�G\X�i
�%�+���b'���E����t���!�RY�᭐���P�tO���/2_>Oł
ŭ��N����g^����X�V`�v��|i��a�;M���?������#g��S�t����"W�%,g�QI�{A͔y���){
��wA�Mf�zř��$G���$S�h�f'a�QTZufT-���z�oyvwĽ��^� �+	u��8,=Fӣa��[��+����6��%[:�|:PE'jY#!Q<,(ar�����m��+���c��o+��8�q���0l���0�U6��X��� /Dɩ�ΩX�՘��l���n��|A9IK�� N��J��Ss��l[%�= q(�\4���
/A��=�W���3``?�^���X�:�[ݜΌg�WR�^%��ѱj�����z�\
�MӁ�gۚ�L�3_x�{{$�q{���L #�ʄ�lvq�� ��Ww�?��Hۄ��1:���������]7��_���d���"\;5���)��c#қ�v��7$�e$ģT̚�(ݻD�p�QJB�� YDI�a��H�Y*��qהF��s�.8�<�|)����n����]���|��O�|Wy�w�*4�/���W�<Lm��t>	�U-Mtz��hvH�C'�ӛC��O.�L�&fԳ���vYb�{I-�q� ~N��j�%���`H[n�yl�"�o���6�<��6�_���<x��፶�'�vh��� �k�3P���uك�Z�����1&�y2`�|����x���D�H�9�N4�D��f�@�km+M�a�mò�k�
=n0,��YmMj��Cjr|���xz>`����"L�
i�g$���M���8-V�9nA@�}���q��.�Vb%�%��V�Э4MϚL*��m�$�r�]��֋&�>�	�5�D���m$ )T�!��O�=h��� �2�u��Nf�I��C���T'�B+-�R�ܠG"+�K��*R��ͣ��]�k�:�7�U‪%'
�J����>0Pz���X����~���9.���0ׄ^z{�� s����k� �� ��I�V����K�q�l���bm�V3�9�|09����
9O/���n�ݟ:���mξ\�F�V6��w�>����}�L��e �������d����S4���4�sr����W��z$�}m�U��x{�G�#�!��k��P��.�/�Jr�á�,f�P�f.���G�����zA�N��ح8,�`DRJ���NX&��¥�lUx2D��m*h�ŭ �A�Z��K��!�D�{^�W����Ӿ���`��0�v����2����)����WFU�1�d��1�4�l�)�Oے���,	v�R�)�9b��;�quU��St��x�X��Z����!�r��sq�W�� X�WN$*F��;��3a~vc���q�o,H	�,�<��0Ɩ&;e�)F'���TJ٩��7�� �g��J�l�S*K�+m	/�W+I����4D�2}���7)�F�"&�����T���B��=�ޫ*0�d����e1N�{�5>$���eD4��l� %B\6ߍQUA)x��"��nCC�GJ�G�c��#wKz��#�5��3�u�60��h�劥����bwhJ-ɺ���� I� L�o�YD�x�0�93���M���ӽ�R���&��J�m�/���~�\���>Y4���*�Ǘ�#)~�`�:��P�d2[�|�0�,>�p[���L��oI��䱅LZ��ߌ��@d��ȶ�J�n�籹�U���c�H!���U_�D�reY]�]�5(������TN�"�aZ�e (��n�,EI)�;
$4�ux�	yEqy�!�TM��
M��CȲn]l���>Q�?Ԫ�P����Au̳h5�(��BpSĂ1b�Va� �0�p��z�\�A%�_�:���E�jT�@��]L��b$;.�L�
q���V����q�b-�o�oʖ�A!����0G@� <�>�\�Z�;};�׏�L��n��ZI��lT~�
��k�k�[�5딊�4���Z��Ʉ�6��X�Hh��*��2[��&Y���X��T4�v6��D@1^^�#Sx#��M{R�Z����Ve��YB�wg8��k/����ҙ�O_�_�T�q��<�e:�9H�DpV�ZT�����-�2�Uy�&bA1ȅ����� S����8����`�,�>p�����q�x�ӊ�pie��W����L�:�=���m��ɻ,6R0&���~/���ָԝ�-y6�΢`�!�e�&�	��в�YF���"�y7頎��j���@��B�*��_m^�t��0�Y�Tص����.1�`�!Q����b����+%���b��b}H_?�9�����.h
�*�Q�k�BN�����=��_p@�g�0�'yo+ן�N��;�כY�E��~I�Üa1�|����+C)������@�V����)q�W����}�zm�@V]��<��-��梸������d.C���~5���cV���wm�1�Vr�[�}ho�tr�O�D�o�t�6k���aQ�p�j3����M=h�	���+���{Y܈�[圇�݋u̲����	������R�..`�g�TԎY�k'?������+̶���2y��c�)K\�1�߾��:����R((B���)�g�ʂi|1:�Jz�a�0�����3<�s�����k\J
�[��K|�M8��%x�9_h��~(�\��<�7�����ERXݣ1��&�u�p�MA+J(������\Ա���J7�SHN��8'P�I=��c�x�����N� �m��Μc�&���`w(�C\���[��_�F�[�S0���X�$����4���Swm���5�	|A�wv��`���1>�^��4���7�v�X=hdb��A�ަ8P�� �F�X2���h�ZJ��@� |�J'V�bO�B���׭�Ӓ)��ƈ�����b�9���]�Wl�yx[)��u ��v��$?'��]��� =����*�or��/��'5'#tE Z�q�I�q�I�\u5܀6Uۤv�UhM����y
Tv9Q���z��I�����b��sT�RC���ṧR�1m�*prWP�'4��ȌvԂ�Jv}Ǽ5��"od6�RƮu=��׌�jb,�u���n��3>@e���ꯤPL�b�&�e��@SvK�ꀿ	S��vL�C*�(�B�G���l�� ��k֫w��r�kY���lfl5�?�Sΰ�l��4Lp�3���rx_"��(�e-��7-
������j�:���s��i��>atP��@3�s�����2]��E7���[�^Rzבy����Яn+_|���7��e^�� �c�Oef�sys'uL���
�/��Z>��h`f0�ܬ~����N��8?\��Qxn�%4�	�/7�2�� >���(��~����$�"�"4U��0=�j���Ƨ��`����6�L���d�d�)�B��hw=�%i}�����`���fs.BbB��v2�jp|^�$ $#�1K�Nݱ��{d�c䨠ؐ3��0(!&\L��o��u%R*K���z�
��z=�x�n�֗ܪ��!#�IPϵ�e��/F��y���,kGodi^v�*~i�5����5uJO.�D0��֘�ޘEw��&�S���u	]���׋<�:t�'E��ޣ8��-fPp:❥�
&<G���<��0�eO��x�Yw^ͪ����-��H���:.{�|��	H#��,U>XI.�]l�<Idq�z =�| �y�S����<����\�;��hs5�ߝՙĿ���m��Ɖ�
��[������$ `W�+����8�h��t�J�
M����U\~���-�v�琢��X�v��޷a_�|T`L�[{�_?��Հ�P�P�gē�2���>W���YT7bZ �i.F��w��=��U��-k8q�|L�ct3�W#���yq��L6��jh�kٟ�g'�Cua��,Bj1���E�O�O
��7�ޑq�svY�C�ت�Lz�b�H�6��<Œ����L���>C,�F'�N)uD+#L��-�o>tĤІ��Y��fS�+�DX��E�94=h��w�9L��>�k�$��n�P�zX��׺Q.���G3�;'�YS��N;�(�H
�%w��e�����/�������9 [�F�c�B�:��KY�-�|l���%���O���`	A5j<�t�������5�S�8IyI���'��L�ئ���`s��蟟�ޒ:�1wᩬ
�k�n����RI�F�5����zC���x������{�&����$��բsz	�` f�`
hQC��E'��X%�f�ʸ*��w��9�.Qj�G�����|�Vb��J4�pwH
}����  5R�ô�~�q��l��x�i��9��������fV�x"H1�k�)qK�>�:�n�v���)C���6��E��a^��])ٔ�O�r#�G�e���,`�G�p��IH!����*G>��A8>��_�M%$mØ'O>4�\�q���@�&�!�e����r� (k�����ѵURJ�Q�#qÅj�*��9�.i�Ы��u<��6�}���.�Ql*�b��@�J����+���btt�du�2�+�nڐ��f�L0�E&��~�3a7�̙+�Ѐ�=��7���-������t޽�	
ܟ�IE�/��`��U�Z�B/�����I^a$����9$}N{�yL����E��ekթtzU'�T���|MK�k7,7t���|)rlM�t�/��GQ����w�.3�<��޿UVn�'���9w�F䅠r$-6?R����$���N��o7��⤧��Ļ�	7C�oxԫy\��ӕr"��i�W]"}�D�_/P5�NY��q�,�e���8�)?W/��;G�]�I~�8��	����[����LC%�T|ہ�D�e��Oȑf�'L�#��Rg���8ˎ�����(��p2�~D��8g݁7+�\��,+?Ǹ�B̕O5 ��˻������O4���%]h�-,gΞ7��*K�N�4Ll]�(�v�e��������M��]���dt,nb����_,��:�@\Ŵ;P#�
[U}�kf��)YÕ���
��|�M]t\+�x��d��+�q(����%�1�j.��fRl�T�*%AL�>�Y�x�K��8����"g�K��@x��WƆLX[+����`�Z�_���Y{p���:�j��֨��|K_��H�Z��5�Zז[����T1g;�$�F�j��8_	�SFM�XƋ�+�\Ѳ���g�8�����;۷Z�|���h3��TV�H���}��zz�@�Ɨ&�į�5����}�<�똰Z�~�{�@�ثW6b�tg\�P�x��6�&s��d$�Y����3#� �����s,JQ�;���#1����<;�-��[ƞ|5��X��9:#��	D�#*:���#�H/a��F�e�x���vT�`��g�8˷C�����g�_Hf3��]جo��W���)R8��O.YõS�,�Y�?1���1��&u�|؝�nct�5���#[m�@��!�(G��@�k�X"$|N���'/Ӡ�u|���Ls2�"�h9���~#(�y!,��2��Z\��B�TM"�K�A�����1���J�+]�H��j~;Qgߴ��o+%XoM ��_fI.C�H\��y�;4ɝ2�S��M� ��jH��N/d����y��ۤ�t2מ=��NUT
��>���4{N�m���_ �.ԉU�q�����f����Fp�����k�L��r�L�m��r�� Gֱ#��t��=80j,X��h��5T�*�s�*E���11up1B{��t�����+�0�"��6���_��~��xE�����
�O�/��&��.�����ߒ���+V������Q&0�.�8P�d�$���Y�n����c��,ƪ"���������9��џ�p�	���H�9��YV*�Ҧٞ��e�ĳn�S�9���h?���Ǵ����L� �O�rg���X�+=��OT����)Q���%��i�{CL7="t������������ߍ��6�5j���m��M����(:�ti�T d���sʧ�����|�^����E�LC�C�]]j��p ���wB�nƬYI��e&ծ�q�*�R>�e�EQ|�pb��8Uo��IdN��m��H��t�ϱ��}�u9�6��Q�x/b�Κ=d�P�ñ�N����W�A�pWdrf�� �JX]�lȨ�*���M��l�%�ȧ�Y��pmJ�5r���2��j;N��=�pk_�'�R��Z�����_?���v�Є^�m���V�OI���J�
Ba����<��d?����O�iR�P慡]��TєuW�r��ݿ�3Q	T��J�KE� #3�dX�ȫ%Xt��ٙ��#��;���b�`JP ��0{�j��?��{�9U����W�դ}͒1.a
j��g�a��,�Il�Hw�f-����~�[�[!���ä
�4ONK��vxD��x�J�t[� ���|�2M�u ��G���F���K�OׁCeG��������=�h�X��L^
%l:�ԻI���i��ʝE��#�i�i�ϗ~W��� �X#���-�B���i�����-߉C4	�x�^��o���F�����K8����Av�3���5�6rNmѢg�/�{B��z����)�`��Z�jl��@@3֒�
3��L�E�7trc>mC���}#����J?�G�b�=����YXG,F����6�T�}�$�����ꛚ��"4��92��{%?~Ѵ[�����c�{����E��y���{��P�kD�=+r�;W�a��yQ�J��l��ϯ	o+���*��F$hZ��R0H�g�@�#�DQ汥@�j�9�y,�KY�!g�{{�����0������>��\���i�g�	�Z%A-&88���i?R���1
,Ϝ����}}�.���F.���iztq�>k��%���ֺV枦�� �>���gU�U��C�B���Cwnշ ��>7E�\���#P�<��	g!�x����n4���dt��F�Iss�~$2_}�_���[�]["���a�k͙M��"����f;P�J���U�2b�R'�1�ǃ(5��t���9/����Fx�A�{�3^�9��#���Ԇ�ܷ��	��~7�%���90���AX>�k sW����y�@}�ٽeW������_a�W6ܔA�Ś!ĳ�ɉ�M�5���n�3'���62Wi�e�yO�����}z�)��6��C�$�edp��΂`ߝV��f�����'�[7�w�G�xy���>k��������]�'�.�$7s;��=�<�oL(ѣ/�q���f��FXm�:hm]��{+飖]���]�	�?��zPZ�D���@趍� R|�O0�Z�ԇ����F��7��dDޞl�i��N���pB+��u;����p����X�	%_�B��<Y�(�.C���{���=BI`�9�nV�W�=��}59y��-x������rvZ��P�5��Q�P�B����ϕz�";�As`�I����M)�LDsɈ�
F�pK,k�9�Q[��������.�Z�G�I����D�
t�˕�a��J�Q`��]��X9V0��I�+�"�^�r.�~P�p�N3�ٸ��g�T�-0�h����x@����s~��v���<�܏�a�1n��9�t}���鰞X��/������.n�z�Ǜ��08��\(��_,E[��|���ٌDI��{H�:��e f4z��L�˚!���F��4Û��c�1��P��u����Y!~,�A��_/����E/��iU�r����J��(+��8O������rP8�Y��㠦a��a&iv�W�c���B��lH�����*B(oM��������j�}|>G��4j��`s��"��o�(֒5y�� �(J2�{�~>GMie_uN��9T�� �}�i�?��"P��3�[!�ft�$�ԍpБ��FQ��{J���GB�[�_h���U��U�C�~ٲ��s`R��$c�j�
&�2��vͩJy�.��8�C��t �{�'�nQ-�`�*]@a+ �HEW��<�h8N�"|����ى������7�������貐g��]	�+h���:׭~x?֣F�U<#��[�+b1�tڕB6մ�
�M=�$P*ƭdy̰�j#<0������tv3�OG?:!��3���<�ZְQ�l*��!|�+�R�D�=_l�G��O��8<%Q��B����/��6���/��},����n^L���G�>2 1��89IR�H����f�'�ݲs���ic����3}n�R#dI{T��Bo�DnN4��h{L��C�
R|D��-=�Y�1����m����6/�"f�w)�1�|c�����^0=�.l}�\�(z����Z�D"m$7�����ĭŵ�v�{]�1�g3_Ġ6 ^Q���E��j�|K5 2���d�F|�sѻy;7*���|F^�;�ѽ�[&�Yfr���lVǸ:Z;��{��!o����*��?S�m��XK���Z2B����El�,}� �<�@T�r��������"�,�d�<8�����6���x�oّ��/틅�g � b��/q�j>���I���B�P E'�@q�+h5i�z�S��'�2��GA��wٱ��+بuNl������S8���_cL��㬯��ss^�|%X�oÞ
��ſ��bT�y,�F����a�>�-cc�F�XO{�`Y�dn���6�!Q<J�r�x���r��-��<���9|�^SH$M�M/��5{J��SB#�ͬ��՚'���������~V�hү�[�3����Ę�owC+^�!�b|�#��(�(ٓ�	�0�K0�-[�Mew�&PG�^&�Qè�[���9�|���Y-<S
@����D�b�QcN���w�O���l���pwp�g= ���)�\�k�S�)sZ_yy�j��^��(ջ�*>�� tȯͩ�e��N�����1�5I�-AT�૷Tm��w!���N{���@�;Ǡj���~@_Y���?[$�8,:�M���FڒR�>3��lc��oً���j�|ba��;�c��I�R�?N[ ӖU�U��Ʋ�&��'�ؠ`�Fx�y�}��&��q�MdE���e�/.6�чYM�����ڝ��V��I93��
@��t���H���� I���-������B�)�|��Py�����;V<���ͯ���(�qF�E�\\���޻S.�d�a����"��6u<�=���b�z�C��#������7�>�`o2�f����Nf�\���`����vK���O��Ae���Ug:�L�	�L�]�E؈<�*��]����<L��UYkfk���s'�K?�x��-"�̍H;_ʇc�#�v��<I(�.;����h��Գ���
����{�u���&�'Jó���-�}m1��+:�,w�\�+#r)��8��rƑ��,����X 0�3���4h���|F�tz�Jlbx��t�+�]U	�E�
�`�Ȼ\��#G���r@��OQ���賁�p�g	��:_�Xh�\ ���$\S�m1���Ta�EjÍ;��񴫈M�:p?�*U&��9�����b�$t����^�����ܦ���#w�(7{B��m�r~�|��<x��Y��!=1�]�O����s�\��!.�g���m���{�@J��+[1^�֤�2y�x"���Oȉin���񫒼vBaR��M<�~�v��kZp����5��+�ziv�}�RCð�G���8�8����F�f)�7��.�']w�F6Ϸ
��YS�B4uc��^x�a��N�#0�]+���_1������_�8ǔϫ�@CH����ر�g���@]t`3R�连,T24x\،w��%t�_fh��-�Q�*؍N���f6�|�m����H�xB5{vl��yȾ/�t�\*���T=���J?փ��\�R<!�V�"�8/ ��W��E���_��������F���~�h&�� u��W� iN�&yG��8N�����t�W�Y��,�`�ϙ������?G(�f����(kqWX����}���Ҷ~G����/���DُF¢?()��ݏ/2u�竐�H��8~Vl���=g ����9�e(��NH�[5�밮�'F�+�m�+>��`��U�ņ�(�o��/�؄X���4��+z�cM�;�F0�h�.S!?��1GSH�)��8�#�H�5��m����|��@1�Pb��6H�h@��	��Z�2�3�7��B���E���mHM��K���{,0h�b����c]n�Y��P�*��U��q;��
�!�s1X�G�zVG�����L>�|��W���~0p���{_��AHөP/p�w�NX��`)�۔F+��o����2��^�sѿe���ޜa�!�O��mN��e;֡��e�q�s΍<b�LQ��0���\o�%�k���-�\����f�jⷞQ��Y�#=��`M���0iNX�^L��?��Mb1�y�&o�r �v�ޝ���~8���f���FL�9]�Su[�<�l$x��D�ĘU�@	#}g�-��1�4@C>�1tǾ],�������f�x%eҳr9��h�)t��n���N�[��#~�/�����a��@G ���Ű���`C�i6�!��Y�8,���V#�s��f�,
�W;v�M�P-��M���ļ;��{v�ږPq+���}V���=���c�At_)eI]���i��`^��Lo��7,��V�r��MZ~(�8N�uJ�q��\Kf$e$r^��N�'��y˝�����r���J��|�O0�Ծ؏O�9C��!<·S��;AVbS��eZ2$lf3����.��>�"��x�>.��7z;�\�F���I��� H�p�o�[�kmŧ��(�Ԃq9M��W�x�ˡ�\�>yi��n�`�@5��zT���:�,N<�^v�z2*���<��{���!�¶�jٳm؛E��H<B�DqTQ�/C�/M�)>�Д��0�>�Ldu �*��>��n�d�%��V��v�@E�5�5^^t&V��=�(����!n��b���(M��_*���j�[4�>P�k����o�z������Rݕ�8�v{[���S�W�2��~�����g����4�Bp�g�	e&[��,� D���߽ ����%zb��#n�6N҆��vS~��� ��m&z�ؠ�� 8s��w+g�B��
�^}���9�!��!A\�nz�O��/ď����3�1Ee��'���I.g��W�_-b����B8���T�I�s��&���ѣ}I�$���Zء�#(�O�az%4�3݌g��g�<�hۦ��X��AW$�e���4������-x��n���n�_̦\5�ڱ:��L��TA�x�a5���Yf%��?�.�'�u���	����ձ`�	��7��L�Q��p
������=��,�Q�!3ܮv����tT��,��QDod�s4
(�1�d><V�v��fر��b	�X�����j�Q��p��Pu���Л f�y���,\�*·W�P�F\܊}��Ù�^�0 �3{69�o6❂��e�����0���T�xh���5=/߂B�A<%#:��MW�;�Ҙ��u����j�VM4�^�[!~���_�j�9�uK
�^&��24~,~�֋��_͗����G��p_*My�=���m�z�e�z<�$�4��R��yr�J�g$�\hr���<{��5��	"�M���:I�\��+�F8��׸�|c	��9�ɍ�V������:�O����M�Mmz�U�_�6�lY���xF��`���]�em݂ŞJ���,�6�=�-SStC�;��]�a����:l(�(^��a�k�׏|�?�^cWd�y6��@3M�gg �5��	�a=��]���l�"}D�𒵱E ^��!c�9y�@x�G@8������!wIx�Әtհ�&VI���JOD;'�EZ�.|�|�q��1h6'�K��, ��?�X/ �FW<ȵKp(����ӱ�1y���I��0$���t�Q"+Z��&:r�9Hq1�d��3dzɡV���l��Ƣ�b~"������мj��^e���RQC�t�XzxVys�r��9��yb2�(� �鶖�4�Q����M,K��c:��OG'~0{h�ܕC�{{�XI��n���A|`lD��o�6�	�r��od�)]�-£���ڮ#V8�6r�Y
\}�du镻��h*�tڢK��kaG@��pQIÚT�� �d�]Om�L�q�	u���gf��˘hPۘ
2֟E1p_4�:\�p���s*�3]����� %���Ϟ1{I� �x�U�j׼k}�f��x��.Ô-{Ug(
"R\P/�Z�s�8!bj��-C���`BU�M3�ҩ�?���D�j��Wn���K�3}������ǆ?�u���}N�w
�W74�D�r�)H&8����VS6(��Y�D��UE����� B�D�f����[����i:)�ʶc�$TmG?w��K��r#j(��,�f-ݶ��gQ�%���>C�扶e\sc�q�S�B@%L�Mǝ],��U����h��^`(�Y�x� F�	Ύ3X(|�:�v��W���p�������+��T���Δ��G�WP��r9vsV���b�hSN�v͋�2�������`�������|�PPJS4RT�u��;U+��8�`Xs���o��r�.�w��/#��|��Y5�m��*N��y�����:��wJ��t+�eJ����jk���?-�(ח���n$�EhV�Qk�]߇��硫ƬO�9j�B{[0�v�ӥ�:��AD���$f���7AR�9$���4x�\�t�m��޽���M��Sw�CnV6�l,���I��6N����p�hi�˄7�V�)��̒�Q���nfزU����;0F���"��&����qs�����抛|�D���l5�`6�s"�T�#�y��)���f����\��1�ޤ�#	m�+W�������μ��[ZB�2�1�j�C��Ȼ^�ۏ�i�7�x@�l�8Y̊���@눹�6@��,��d9Dc��h�? 8l�6���o܆��5�h�g��cY��qL	C<J��L<�Ԛ�ǈ����+�W���H��W�Ak$�Z�br ���X��)�l�b։����Ŋ	�\?GNQ�@퓴I4`�
�8J 7�s� "h��Ew4-M�PgB��n�L�m�רüZ��R��G���Z�7M�A�nnU�f|�+��lB��ot��7Fy��ÞS��4��f`��@�ˍ2���U�9G�Y��}�����vㅠ:���e�neYg�03���-F��X��1���c�
w�I���S�k��x����S���Zk���!c�Q��2a��d.�OZ*�K�E,I�o���/-�kЁ��^����Wh$g����h��$�*����.������xz�4�*��ȕVn�1}C��[�]tQ>S/���A
�)o �I��bQ¡�e0�r���ZI��k��J~���2UnG�6�*^}�qT�/�g��na9V�4-���C��C�mkjɱ�J��Ֆn>hJ"�i�"~'Hf��IY��k��||C���'�~�S��O��uXޚ����b��˴Ae-��˧�QsQ��/���I�4��Wm��I���� �h�b	�U���O����q����{� jRR�3��3YU�n5���o��S��*4�G��~�W$ 5O/�u �;�"!�������97�5'��/d_��ܩ8W��,B��'���{�6$H��&Ek��?C3��U�7�Zӥ�����~~�� Kw���f��s���9:�U�E����?�2|BT�}E�n��Ӌ����J���^z��>�d*��K� "�iVq!��|~���=���G3-Jea��ty1V�b�xm�ٿ�b��4�b����,�*���keD���)2�A������[iq:�Y35.��,Q�-��7�Yw�b�y;B�F�7d�M��\0� ��-����`��bo�m�[��PEV������qo�g�쐁�GBԨ���� ����hҷ�2O�IM����0YŤ�#$x��@0���	����^��|0�'������`B[]Ӯ���L�c^��wҽ�H_��m�-�K��ˇ4K�7�:�%5O�����#�T���U!�b�˨�4�p9W �J�%���m�#�f�b:#�daJ��ViH$-���`�ٔX:v��G��0����a<͎�g�4��z�uM2�e3/��iq_���Ю
�\��_%����/�y�����j�@�1����DL!�ѺV��a�����l��AK�$��	X\9�Sl���F���^��\�؉�=r�e��T*��VV�����U�K�tB�F^s�	ƛ�miVs0�?�&��y0f�O¼��K3����3'���D�3TE�� ���@Zڼ���2lɚp(��V��gJc�]���
��],��'�x$�El.�_ @���'O��ί��c�?�z��_��\ť ��g<��o�'t�D��[]���@��y�Fh�nb �fD��"�Ñ	8L�)ZT��~�Doh�:��87C29���!U�����n=y@$���� Kj�v��9d�wq�y��d����I5�����ͨx�ˢYB���������ZJ"��극#������=]�ؘŁ�Jt�!K�;Z��mi�ۚԟ��I�|�+���O�s�0֬�`�W�"M?�ܩp*b/�-�n%$!-yIQ������c����p���䦝x�B��:�}�_i�v�h�.i��{�����b�~��35�Y���(KA�Eb�l�RԾ�D��ﺱ(i�B���/.=��\�05y�L\M1:�X��ABfs�I#���%k���4�2]���o[Y6-/ (��nY���!�ʦ���=�Ǳ��0�p�
�4��f9b�#����ӷ*{L�~$���P�����<G��K��p�N˵�n2E�jV����*���>"�����D�l1ː�b`~�j�r����*A� ��+�q�v�2��6a	tQ�/����-j�G�4��PW���m�Xv���ܤ�4?���������6�Ϡq��G����[��9�xl;`����+|M��%-��xp=�D���hi�͊;��HD<o��e4���r��A�E+�-i��A5`҆6��f>�!���]����6�	��5���Lփo�Y�n�汱\,1.B�����s�2�d�+ȅ��uOm�KkrBxa�[h�M0��Y7d���	�8�M�ǣ���RL�Xg�msv�l\Wr��S5�{�[dq4SV?��	���ŋF\���������p�x��Un.�h:�[���`��!��a3/aI��]��s��2�b�h�?9.�X��0��c�y����[�[7jJ�cA�h�]�F��'uV��p�r������쬰\*2�i61�љ��	���<&�κ�_��o�Qn��r���s]ۥ��u�^j��������g���5����+�|:Tl�و�r�Fi6Sg8ck7h�����3����B����	_)O�ș����1+�B�5��ދ�+_�r�x�^���/\g������o{��LU�b!�=�.�\�[��0&s�L$�1Ű�p0y"u%�X�:�s\�:��x����֘��pI��
2��U��=�a������c }Z�6�&��)V�X��%b���E���1�6.��f���+��T���VM�p �;��+s�G�ɪ*ǵ��JT�P��fm֓E��{䲎r'��6OL����xS꣤k��w�bl�o��f�ڙ��>E�Wu`���8k&ѺR�<�]b�E^O��
o����,ʋ\��p�O�f6�#���egU���0�O�gй��(n|͝�EZ��a=�:��]^�v@-�+��L{Ou�m�-��B���*6��u�(ed��wx�X�e	�LF����n��N [�	Lp�h���Y�7u��?5�s�)��Nxf��ORQ��Ǐ�B�Y�V� ��������3s罦VP1�+Qv]��܅!t�S8a�"��#�3�H]"%�j���)<�!>�ğFLf
��{�NUZ�O܁b�n�G�\j�7�T[��H<��7O�V��O�R[8r��*4���)��mi���W�ۻ�p:�M�%K7`|�>�d�mҜ$ǧ���#
�ޓ�&��!+�*��~ac� ��ƨ�C��yo�9��g��_G����0�B�I.�HJ
�]��h[`��Dڒ�%�î���-��m�]����"B���쓅�A���/kׯ�cZ�2�N(�����+����	�����y�Ʒ�B�6�ÊeuS�%��ejO�w+|�V:�?������E'�k�*q�wGA�YQ�[�*��*oD8�^�	j�M.���K5��}o��]N�݌�>�;_C���h�����#���̦Ǯ����?�b
Vr�C;*=2{X �DtD�W���nsRѻ�L1b�ksݡ �@p�[$Btvx}�y��(B�r
�~U�S_���E��_f��1`�:�oٳ�L�w�eoz�U�lg6�і��[��Ŀ�E��=�K����GԒ��?,b(�v�����l���D;{���ÎH�^	O�d�����ǈ�>(���[u�.����5w�y��t6\yۄ�=�Qβ����wi�n�.�9���:�L�eH��!�����_/�7D�^�YFzt�?t�����4iͨ��R�R����i��`�w�A��
>�>1j�:�bT|2�2�rW�6oS� �'s���v��w�E�<��Sz�P�jQ�}�⡟��+S�������x��\�r>�r<�b�H�sҳ~h��x���i�z�#���g�l��!�t�-��"�LU���~-5��*OdÏ�R=Ї8�� �\�֤U�N~3�axχ8�����9b�B��M�Lq�!���9ū�`�D��o7}F��^�y�B����PD���3J�\��!͘V�NeTG͠����F������=c��H���=z(�Lg"�a�X1R��An�r{�ո�9��6����ɱ��b���Hƈ}G¸��9@�����ikΌT3{N4)����ޗy"��eMiTt/č&�� ���� �j����R�y܅1���ά~v�[��?��x���B���p!�Z�K�����^�.����k{y����*!���#u��J;ٻ����
�w�9�Q��
�+�� _������#�����\��S[O\�h���ߩ��8{"�$�d�Ԩ�9rQa���P�T���t�?<&�N˘�L��!���\��W�6$��W��Lv��o*L����~�զ2Y��(�0��&>$����#i��0��A�����2r=� ꚿ�(!�}w��z�ā��Y���3Ќb����<�G�\���'��f����ۏ��(�;���"�����JܫU&����%���r���7��E> �=��g -<S^�T�B,����eQ�q=��m����ĥv�/�h[U�O�����v���WK��-z�i��q�wTJB ��)K8�0y#!#���OR.�re�K@(���h|bO���	���x<zV;�(8fߴH�Q�W�P�qگ��X�D��@_�3(��»Q��%��l��?_R�>�*�!Y/���:�VQX9����E�w�5�kR�E��H��� *k���"ŧ���5���~�侞���ɽ��~`���n��ȇ8��)F&>pq�-l���/��N��	^�}�s/�MOV�
5���c�P@CTL]�^��5�I�r�_Q�|p!�����l۲f�����Y?����@Q��wF�t�3�$�O�qɿ�{<Hm��<��YW��c�ܛS�V�7D�$���;Csx���v+���&�z��jX���������y�+#X$�~�g�֢M�� ��5�|�.'`�cw��fgϟ�"�ъR���P��Ų.�q㸷b�or�=�K���x�lz)q���O��7�&k$8�d:]Pr,ip#�5&Y���~,�C������t��s��c �"|]�1|L���3��nܴ�+�����8��Qs_*-[��c[��Ԁ4a����t�((H�q-j���Bk�7��y���-��R�OW#=��/����w�[��l.�\D�Ǫ����_oU�<
>�U��G�/ӟ�����q � =�u�%�Dխ9BCU��\��-�ĸ�,ŧ�� /��m1|#���N���E����7��KEe��]��g(#cc3��>�)����D����-$+�z�M���G�ԧ�s�\����KL�J��_�ת8OY׾ٱ�d�<�p�iҫWC��7 ci7���Q��,��@=x[��;PΜ����pd��U�W�Z��q�:&�"��T�H�1Vl�!��F�Ѣ�[Z=E���w�Y�E��r�v��tV]NL�L��1_�ʶ�k��Tz�9"�5��^O�M�bc1��d(��DRh%�i/��F���|}�L%,,?���_v�iF�*��8�(Rg�mRl������@�쾼mӆz{lk�B �+��Eք+�+�h	NE��٬l~'�}t��7����P���v7��7�`P:󒠍s4K�ޡC̲�}�_H��"�*;F4���u%�]����0��&x�D���(��W�GK�r���<�:��A��i�~�-&&m:0�1[+0�x[O݃eܿ����ǂ9C��w�!v��K��`]���e||�x*�ML�w5Lk��+�X48�W�Z���ua���!I��l8���d����~L��3o���3�����{�D�|�x���De*�0���M�70A@jԠp/�����/�+P���4_���\A��W�! H����{Gϔ��t1��mr�]��mL�n��B�>�Ȫc�0�E�����z�	�-2�Q7Ai����J*��`P�G����X=섢���Gs��;;�����5��T�E۸4Qw̬��xq���톭#�TϾ��I4ͼ2��s���H��j������ѿ��Yܑ����l!�/r�r-�U���|�e��ߕ�4aO�"�Q7�{�@�y�O`�S�1���ɩ��6u��К�V��#����Fi���Z^5�EI%"o~Y�Lj*}���:Y�v��޵�����3Ul�fg�2.���e��'��f�h->�J��P���Ի¨�������#j��+�/��V��0������#��I�t�����f8��{�:p�}�]����%�-0a��GQ�"�G]��h_b��ڸk)|��	=ُ�B9�چT� ����#0��u����~ʹ���1�4�^�~�w�^L��}�ߦ���+����dr��GJ$�XJ0�z-Tl�H$�X9X�0���{��@B�&v�*{{�E����3F�-�a�i��G=C�g�Y��8{�8T1Cmo��@2_�f�Һ�u����(H-R��U�7�Ki@�[�x��Ff�2��j�Am�͒�-���iv��C
e�̃�W|�QaK���n��& �I�',:�$�L���y>���z�����tGq���i�t��Xd�5�~Ë�ע�M�S��;����Z�E'%��u�e<�:Ŭς,j�M[���c�P�3�[�#F�N� gTU��\w@�R�.R�>h���˿�W���3)�X�qO#��� �î6��*�Ԍ��ߖ�(�qU�%��:<���G�v�?���b���zޝN��C�/*�����*sa@��r38��B ^��޲���B�KۏD>@������ݿ��Z�Mx�[�t]��|�����兀�o3qe��ԛ��4S�	����F.o�y1��`�4X��ϐ���,���)�æQ�o�w`1�#�19��������KqT4�/6��A����n���~�n�����CT��_���t��᣽��,�㗌�fr�.��1���׍�έ��﫶D�nc)i	���	Xب��"l	�?|).�y�����[?!O'�%ɤ�c��qT�=�V��C��@!�&�!D�sDP�hPR�娏�����wE�$�ܟm��A Y��!�k�	x�~-&�j�k�)҂��i��᧤��]�FY*X���N��59})���FӃ[��5��E]C9�{�7�a��	�$���ZE����,-Tx�F[���u����(�@c�
��! ��GE	5����C��o�{f�����d<|�Io樭|�Nm_F��b�F/��?��<B[sC���5p���ph��	��vS%�^�A��Et�Rő=ے�89xg@�ʓ���#�Z;��R����!|-q��v	��gA�J�E��c5�R�w�.a����4����F�("N�.�'c���H�dh8��Xb �l��CM4O��ųT6ҷ�w~5¯�*��	u����z�5k8ڒ�(����[W�4���%&<�����*}w)�&�������\=�%�����܋����jd��*�
��[�`�yۃi����G���u*l�8v[Q,����؀�p�IbVC_c�ˁ��G�͜�9�IMDǖ!%^i��_�� ka�I��;���L������4tdHI�0��%�,�v���Z�]0}{P�̹�vԵ�� O�w:Ը��ǰw�i�dȯ,;����v��QȾ�XS�9��\Ǣ����|N�zT(�Qc�v�[���^����W.��y���@.$,�qt���W'��N�
�����P-y��՞�Z-E�!�
�q��Ү�f�1�͠ZJ�%� t�w���S[���|RO�7��݄�R��y.]*�kn���3��c�t��*���g��Ş9$@��7�7-�#±�0���%�Z��Zo2��}�Q�ʿ�um�i�s�E�j��#���m����y|ڒ�}2 ���n7�%qD�	��a0(߲�܍����r�% [P��-&اAR�Zخ��v��O�����jG�:4��At��]�P��9��0�_��T_)7�@i�u�i^|Hc�E�DN�ٯ1$"w�����x�E7��sS�rS�
p1�QYC�IbX��#_��#qRY�H��	��PG�8