��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�APq�lG!7s�H=s,,R!���#���$aFͿ?J|Kf�)���	̚�踹j���#;�uv]>ET�	)�;�f�uv��K�@�q�5Z9|�<�Σ˲:�������P���6����}X�YV~��n�2�l���X�9� J��1BH'�P 0�V���6~n�ƻ&�0&��x��M4-<�'��8��+]	��ko��T܅�=2p{���f�S3�'�H�����`�z��H��[�s�Ҳ&��6l�s� Wۮ����\�z@7s���ިUo�C�=nR�Aw.J����_��,��i�	�(;[���yh�[ͩq��J�|�7 �H�>�R���1�����,����±o��97%e)&�5/>Xv�)�)�;2 <���sXy.�/�Rb�cG-�ZkTÎ�]�:�Ȍ@Z����+��(��E�ICS���͐.;�O��c��rY�Av��
\�����P0Ә��L���,�I5��&��x?W��L?��G�e) j�_�}8���v{k�+����g����AZ�C�$�@�+0���o�0Ho{~���x��������:C8|���f�d�Z�d ^��{� �~�����Zav������o��4�,2��
i�o�h"��Z0��?'���2^ ��7���k�Ղ"��@S�c%7�d7M+#+��R��@�$eg���"�bl��
��#��?�:F'"QR�'?GH�:��|��� Ŀ@����ݹ�I*+���H��F�ރ����'� �Ҙ���Z��i�#����>���A�`�������d�h4��(�u�k^Hz�fv��q�g6)l�Z^�;HT���]�����!Oa�[���	�ʡ/�ɋb_���X<6J���	�/�s��	 䥪D/�-�HLu\ֶ��A�
��'� �ɨZ�pDB{�,��%����Z>��_	�(~ٌ;���I�3�Û�6Bؓh�HJD7x����x�P����1Q�bז�WV��"�a�s�iI
�xt8�����z���h ���{��*Q�'Ѵ����^#���:@B%����xsq/�w�/����թ=�ɗ�����!-1u�{��>��.��v��y.�s"�e�h��B$iy"8m�3���qQ��
ڷ�-�Z�9�3K�j`h����q�<�N���B� z�b>ț�����q��%���!�K�ҵ��J���sR�Ű�k�y�%,Pޟ^���Q��$�J�ژ�^K{�m?�����8�(��(֮["����h���k�U������+sAEu?^�3���G/�����b[���$�`����b���K��_�	!'�ݚ�np��A0$L�%i�����qqR�<ss[D�zؕ���涋+n�h���*�w�N�X��>��`���뷼��3nt"�ʞ-�"�UAq[�� OsHbp�u��ŀ!2�.o�#h�݇
!�A��3t�(��>�)w��!�Xt��<���8 q�Z#���І:5urX�|�;R�^�mw�����]y^���,��qP0 ����b����B^�]Ԋ�?3���>�E�|��� l���<T���i[0�0�m��]N�Xy.��mm�	�lr�P#C�� #@�'��];BtN
����~������iؙ�˕��y��A�`��������n��M��q�=/�9�0W����R^/��S��s�V/C��:<yK�Bw�����b��ؙ55��
����}�VK���QI'C`�,�R���0J���+�����c^G���K	���+pY�6V?&�j�� '��)~GW�7�b���ƴ�f��\��q8SC��6R1�)�쩣xN]'�0�� Zl4W��~`�^��K�S���H�#���n��/�ɵ���S���p�v�.�H��:��/a���W�޻��v���h�$�r��]Z�NS��#��ˢ��s��X�{A塂����$h� :�	>�JN����D��=��%�VPL��S;��M[/S�?	���Q7���LM�Y�M��e`~�4��}l&Y�1�`L�V��~�u���ݠ������.���!�2�����l��´n��5�lu�ż�H��K��qmb�IX�3�U��d���=~�;s���L!�P�T̿#mԷ�t��E��G���I�pX��`jb���'�������s5
���E-o8a��8�z|�۸�ܤ�<p�@��E�� �iH{ ɾ�ۈ��K\�k���#F=��!�R?�����ω�3�V�P��H���	ً]�h$ ����	�2���7�����\�4�3_�.�UT�n�6�:?�;�Q��~#G�9VL���*v�SV����|�9��!^��Š��|E�a� G�dѺL���&���-��W}��ZVI�L�Rp�kw�q�:�6V1�݈0I�F�<�q�nc+!��W~d��fc�q�-�~�`��T��WM�SW�%��Xc5��Y���\�18��������f�\!�W'��P�f=�+�7�H*���ow�Tix)�ٷt-<y �'R'��.ء���{���j>�a-Z@�����ꗅ0�4����2���d�w	x��P �6,
��Yc���!ѓ��$��D-��2TO���;��:j46s�WG���?���Wo��5�>��ȩ{�o�Wg?0޶���0���X	����J3��t*A+��FK��b��J�o�}�!dŎDa��~&|�h�L�[Fz���d�d��2^�zE�����F@��-p�
�</�;�c"&S��	�.q\A�c���Ԛ����~�hJ~���(�mf�G:�΂Z�6�'T�ᾆe(�L$��9W���d��sP�.-��C���e���j<B>и*�m�CBJ����	k��.4�@Z]9x�k�!�K��7R��|:�޿�ZXߦ�� �y�A�w�=SH���3C��,��Ӛ_�J�ڂê�ӂ�4M��%E���G+�b��X�+��o%۪�n�Y%��ؖ<Е$02e��*��,b	�/�j{���ě%�Y�5�PٿV�#�(r�PU ��C�o�bi��b���m�%�������-�;&d8�������#��so�{�ޥg�J%����&�	����g�9�&}O{ε�}5x�ZU�M4����t���g�.��z4�����'$;};�S��܃
�G����g]�8��G�@�x-PO�y�Zr��_�|0��ŏS+yT�"sy1r տ�ލ;���A^o�Y�iUeB��:N;X�����3&i�;�u���˼���r��Rc���K`��$�	p=-˺��f���M�phNV s�]�K�2�gR���w��b:�*gW���89+���n~��7Z&_7O��-���r~��9��A��UV'r	��z�]8Ny�L���Q�{����r7�x<M�B�%����Q3f����iC�N�b��%�#�V���no qcO�]N{l��S��ǁh�v��ы�뫀/� ���E�q�ygM�ܞ�^����x�˖�&u�O�zb�䧮r����3�t}TַJu�o<:�]�n�Nܧ̞�Wod��C�Գ�k,8�t�>IS!C!1���6k؞�X��+�h�$��?��ھ]���^k)jtr̦�tn�#�v.|s�;��/�l��/�܄��M�1~Ղ.��ǣ����|3�[7:��j�[����:�ƛd�!�{
�WD���1������>�_*�����gnۆkh>J)}X"�o����!6�V���.l2:�*�X�B���-	�.ƙ�1Zp��3)sh$��M{p:N���B��̾��=FqêJ'�9��"~��W4�H��r�/Ͱ���!���3��uU�h#�kIS�j�#��������ZG>�E�y�������w7��q��V�ʐ
W��=��9n�J&��%5)��̓�P�w��|�&��utF�,��X(������i��ux��Sg^�4�ʻĉ��:f�$��F'�l�^l�̏�M��&����w�K���]e�EyHݾ"�g��wխ"�D��X-Q�R;"���.�����'���|k6�jF�O9L�Lx;r:g�It@��){�{ sއ�m��ga���3���٤��RB�Y���Bl����J��A)\@��oF}ʾL�e��#��l*�%�l�1�����r���X>h6��MO���7Thw5�#u�b.��|~��2I�)Κ�<�%��OY����c�7FT���d�=HG���K�`,0�t�~/z���?�.�m��	
�| ��qS5G��ر�{0�Z���O�J@<�����D�=co	5I86���y�\� _C��oٟ?�'Ō���C��ŊD�u�1���Vv�
r���4��v�"��F���+��~��A|^� � �i��HN���0�4���3b���=��b�1-ƾR}���t����T���,�12S}c0�T`�����o��"�F��2TCH�]���o� ��&��ǻ;�qK��>l���z5)ʘW43����*:e��,B���EK�?>�]bi��<
9�F�dw-��\��c�"����7�-��yZ���E���Λ�N�ޘs,���"w�?���.�����
�[A�W���|й|������N��p�.��I�}����K�xl�@���'3���+���3ߋA�8(��,����K>vCQ�#q��Hܲ���h�x����-K4��L)W����Ƹ���-��E�+��ZҔD�7!�}=p��22Į��H�p�)���J ��h�q��Z�6_�ސ�BR�M��������\�SAQ܆L{��]���D�;�����!JYO�v��dJC����Q�H�xS�`��
�������/��f�2��,\)�_+-�o1�b���҃įΓ|�����67�Jz�iKHE6����g��t .��Jn���[r̓t�0m>й �W�vk�P�v���5`-�^)�w֒�a�����Bj�nD�l�50�8�")��J�o��k�E³I�q��?���� �y��5S]V�͘��~G�\8��V��s�ԃQ�[r7n�]}�%G����Nd
��8�6���
�X൞+�����#���U�rLD��_Yp�^�F�&8VL���V����͇9$�a�l;o��%�)|�fF��:�C��Vh����X�w�H�&� ͅ3y���͉f� �H��(e��-RҤs��q(eoa&�K� �_�(�N�f��.e ��$1�OMF��d�X����i�^��e\��}����8�A؁�T"�|�c	��2a����y�Y����7V?_εG�GzYt�9�B�"X|��{<��1��B�Wy'd���H�{�����˛>@�
�� e��:fʲ���y���bO
��浕Bna���4����~M������2�wY� l-�þ ?Kx;s��PJ��h-�*�J��rHs8i�3;���t��<���D�Dk�l/�˗?eHh_f ��-Pg m��c�('9w]�v�ɆƔ?t�;ى�ˍ,V(�@N���*�۟��`����c����
c|^��?��%��A �T�yJ��:�N�D�D2�l�Zx�����{��u}�0�"��vL��{�O�$��徦�O�
�թ����z�6�8��s��w�YIA�ﶴ2����"Ey���޶;{�zR`	�+S�>���=`��q���P
o��8L�=���:2=������GoT���pG��&4�c�����E���k�{�����:�n�]�A�1'��CxDk_&c�Fk��va�O39=KK����l����sL��M������1�B`��GP��*�ӧ�| �ܕ�#PY�j>p���S�ĴD�=;�|��M�_�;"��<�l���|�İ�[���c�W�Kxl^�FͶ/Jab�	9�����a�ӵn�J�Ę\���M���ݷ3o�F��d��،t��v|�#Vg\,������Wc��<T���lq�&m����F�JMy�	�)�A�y�x~j�/9#�Xn��z���+:�l��7�bY�I��P��_�|Ʀ�[�_�)�0�~kP�6!՞���)�)�y!�����+�0�>�W�@�����*͎���r)���Č5�]y�Ӯ�-�1�jt������z�ـjY(w0����Qc�B��9k^�o���b�!�����ٷ�~��V��VL�|�ϸm�r��f?Nb��R��-tD�6C�j��UW�K�篈 WT��'�9v	�NO�����r��b7K���K|��	�G]	��[��_����	3��/&2��w����[}�S���G�T,��y���<f��,v�5�<��bγ<WF�TH��)~�,h��I�:(UH���Z$��{��b,��b�p1+��f"�-�8a��]��s�Y�����E1�3���<��!0�����d���S��ߖr6$��z�93�ƵuN6����=`�861Şe"�ˠ;YK�R�uu:`�ۃ/!�O����Z��߉��'�1Y��t�TBSr�ۚ!�@P�=��37�ᠾ`r�V��D����*�ʋ+}�&?�,����E����1p,��>�2��8��`A�8�iA0�
��`T%C�C�E'�)/�ȁؒ"�H�+���jUH�(2B�3'�:����无��a���5+���`D��1`lx�X��ك�1�������d`�WZi�-��),q��pL�Jמ<��-�f��Y���M����-2������*�u6�h ����l9�1Nź�g�i|bW5'��?����HLz�G�*��5n��/3�&�)�
W��m��W�trx��c����)�d��V	~3�$UY���S�6�����������Oz)�Y:�F��}��ez�q/�G��b���<ZP�̨�"+�UV��ca��N����ķQ��2�}5~±����63�eP� ���{Lz(��:S�?^8(A�^좈���yj����7�]p�)�4)������Uz�������ڰT=���vD�\3�8�����BV?�͢*���-ݚ��[�=�,�۵ɠ݅�������k��w�� 7ɿ7��H"��;9zQwN ����3TEir��ӈ��+����{=����۫��h�qܬ:/�e.��`h������6�G�>ͯ>�)��&�k  ���*v&�4�͙�i��2�UaG���Ki��	f�t�.��7��^�L�]� ۸�R_8\I7�A�1�P���-���o��0%=���o���5+Ee�.��l��>��ԩ�$��ZiK���0������4�p�C �-��=&±h��h�n�FW��)	�ݝVcޝXЌ&���{�����T|�ũ�A�����
N����RK��(	^�#\��f��1B=�/*C{�B��{�~����oWEoQ�u&�=����p:���U���/�<�^'d��!+ћ�yW亝�� i��2�F���uJ/�<1�f>R�<��6+z"^�cF�y�c�u� UV�����pyb	�F���wX��g�����T��nѠ��y�[Ӛ��c�.˻�䆎��팼�$S6���;�+v�nJ��ΚB瘭�\�?��-�����{��^�T/��L3( �}8,劉��y�*��?"+0���/��3|��ZD�5���@�OM�^����:g;h�i~�ú�	!$H�q���,O:.T��8���L�}��x����3���p�l%�h��
�s>�`F�U,0�o��ց�)y�����myr�&�@��y��8i�v�Ӻ0i��L��� )���S�t�$����mh�.�XF36��$�ei��GEd%#+�nYsh�Q�d�
���0)��������wZj �'�O2�~�,A|/`kX�wߠU����f_��H�:a�U��`VU�F$�T�j>�� I�._(흈_�H����1BW3s��|�m���M���V_��)aYGh�m�<��ӹ?�Hi�I�g���5��s�H;7Qq���Ģ����{�1��77��\��T(p�Z���:1�ުVk�G�G4ص�%{A�]��Vω�A
3��x�C�/.�T�I�����ơ��i�W�1�1�)U�	�)i��dd�2�:Ⰷ\��#�t�Mu�/fy _׸��r�['�����5�*�F���Q��g���V�N�Տ���wQ�&͵�|Zp�v��	e�t�o	��b����,�%���rw5C��䮃
`b�'�X洡�O��j��e�3}������[Ad����%�נ�3��A@N@A��l�G?L���E-
�3�a�SJ���PV
��\`���J�|'��L�5�g��B	)����Fg�~%����V���ƥ��b��G�����C�He��ǟ�޴����A�uOQ�H��ãc2�0x�ܑ�I��4uN��F�>�|�L��2�N8�gŵp�d2����t�����R�8�������(CT��q����mv�k�qLa��D
�G��5�@1?�9�e�b a��4=8&������6?��`3�9���=��J�H��.�%��]/y߻jA[�	��r�5�3K�J&8]N���%k ��1�fV^:n�ty�����J��uPM_���8Y�@D|�n9fL�������|B�i��p��M*J�3�Dڱ��CQ���7遳��Sd�RߺW�G:�������L�$ۗ�!�{��0�z��W�+G�{�pn�s�Wd��������]�]:M��o����W�.�dE��0�N�����W���W�����Vf��?�w)��J@�ɾ���v#+&H��>��d�Ĩ���	F:��	S'~�J,�V�!G1�C�)m���S�cc�\t;��E',Ő�#��L���¯$�Y}%c��,���u��p�iJ��}� jM�.O0G������n8M��-��d(_� �^p��H@�����l����l�֪~a��y�n9'7aE֓�t��@=��p��R����>΍-�v�S�q�R�E	���)�Ǫ�m$S)3�(�^k4or��FM��)e�i��L*��IɌѣ�cp��?�y�uLTϴ�_0@)��a$���(��&;N�Q�]�R$7&6]�~�	�<�4)�q?5�9E�|6�E�ȷ�Vω��)���\"��\��i	��� 굉]r7��w�A�l �����/�z���aXo����X��L%V.�s���JM'�z�G���$��w
W��F{�WPw$�r �qq:�}3��'k�IcǞ��Q����*ORK�dٜ��~{���W��ڋE��o���C��blx&�Nc�8X�(��ʫO�NU�b6U9´Q�a0kX�o��?�?��%�*3+9Ԟ����� �^2�=��H}f���� ؄����E��3ުd��A�xs��ꟹj�l�%-�ª#��ǥ���L|�y�}��w6Nw ���b�.j�j�_N�r��LWr��M�� 5�F/�J���n�@���NeAA�:󠍥1�e �w���*co�KN���,��������W�/��cW�f-ܸ��{��Sk�9_��m�8ݽѿ~e�@�\Zdp���&�#d����8��Vn1��R��BFg�ؖɇ���!�4��dMl�ɻ����#�����<�<�J<� !��L��3����HiX8&���m!Z���J�?�ߝc�,�DZ�o����M�G��66�XNs;�~L�ez�1�q�&���˕J�Z�_
����Tej�iB쇐�k�y�u�Z0	�}�/��.*�v�^����^���js}��h%w:��Qi�i�%9���Af��֐���qGob_�@ؚ��綏��UE�]��g
A���=����,�j�� (*��� ;W5&�T0�%����U���a	��Ģ~��Q���ԵQ�V�}�>Ϯb�օf�]���݋EsთHnM����(��F/�*Wy�I�5���7���`/,��`|<LL!k�z0Q���q������'��q�a������c�b�b^{eZ�� �j*����y�K �	t#;���;��
C�C�|�`D�ЅvGz�6]�_�"��L��϶�1��eb�[�r�U��g��;�t�_�_