��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_}���l�'���(p��9��^P�m$n��B�`~�^�%�L˲�X%4Ƨ�$��I�5�z.8�"�hdF�����D����֍��\���(7�BW2�����KrӮX��\T�� ��kh<�:�?�b�.G����%n7�B*��{��n$W�Q���t8P�\J��t�q�Q�B[=]Q�(d/?7cb�3u�n>{�d������n�'v �̭N���"�`s�'{��=���g�#�1���f*�a��(��
`2�
�s��=iD���,X��ž(e�f�Z��m�����ib�N8����1�f�|Ia�U|���'�5�����Q�L�%�-�L>K�^����{�x���V�o��j�K��vo�u=�7@�i���Vun�c1�	� ��L���G⠨���y�+Ə���q?������)��Ї5�C��^��<H�E %ھ�2�]�v��;�"��.�Yr)x�<*���~��p�}Փ&� �n;Y����Hw��ЎҺ����-l���ҩ�iƠq �v��=Ԫ�Bu�2��;�s�)�Moח)^Dx��ͻ�5��S�O�s�F�o-N��^�#��k�sj*�%Ӻ=u�����R� L+$1��Yt�����|���W����3��L���w6�+��z��BW��z�:�qz؀]�t-�e����#@��m��L�=yq�ʄ�.j �x���;��n0�,;�$��۶:�)�L�B�n9��H�4���?�hwB��q��kd.2�Q��3ii��~B2�l{9).�{5��X��d��p��H�E�r3�!�_uԾP�Ҋ��u���7
��_�����+RO�8���5;��C�}�L���gx���?ދ��}��o�� ��0, �x3u���(�F�G�K#�l�B-�LC4�Se~�-$�?�M��Ed�x�d��[C��XL$�2�mӉG��T������&�Ϻ�p�3��#P��S�T�X�"�Y�ţ���� |N��	�ޱ緹rY�I���)=�K(�]N�����=4|����Lt� �"4kĥw����Ǩ�NRz��;QáN�}^|���:*D������Țܟ�;��xKN�Z�oC�DFI�&X)�8��ZR��ɱ#&$��t�aJtCt,�j0��7mm�$�EU����b��7�]���?���6p���:s�([�DSI����J��Y��S�e��)���鮦bܳI8��[ؐl'�/8�Jt �aƻ�4=� iM����hH�S$;.�톺X+ )��܉^����J�>�X�v��\� 9?�ǝ��o�O����3�������b�""Ǒ��;�tڞ���38e�y������_��u�_KI6G/&�5���	��A��������z���,:�>��{� (0�5�������8��$?-:l��bIl��bأs�g���
I�t�[�x�`�dQf�B�_6�7w��wԀ@6� �0��^�[@���E5"IG��� ~�8XЂ��]>A�	
�`�������\�-#������u�*�����=`�w��&��1���A��@���y>�S >����攃Z��6�HvR#�y��-�0�),�18�}�:j������ṅb�tl���}����4����eHҦ^��4�ja�w-�ݿ��O��堺�P^��6���d���A�V%��R���j�9��Ȍ�b��M��O�a�W��ū�N����|n	G��']�����r��/����^�c
�ٶ>]�a_ �k\7��`K	�ʥ&�|?�;�Ӎf�$�dՀq��MTLi�#�}:Wk�������H�����3a.)`�9?g.]������V�{�����p5.�T<��	��|��)�ä�o�MiI��O�VLb�����+�$�]��6c�#.�1J���(��R���p�h�Q�l������;M�L��Mّ{L���ư 'Mؼ�S0�+�/-7~���7�&�D�5}��fH9G�b��a_xkQ�(�O�J����ޡ�5��.l 2Đogp��
�4��]��)m�Z�� �Y���E��-Y�g��^�D��ѽ� ǍO����� ��
C�ſ[���C�����P\�swd�V�P�^���/�+fHK���zWhQ@�`�G�vr�6uΌO��Y�G��Z'5d���*SJmV��"�E8���G���
���tL�����-��iQ;˗Vt�q�O��q�yYa����W~M��$�E7P^���Y3�@@�4?".�,X�"z~`_�m��ɸEٚR�����������T��H(�lsv�����H$�#6Ke������~�W|Ko[L>�:x��a��d���t2I�5���`���\���J�}��lx��|N���շ}�zd�ԗ�x3_�N�Fi�(�a�/a��~�+#�?c�
�T���h�g�تc�x�&(ݥsn?��_�c��H�����L�"����k=��sc��.zze�S=�����7��#��5!�@Ϊ���ܝŇM��r���,U�W��R� @e?e~�[w����vXV���@Sm/���<�)��TU]$��kq"���������&��ѹ�|W&TgOC�!��.�t�]8����Q���`e"��z�~;���ՙJusՋrm9V�`�QM�Wj�ض��q�I+6���,%MM�5��U�B���W�X8 "�oC^��Ρ�;�K�ov��y��E�,��>i���j_,��U�_�+�^D��3��K�l���$�0��ژӐ�H���6�������/�#y�Vb�$t����uI?�V����Y�M�`?\.?�r����q+1�����8[٤�sK�=�t%�O%�SU��<h�:��
��������ؔ�'*kvr�*�=�O��1���ⳃ5;Xqٳ8��*0\�M��K�
��.,MxLm�n��m�3��Qq��1��*6���S���7y1�,�,� >n�};��1?Q1��?TD�zZ�2G��kN�^��r,�t�����
���᷶�據��a�&�N ����ٻԍ��\�R�-�F��cy��y�5�����C7�U��k���,�,��>���I��(Ȟ�JD�O��x�Jh��&�`�o[��f�e����%��=��@*�������lgL(�&0pU�^��'����d�=�� %}-|���gq��oV�l Y�d\c��r��s�~je�g.F��J0{`�q�sZ���8�}MӠ*!�T����jf�り��k�9}��\���W�'�L�<�
|����j7��� ��P�-��W��)�6Ǳ�Z���j�P�� ��n������9!M���L��t#Z�95W��|�r���������������i�e�q���9o�FU�r��6�h�WÆ��C?�K�\4v���fj�?U�S�U������D�&A��_]��9Ӱ���"���'ҋWm{4A
�z�E��٬������h~��T{:R��x;U� =��Qv���]l�+�:�h�
�3�֑K� z��ќ��� �p��Ϡ���09 �쭒sU2�[�2Mޝ�`��7:��A��r��(����XqP�Z2�ޭ+���7K�K��ԘF��>8j��HS�@grU ��|���
� }�2���:u����u��i�5��~$�=���!^Y@[Q&fO���A��F��p�'��R��
�4,#�OA��
���3a���V���>��_�O
��փuL��2�1���+`Uw���a���(�]�p�JG����+���[}�S���	��j�bD�A�Q #�/��	3�N4��y� _s�8o����g�h�v�e�*�R�*���6ŗ���5ĭ��/���{�u�=�3�1S����O�	�U�ޖ;	(�DUWZ�eT�eo9KY��
Z_�P��o%���u?�/��d#̦�a7/\��0ѯjM4tj��)VJ�w�Ex�������e�� �_�],:��ƉB����&P�¹�	���ٟ�0�Ȁ	��hCv��V���;�d����x'�f7)�N֋�����[Ģ��� �Ń�=h���~Xq�Qy���K��������d/�#����>pi���z>_)iw���z'��o��=��£�}y�����>�^D���U/�#�.��Q�/
@_�H�<�Z<�ý��A&�,J/�.�D'�VPk:i� #�ɊuNG��� *��H��RF�S�K ��5��9p�����V��/=�!~��5�H;΍����t��ߏ�geYCM��ԫ]����2�}���+��U ݺs�C���D����r��=��6t�q�4\(5rZ�p�؛�`֓��ի���r����,ף?�NXѫ~��]��{_�W����t�I1�;2��a��=�(����K��=%̌��d?�;+��Y�#$���R-9�h��%�Z܍�_��2���_o�������R�	p.�y(��Ԧ�j}஧�SΤ�k��Y��0A:*9�Х��`�4G��ps�O`����j�M���H�(�m�V�g���UD�w�ɼ�Z=@͖C��l}��7f���%]���(���Yr�ѳ�kо^��Ʌ��O�d�<�����˾��CTL�s�ߠ%_�6U"�qj7x�����NL��_9�>�	`ln��)�/�_��f���UZh�`�1}�KR�F�U�L;mCQ�đʼHe]r>�r����}��I�Z�{�}��aL/���XStߍ,��@�t��U��`�$(���8����<he�S9�z���n�k+��>�#�W)���eYV��$�L�<��Ν�;�"�N��7�������5�N�\aP�W6f�z��"#/��Ȳ�l���"��;���qV� P��K}��4D�a_���#�̓Me�d�e�;��N�]͟��C�a)x��H5]{T�kms�T�?9��_"��;q�6m�١��F��/x�e�|�!�H0��ĺ�X�+B)��7q���j]�$��C�ѩ_�EEn���I7�����!ˎ��J�p�&�&�>�-�-�[!���d�s޺���40!������@�� �&'��H���٧8�i�[�{�V�W�R�/������*	�|k��Cp~7`×aW��{�0높*x<{S��ڭ&��I����rlv��� uHA���.f*�q��t��
�Ե�ef�MH��i�8��:��ϸ'4�\d��'���L������]�?�h{$Є���0�,��i�1��FkS�i�T|q8ц�	A����)_B��|���JX��ʤ{��e�ݺ���H�@W>�e��$a!��J��c�	-�K�!޿����?��a?u�Z���r�+��p���X��i��
h|�`�o��Uk��ె'����������O�g�B>t�v!<��W�C�W��b
F��6��s'�ߞ~3���	]p�X|�x��z^B�/!~%DCO\�~����^!���c5����$k�{P���0�#�e0�*?F|��':@Z|o��V�g�J~����láAz�~���U�[EM
�c�`��@v�٘�(1��AĤF��gcaL�hIGH��j�����3�S?�~K0�����9I�|��8VL�+��đ·^ZY�fBޞ��k��ƣԔ�9[R̉/D��7��=x8�����f�VW���o��s[V��������F�C}2n���+�^Of����H��lhaƘ���OFm�s�3�&`GI���%�+l�{�"�{}�oC�?��O�/�K!�ŷhlM��y�z���<#z?�G$�e�J:^�����\���/��Q�ܵ�Y������Lr�k(C#:���;YK�\wt!��k[qs�틇��|*W>_T�(����/�.����t�]���5%��g�avB�ח��o��](ތ�َ'm�t�m�]T���6���ɼ�[t( �f:_謈8��#>*���u��v'�yl�r��� <`�J{W���H:fO�9�J6.>YF߄�����B�UZVۖ	fM��d6QT��C�P|����+�C�r����Z��`.)�LL#����O���;ݨ`h�h����	ױ���Fj� �`���i1��x�)��.��a8���v��92s'�v�y�-�FIp�F�"�F*kb���&?�8>�;~�LK&�dڂN:e�S�Ʀ�p�	��n�qY0�7ޖ�6AJ@�w��/��Qy*~�1�.\#qZ+�����a*	�Wm���SZv��@�5S�`�+:U,�GE���&UW�&��]��!ԐǑ�h*�^�D�=#�>,���	H�m��i1�	���y�7��	üw��Gw���5�m�d�>���#|�^~�ك��Ikr�d�z��pf��0E�ǁ�懭��~�A/,��\]������"Q�ϊN@J"fѲX�E�s��L��;�՜/�>�)�F*�f8�VA�&M���2����L�\7��d��l.����(VbO�6;���E[��}��E�w�!_�}��;�`��_�:��*����b�rx����l�&��2�6���X�<�j����8)��m�t
���-���1�W��$<�D�_����	�I���lLA�L����sUԈd28���\�o����2pG9Yh�.��H׽��{��V�W������\�:�!���rP�`�� ikXu���+9��:�ĉղg�}��NH/�S�&���(�Pz�]�c��1�7�9��j���`�%w*��l���������쁴����7��Ղy4�Ҝ�9X��T�������Acer�[�ݬơ2R�T�T �V=e�E�)7|�yb<Ye~?r��'k��aMZG? �e�6�Sbё6�*�t�J���o�t��"�&75�v��n]@/��Mhm���8�7�Ћ<�y&��`\���������72W��U[�Δh�@�#�n�
�rPz��]��1ZbR�Tv����$�bkfX����;� �L�A���!a=٤���*��U�� /�]i�m4��s��IG��*���
e�*�����u�|�H�f"�H1_]Z%�~q�QU�:N�&����7����Ac��XY�-k*L&N/�
LX{���_���9/&��O��!��WI�L!O�����T��>�Sߪ'_���������XıQM�9s�ս��Pwrt���ٙUB2$���f�o)M�'M����~ߜߙ��b;҉�+k�!��E�7������Bg����lK-� J�#�/B?�a������!3	�J�FU���=����<�wz1r�0E�ŌVWf��0��Ȱb������S���z��f��w6�Ј"�2{����́�8�E�{W�ޕ_�-��_i��F�T�G7¶|���0��[�r�?�4y5ԣ3,TB=�:{���N8���q;ͫr��r(s8�?SP����o��|���`IJ=�Lw����/�&j��(S�'��}b�`y=zȉ��A���ԏ�SI*~
C�9����ꃧ<�`<���ʩv��w�Ķ��B/ ^1.��x�c�[H��|���L}��I�mC�ܺ�u�H�gޞ�%�OĬIIyϋ����ZW��M�zEre���ٰ-���X�礒E3�0"�u'��֎��aYL�J��e�bs�.;�5�������?Ё4�	e�/`uTo�3;�Bp�턒��%.�:6͐ɸTF����N���2qK�V�|���_{!�_o�Q�������wl�z7?5	��)ޮn�Ӕ*�0ުPi=u�����9�CM���>�l���N���:��>����VH�����>�]F V*��PJ�M������"�o���h�N�W)-�:�i�>�d�/B����x�R�Da����`����A�F����@��EB��(T�.���̼@�:!�d���,	_�q3���Ƨ��-O@|������쮈3���s/?1�rK3H��r#����Ů�n{\��+�^�$L���2_�j�P@f���c�^�KZC�#K�/��p��0����l���l�wu`��:K�nA��¯�6h<S��;{٧�����i�����ﲪz����E|Y1u��CO�����\���ٹ�}v�a��7�1&z/<	�R託�ЦL^�K���[�, s�N�|y�����yc��d�3��q�/�Y�P'���(��[����|�`
=�kjZc�y?�j#�7�Z􄫄�"ç>�L&᪎;�i��n���o,����V}-��,<����p)�T7��-�ٽ�2�R�B����
�q��d+��.S�D%@bg�c�9/ֿ]o�"��j��$��A$!�?F,$#fluy��L����o�2/���zx�O�-,i��3Y:�1�����}��o��/�u�?Hc�xW��]ͼC�gptĹ?�H�}��.�Q]Mn	���� |Я�w�����V�xr\��/R �#d��,��f�'#cC�!	�Ѻ���%�ų�{���q�� l�6�c�/x�g�[T�忛-�x[��Pq���7��I���(:$47q�=%%�i�S�����G��� �C�n/�&��$t6/����w_�>�M\[�>���J��򘶨��Ok�h�hU�:<m�2S�Ѩ�/��f���d5��V��'A�#�Bf9K�=�n��Ѯ���r�f�Y�h��?C�y�U�a#" �FJHQ ��)VCX��� �/)@ �K��`O센7爮N*���f�f�\�$v��T\9+����r֑R��D8�/�
�mb�k�in"dE����u%��Y�	���!�J#�V��4'���#j`r���� �\��3���D�`"&��nW�v.�)����߸��k�P�49�.�U���4�}aoBq��.��0�e�
&���!��}f�|�`xH�v%�v^$�(�~�K�s�s�%=��s��(~�QJq�8I�{$��:Ig]s�IU)�Z.�)�G+P�#��h��lO�w�}݀��`B�8(��{6[��U�*��,nn���/tH���_�\��Ȳ4'C̃�m��n�k4��;� �0�����ǭ%o(o\' �g	S׎Ӷn�O���|7�����"�~�w=��e��o�"���jĥ��pƳiPt��-��=Y欤�۷��dtmp�-�ϭ�L�kZ��U�I'$��H�&�������r4������&㈭�d`4:~�w�(�� �C��j����X~�I��z�3M����kN�z��C�~0�WRL��0V�)�W�^�wI�X�V9g!�R�p�����S�k=����>N=�J��N�)���,�����%H���[2`��m��XW�Lk�u	�O$��P��҉��a��_�9!c�f����^�b>7M��'����'��g�z�q���B�Y�x�:�S�=V���^��t��n�]]�� /)�O�ՙ2��@]����*�8��~�_���g#��~�s�=�M�G0rD
�ie ���������7�N�Md$�LH�A�up�QE�@��BGވM)/Nt�Ev�f5��hL/��P���~�v������oK~Ϊ��[�S�c�^]��Tl��@�3��%�ۛ�x(�(.��j0�ja�5t���6Ē�F`���o$F�7����G���`�9n7�հ���z7��"(�T;�F[�t{���Hc��ڟͦ=Z��B1h��s}��	d
,n@��΢�K�is���sև��H(t���/,�����v�bV�Aİ�%eO0��7@�����6?ZY����=."a7�?�
��N?J�6²�x���-� b�rϗ9t�[���[���V���I�׆����?�b9���Gu=#&��mu�����{��h���׋��V�2��xƀ@뜻��=5P��|�F��[;	
�C�W�+�/'���M"dX bY�K*�������j�R��K��4
6Qk5�0F�� 2����������J
`iöd�A�Z~�7*)���W!�
`��t�Fb���.�����:��7}h��J��ӻ�CB������Tj���NX�p1�����	�]�z|�E�~'�������ɾ=�;IҜ��:3"������禐�/�JQ�+}i	jS���	�[�V6D�^��_�������f��[<����-U�g��x}S<!��3��d��,���)дG 
�!��]�R��7%葩�J�G�����:4�QW����t4<LC��v�R�aӡ��T�u�|
3|��%w�@��)?�[-�T�u��76>w��	ΐ�;'W�ޯN�8�6T2,�s`�Z��1/��,M�N�4Mu�.Q~��b��zǬ�5�<[�[�˦�p{���*�+�0MVo<�HAuZ�$��U0t�Ê��r����]��v����P��Q�%����l%��9�^��q"��;���
�X��v�F�Oy��#vs#s��?T&�C3���lA�����?�ddc�
�֦CȌ_b��x
Y�sΜ�c/\i�=t�K#0?W���ȅKG�%��T��0O������G�-U`kB=���ڞk�	��_�Tr\�h��]�$����&��+�i��ÒE��~!�|�`U�J�;���=���U�A����"�%}�,  ᇱ����Ѡ!i��B5���quѴ������y��7�#%��n�wL�a��2�Z�q�닛-��>��sp�a��&�S8X�lUn��Q��
�l=� j��Ʊ�Aa`���#60���f��n_X?������Ms��<t57���0���uR�L�~:c�zlB8�ڭm@U��LS��Y ���B����1O����%JkjL �<�Oư�ṕ���ꚾ�n0}�j���w{\O���M/Ni$76Gj4��مJ����}�|» �,�¥�tֈ8r������ʣ��D��6��j�/%���Fu�T:�"&��mT������ԣ�M�j2?��n+�j���0��~U���˺�#1�r�i�#8�2Y;]ń����a�%{j�tz�٘ry�jЄ*�����3�: ��.7�wV��/��¡��'��ۡ��ͫ���m��'���wj���[�e�P����$���w6��e	�²��q���O�'��#�T��R�(�	����Y�+�9%j�"����mBT�<�$P_-�]&t*d�Ѝ*h��W�r^_V������!z�f�n�IQ�}6��%��S!��^2Dk�F�H��B9Ǻ[G�so��+�_����ז��	P���D��O�E�TX��x=� �$��3Y��)�[=e�pZ��o8�A'���%{��E�S/=U�m���y4�u�ukj��s�á���y��q��B���ܜ�Q��:E]m�t�r��=�|�|�~�Ԗ��r/�S��V� B�p��6�%N�JO�U���b�G�s��DWƞ=�m��^=w�j�8���N��MW`��'������k���n��;S��-���Q�-�T��{Ȅ�e9�Gn�8�=Z�S���X]�8̗Òly<x Λ<���("���"H�7��q&�}<�"Ý|���#Ipڀ��1�V�G����=�w�����x{�cP�����;c!�����1�?B��pj��4q��O�|�b;���}T���[*�kJW�ѺL�pf=���%[�
RL�I�� 2C=��TP�s)6���l��������~�d~�W=����Eg���;�����U[�����LV]����F-�|��M�>�fDC�@�1 ����+�:�n�a����T���FЩ0z�	j�z�44K��CX4��0=�A��Dg��W�$��DO���t��b~��9���[|KKrMQ�2iTm{;H%���$�]]jP���SAv�x�\;��ҩW�f�[쉺T��u�>�-����
Y	e@�G������ Q|B�޹Q����b���Q�T֊�۴�X�4�CK��B^�S{�ϳ#qn�l�y�[;}ڒ��@x�n��?])� �y,7�Ы��H(�����مb�м.�Z��A�������&�����L>C(��Q�j17;���5,Zl��uw��y��g�:�!��q9��{�PD�?o�"�v[����FF�VT��E����d��?s���\�11�A��Q2�����_�i��&��,GÔZD��y�e�(O��'���/T�'�NX�=v�����t�ʠ2��ҪĄ[�w=�g,�if�u��l�Sh/��{��&e�#�]�"i�f^!��Q��s���!�xN��e�hE���Z\���t4�ǨL��;[No�p��S�h�s���6^��� ��Wy2;B��R��G�/ð������)�ez�vFz��vq�#-�N��ܺ�,�j48_>�>���� �ܭ/'7�'�i�I��$����|�BO3��S�'�#��&�w��rm����!et�kd\`��7^SC~����Y��s֨�kS{8�d�rW���X䔉Fw�`�������mk��nn����������N�=�P��!<��_�35�Q:FWx�=��'��܄-��/G�;���/6�I^�S��`�=_<��ݓ����m��j]�O���l��h�~��Xp胐j�F��U��n���7(����c#�����Gd-���t���?{����"�__E�N�Zٯ�^*���y
��˺���κ+�it����v�[��0A1�r6��j��-�~n��4Tw�fE��"O%%I�|�����?�Q	� ��2�
��n�7,%�Z��1�gu�Ҝ�������jn��?��,���B�����g�ܧɌ�)\�����^���ze�h��?؇��݇$�ǯ56݉h��W4a���dP�ډ K�k5�,i��R[f�b�@����m��d�R�@t������Å���W�y��^�.�������(x�����^�Le|"�ϙy���(\гI�w	�^��g@�jf��걓o:`f�I�M<�N�HL���S߬%^�%�9�X�á�'�]V ���X��!w ��1��Z��	�E���L�B%��,�����Z����1��*�͙5ѓ�Q:��U�D ~�e{+�"�7��r�g-d���� ��x]O&\��V!ݮ�UiI��Ǖ�*-�f��P��iZ���z嵐mt�hֶ�lv�v��.XW],�k��x���mj���ޟG�czBo���6�b����ۣ,¹�
�=�z�h��LkB,�S��Hd�s8�?G�I�%�i-l%M�Re���~�.��n�P%�s�Şp%;�J�(�Ј&�)�qX��f��ؽ�D�X�Բ3�ѯ_�'���3�Z�${��;��P�a@L�6%�*Ĳ��$�=�y��왡�#�����?;�4�@�zZ��UҪ��R;G*�S�F#�a<��UDܿ������+	����ז�#��q����~�M��J�H#�����&|�2����/x�,������8N��sb/F6���jAh;f�FHRP�[|����vX{c��`e��/gN�<��.����R7�ƺ� �˨9a�z�w�d΅"��Li�+�\u=��'�3�J(�jR]�̪+wD#�1(
�nL��(jD��A�%[�D�5����K0xoƩK���a�h�j�|:�f�vݹ���X��? ��&�ύBr,�l���t��=�5o�Y0����-����0|�n��g�O]�W��V�<m���&;�e�b
qG���.���E�ʳ̈́��ϼ+���-�lՂ�GA(��G�
��jfځp��#,p����΁|{���v`{��lƵ��^+ǡ۳�<����n�=[���AN�����V������w��`���!��9�N跬�Ar���),�@e �Fª�&���$��gҟ�PBJ� ����/��Y}L��;(!��iw���|���of��n�*Y��`B1����Ә-��~��V􆃨ʧ��U�����r.6uMӉtg\ο�
&���H8��;�s���ŏ�[L��Ӝ���⊏m�5��=ţFY|5�|>~��LX%�և�p��b'Gcb}Έf���g2"���E�ף]bF�%ĥqա��Ya�dej!����,�E%F��L&ݖ�Y�E�Hf�y)�jBD�c���"���7ǀ��^�"p�-а����=��v==ه�s\�7�����7��k����z��lK����Y̔�+�m��s~�w��^^���5�l�������8l_5}�� ��d��L'A*�w��E����?�H�����-�/�Ξ3�z��e�ɋ\\�n��{���fD�u):�!��y�>��Ʈ��	"��� *��ău�7��<:�(R٢�A�\O��{_5�VX�k&_?����6�X��	E;e�����S���ہ��^Mt�F'���ԩ�?䅸.�̴x�����d���k@�Ĥnk����P�!fЇ�xlC�r:��5z��]�%<,���^�&��z����Gh��ˈ�i�c�cL+�:�HJʙ��:{J�!�n�@�����@���
��?���"��Rۣtّ��X�p�����i�R��@{����X&̫���h��Y���ϞW��$:PL7��t����2.!�Y�f����S|6|�Z�W�h�y_���W��@���V�Uy0[��.l������G��rn�4 �R�Y�>��� N��f�?S*�����r�`�ȅ�^3��ts���vV�81)�t��s�ج����G!���i> םQ��.�`	n�~B!O-�p^ĊbayL#�N�WD�;uv���>d�xNe�I�Ѥ��2����hY��<<���J����Y�a�m��^�ҋ��/�-�Cqo��$�-�D�y@��E��X�ѲNzߕ�V(�z�X�ء���t��õ�+�o7K��y�Ёy3�yp_�L)n��BRT�B<-���'<^�i���MHh��p�j����
�D���� ���/���*z�&������gw��(�SE�X�*��Tax>_�?ɝF'���bM�b�<ߛ2�ĕ&Ac����vۙ���"�2KU���'�g���������)1�_� \�|����	6�>��kP��y;�}q��*��E]����پ;�h�ƀ�=ԟ�3E�k��L��Hۤ%^`�_�����0��R<�*��関�\dAԪ2+�k9�ʳ4[�X�0��+3Q8�c�>��L�1d�<Nl)6���b��=��LY=����܀��Rw����h�W��k �)1��\�te0(ڷ2t�m��m�Ϡ�n��&jGU�Y(^6���L@~���,G�-U�U�3`��M�D��Tq6�2�#�LJ�3�>b�s�d�T�����K�����=�BF�s�-dA��ʋzv��ry��C�h
@��]ڦ�6�V�6�{vA�r�����[�f�{}�ߊ�&mH�D��rW�7�
���[�O���e�lϭ�ڂ�-	iB���FZ��"�y�)?�]*�@Sn]�����h^j׎�����O�*
��⺧���u4a�*A�D����xzF��ӟ�b {1���lȘX����}K?���UB���9�����������sv��=�=���A���i�?��X�b�tC��3�f�A�� � ����"XX�����k/�/4O�K	����w��ҽ�[�H@k4~r�ɪ�L�#]wFRpD1�o���ǁe�`Ӗ'������3�Q����M��JyC�˟�=����@���v�ݦS�[���N�c������>5��D�%i���Ӷπ#�j��嬢��|�t���lSm�[Vن���:7����˩yH1.��y�=�F�-�hj��������+��UN���L�j��E_���;�k�r������v�c���-jX����:G�t5x~���.?;�6�Q�B�ӛl~	��ǚ]4�^bS~&��׆WV����at�SɟR�2�G4 ��LaH"�q�<��NR��\�j8��H���@eaK��L�|/��|^+^v�t�\����
�&}���E�؛r��\��ʍ��"��:�e�
�Z���#���-V'��N��M8w�����j��r�o���x5Om�>e;���f�cc�#_c/V�1~�UC
����i�R���ƌ!�v�ϛ��ۆexp$� ?��憋�)Tcq�]���Z'w�|�wZ�ERUe*v��� 疀+L�0�t,%��b�G*���0�`6Џ�H�N<��6��X�":k��%*1iL��w�;���R�H��u�U�1�Y=��I�F2	NY�rHp5ЦYg�p�vf���������� G!��s��>3���M`{̦Ë����`Xp�Bχ�O8��N���X�.���~k&T'�i�vM������C�a�L�R�<DM)U��'X�Є�1 �S�Yy�f��k`Y+m'f_;�<�F�(�Q����Z��PN� W��-�t��4*��&]}�J��co���2>)�>Tz(�B쨨�وuq��Y�J,�|�b�6g����Ҳ0浚R�ߞ馵�\����]�1��IF��1�ή\��|�,P�k���}��<W|��Fs�6�X�N�)�Q�f���_�0����2��F���%?S��~�@c�[8v]�ĬA;w�z$2H���לN�Nv���L]�C-REw��,��ۚP^,O����=og��c�h�@����K�����s�"�p�9�R���sp�M��,��,hnŬ�^3��fLP15�ˈt��@k\��߬Ug��r�+/=4�����3�3#�~ ��#g9�1Y������FH���H:���851�w)���v�Ƀ� �͎E�]	\Q�������q�R��cʟ���04@�Ӛ��9rC�m_ю��M����6̂YDb���O�Ŝ�:cJ�&���O8���OXX[�w���Y|�M1|Y��3!dTr����X�gˤ�=��Ol@�N}Yf����0~`�p�&𧶇{Cǁ�a��C5z����u�ݜ_�|5�Q���>'�k.\w�t���>Gԑ�(y[x�E���q�v"�J#ו/*�+$����z���h���XNq؀@y��1��ޢ��#�to���ڃ?�-綤�� �w�K7�Wlb��kf{gh���3�q�L��s8�bQ�zA�-J�aH����j���Gl���7��O�	��-l`؁�<ע���sz�}%���	������K��f��[Q��!T�g{���U�2���߹�4jyu���D�@���_�m���7�0�˵�a���8Э�4	�s'΀IB�O��7�jp���e�z��{��~����1�&h[�e�^ڪ�Z�!��)���-�+����kq�-�-��ֻ�H��˟�e6��(`a�; >���fFF:٘$Uj����R���}��X��i�f��+@����}�ǭ��^��-�wg��O�T �wa���$�I��6�>߉~�.�2�?v/�Brٌ���=��*�쩰���W��C����&U����Y��������(.�b��@� H��������: Zy=���EX8��,�ˠ�Wc�^�P��Ԙ
�dC��a� �B��1��꽸b|�W���ܻ�U�[Y�_K�����
΢�X������U�yV��ڏFpJ2t¼}�R��u�F���0G�I`�����^��&��
n���}�4f0	%kK��L�h�/��a��g}��:�Y �_$�^Z�)��D���{S�`���ݹ����~���Ϥ���v�fWuW�㺌IM,N�Q��ۡ�����`��w��e�m��☵�<B�ǟ�)u*~f[ĺ=����M]�g�JJ'��4��wc4g��:��2�YD��N�˷u1%Z�7d��gT�0⺓�|P  �\����E'-Sv9�H�ztr>�n�r� ~ըs��KR� ̏��_�����k#�"��B�v~�
">���-��NrW,�fָ�I�[�(�<��׋=<�W�BĵS�!�6�����k���'Z�16$��Ѳ���t_2����$F���@`0�	���,���.)Clۖ2���hT���B�!Ŧ5�}G~�� �'x�.Da�	��x����y�+(/�xL�@_)�������MI��o�\x�E��^p�*�"U.>:��lum58���O�]����S�Ň�]io�R��>�'֤a�E�y����=����q*8e��Ð�M�0	&��Wy�wٹӞQ�<�e��T3��lDlq닕�W�r�Y�	�i5��Q�vz�	vj5U�o)�jK����q*�����������[��^uҫ���7?.���(��e�4i:�r���z�˚w�e��<�_S�xe��{�
깾 ���ڏN��3p���nҘ�ܜ�{4҆K����d����R��k�9NYϬ�z5���Z��������t�#��`ôopt�z4KVA����6����կT�X@��< �V��_1��A6�d�P"4��.���'��Ok221�Ԥ�v�$O�
S�l��R���MH��)��:�1*�k�T�c���捯n'-���F=�kxÅ��ISӄ-��uZ��~�3��0�������-�<�-�:u�x�WFx��L�M0����6�d������1l0�8
H&�5�&���4ĳ�]�2���e�B�A�g�?��_=v2�|!Op�q���B�e0�G��$�Һ�UϞ�Nzp�>�'l0�8չSB�M��O�TD�G��6;�Gb�]A% 7Q~9�U�t.
E�ax*+y�r͗����g̕�΢�o��ˠ�t��������艁ճ󬬉���o7M*�&���u ���GɴP�Y��C��)�|� )1�D��ӈR��?l�=������D�Pk�"㝆R欇ϊ2�P�D���>��y`ˣy(i������5Kۙ�doy�Lp�����������2�M����1@w����)�nz5f�s��Ժ Ǵ+M�Y�(�����M���&�]���,*��� ��صS�^�^��<�����}���a��Q�!'�����9��4��֙��X�e�s}�C�6�k�+&��������Y!�l��_u�]ҭ�2��]�&�1��y����B���%NŢ{� @T�sHu����\-i�G���QIO��[�Hj��''�N�0�#���UőؽY�D�t����/<���t�ܷ=u��^i~işz�{s���c,>��ڼ�4�l�AT���R�a���`^L��:W���9�0��?��KĆw=�8�
�۴���a0��EM�߸�M�''��MO�?��Rƃ���>jp�_�EmH;�?����ط޳Jm���	��H����}`��ǣ�^�>S}ד�]26�����S�4��W?�C�����!X7D�������yz'���Ը�+1��gV+�вx��X��t}�8l0�h����ZČ3rcb�����D�f�����rX�9J�搞f	���H�U���]�:`��W�w�����M�n��6��`��S�� .*���#�YN!��D$��B�^����X��?t�E��a8�z�8f�7 �i;,��ugk��,z�$�0�.oCj�c)�Ǘ���e�sМt%/��y�Zԗ��I����L�;6H�9h����Ò`�ג�4�9�43l��!R$�@�h������3���0��~η�˺�*��ȶ �.5�
k8t}HA�!��0ðK�I����Z�RU����s�j��D����-C�����y9z�ds��Ð\��b�^[6���yiK�k�N�#Ϊu9����+�.n�L��=={|`^��hl��7�N�� ?8�*uh�m9GP�H����Z��p�� 7��u�Y�ع�P岂������hF��er�,WԬU_3�3��n�ԶEM?&0tS;��w�c5�V�8�+��*��ճ�?,��.`{RgN���
qFV��܁�P�Lo")^{�.��	Ĕ�*.��X�<��w�&[/§��_�+���h�F��=cȭy*�h�m���e5ֈ�<ڵٍ3����1���fng�pż��&Ru�O`��&���:� �}��ktV�\���kH�kkzM�[kZ�Ԓ��~6�Wȅ'_�X�r��.a�	�h��B�T5��]�4�$� ^�H��2�F�_LJ��ae�w�ih��$�M�f7r�H@�r$|���"��c�V�����2N5ǧ�&
���*1y�L�o�U������SNX$Ϙ1�ާk��&b��p����r
e]93P�/�%�"O����WE��k�z�A6~�'� s_vC��d�������N�0�%�옾v������m+4wd��Htu��=js����'�q�;�X3�B����b{;l�\��=�D��-��ƃ\t�ʾ";��6��������۹/=,�F�G�&���E�^<L��������2n��d����1���}���f����`�i� IG{&zr(>�. a�: �����<�;�l+�i���BzZt�&�?��|�(��l�9�/����jz9A�7���\�M@�k��s�*̡k����,�l5���>�D�Ҽ�D��˫��ω� W��@^l�֣���5)�+�Dŭ���^�)�AX�<��,�����y%�z+�k�;R,mn�P�}�C�8�_׌�(���vL�����R��n���b��-��g���!}�-�G��Lƨ��x��%K��#�8?0�d&�ʠ����ߺ7L�KЪ��>�L~�a����@���
��$?%����h�đ�ײu`Xpڇ$5#�7�h/��V�jF/eنЊ ��\�`����6j����jF�� �Ō��Q����/6Z��W��}����Q���WFM�42ej�a]��S�u��-Q��(�� �9�ha�~M�P��[�mؗC��#��Bk�X��^>|�����|�#z� ����kӞQ�-~��p�~�@�{�W�21ҟ���{a�>6�Pv��J-s��UU�S��]&�`�yWeq�\��ļ�42�)����C+*I��wW�#u�,#� �Z������L�J]p�̬�2���ZA��䅈Պ����S�8X�*)��I�����A
�䰖�xr|�V2\`����O#a��`uqQLE�<�E�����T�X���b��_+c�1��V��* 
� �z �<������?��ey���}~J����|�����Az��њK@��lLn��%?�����/,W�:����r�A��@�m�I-��#��i6'���R��f�� &J��{�v��PO��=���g��Y}!5�L�`��ce'�w���B7Y�q�����lS���w[�$#��b���)��7��U�S�u+���d�څG�^_�`4|NZ��L|	�Mc\����u����N���+�yT��X͌���AVn1��*��D�?��������`j^�좤��+z�Mŷ�מ5I��f����&]���'�\��Q�;

�A.��������Κ(��ay��ڵ'�>$����)�+�X3��B$`Bi�;z4�&lu���A��B/��>�˜!�]|�Ad-Qq�m�p*����fqN�1���T�;����f�G��m��]���8+�Ck�E�f2gu��V�]��bhKo
S	��],��6$g	F�W�2%0,�
X!g���
��H, ����)�H��Xħ	�w�i<��(�/��(y��%�?���;���H��+CB�w�?�$e��׷P^�9��4�w���Qe^4��hHkZ�x:��
��)���PѸ�j�zf+FU��x'�3KY�Y��\�p���v�a*נRQ����X�HpY�{"CNDMKBS"8�!��$֊�P'�� 1�f�kd���ނӎ�xxh,��nqnݗ�x�"��G3�폪��!������_\3��*�T:� S��6k
�H�O)P�x]_�ֵ�VF��:�+���;�]}�*'�H1g��u �#�>��oH��Z3_
��?O'�`n�YEkS&ta&�Xں����}�և
��?+���N��l<j�7�ۨ~Pn_�N�m	J�����:߇�be�������&�������ی�g��Q~2=q�Bt�Mo�+�㎦�/�m_���