��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_I
y��������k%̜S���9('�X�@�'�X��m+��G������g��d�:]�<'� F��-!�k(�M�u�=X͝c���/���A�l�8��'?nZ�]�,�u�������k��ᚘYڏ㑠ڲ]��L���s��F�N��o3KK�+^_o;�_3B���'���f��jI��j��ŪD����8��3֓��p�O�P�hD�����ץtT��Wp��ZӰ]1�b��#�A�H��,�n�ʫ�I|�_T#{i;��5�$mX��b�"�(���<�B��p�J�O"R���Cr�7몈K����r��K��ΐ*W�`� �s���2q���k1wA#���k�b>����8��0~XӋ�ub����?�\;VQ��!�o�U��u_3��7��"�o r��-�ڙ �j��}��q�4(��jbu�h�b)h:������d!$_���E��FH� �%��?�V��o��[M#ߕ�>*8N�5DIba��lm[����������)w�3����#Gk��y��~�*�s3��£�9�eC��>��U���.S���u�_��D��1#�����\'��v���O!��M�,$�* dM��Me쎶��ʧ<��p�9:�`��[5�^�`�e#5{���% [��Dnî�]���3^&�'���l�z�t3�B�Y�ׅ����r��Rc���O;#��#B�j�R�&@3|N'h���Jޒ�1��j���%�
�on�{�����}��.|"�R���BSaN�_+@_ʺ�����3��C�+T`�e� =9)L�#�~�n�s}y!�w��L��� !A�+__B4����u4��Zͩ��!����V�'C���2�	:wǺ�K1$%8J|�WG+c�"��ê^%s#���S���l���*�l�<WUy5~���j&��-����2�a��?X܌Ώs8���QM{�sO�A.3�g�������$9J�4��Dj� #��հR>��/ꋗ{$��~��3e�
۲������N��p-IN|�p�#\���,�h7Zx�¤G\�u�(y�Eb7����-��c���[���&v�8��s[��n�������-�=i6n18���hKrGҶ��
Xr�=:��[i���="͞w_0�jf Q_�a���K�g�	"��as��B0�v%6��
gƌ�ñ|@��m�N
Ga�YN�痣>M"�q�`�w��nr6؈N�����Dh�Ĳo
���6���F��@�[6w�=^�٬�@���#�'��X�1��{f5	��arv���Z���5�&1��9�j���ﺊ}���4��V� �.�����xyw������śƣ�Z�^<����y���.�
s�~����Z��&��u5�`:�룅hD���,���ܺt�ܰ��-��!�Lk�6]��G�!�밮F&�)6�Z�,�=�YE�[Tk7Y����:�����BJ6O�����m�zL\�Rk��T$����p��a��K�˱�H֙K|ߖ��Im�@�8����+!�K���
kD�Bկ�x�<�:כ�Rg��=5z�9�;VA�A����n��������/z����PT����X�v������	O�Z�e��J� �XHH��6��	&���+T}0>���}0�)�����S���{فvU`T�NfA��
G�N�D8�6n���&�yuNgd0��NE2J@��&NT%
+O2�1a7��_�����3�|��{J���qG"
��&�o��!�&��v���=�Đ����BR�f�����HW{݇\Zn8k8e�+jR1ڙᅰ�9�'a����S	y8��,_���ɫw~�8+�;�/:�ruZN�����f����cY��'�7D�{���1`|�v��L����e�����6"�xN���~�!O͹Ϯ�w�`�`}%�����?����zk�3�$�'���Kp����Y�����(��In�^!�F�k�ܯw��?��5�p�{�oFw�ǎ�h;�p��R�d6���͇���v��5����P���*W��b�3�I���/���9K&�4.�E���z��������p�!�1eU��z�Q�a��j���k���G�2LiG�O���[���~S��_m�G�Ѱ/n�55.sZ7�Öh�����?��m���WH���9r$W}����aqdH�h`W�D���dU�Z��̦a��EV�u����\x�����PK�t�L1�v;�X��&_�'j���
ݦP�H'�f�`~��NC�z-�;�Hc� 9'J髨�����ݚC�{��&���^�Zze�0�O�� �9�/g�t�	��n�(�h5T��m����4�V4��f�hrb�\��!Yh�A��S�&Ѽ��1h`�e���Eֶ�[�9�J|р�
�h������~߭�*1�WT'�_�^�M}�c͘E�Xޭ�Nt�5���c�`m�\�[Ln��]���ot+�&�-�\)'�،�M�^�� f@Ї���/�!芛�l+w�w��Ui�x���+* n���%��d%�1�07�~�7��h-qm�}}M�>p�>O��E�6����M ��e��
J�k!�*4��.���1M~{���0IC�*g3��kl_����l2��н��_{A�,Lf(�?���պ��CyC��z��3AI��P�0eU�]�3����hI[s�I�e��]3�D�ȋٿ�Z�c�ɏFk��B�^7���@#��@��fr4 �E���X���?��Fޯ��<%룃�U&�=o4H����H�������԰X]q� ��:�������ص��������ʃGџ�2��_�E#�`�ɬV� u\�n�Y!=({`f�-����F Ln����1��=_�,d>���"Hm��B\ktwy�Ym2j3ߪ'�]>ܷ�T-�l$c ��l��K�}u<�#a��|��(�Ym��M��H�1���m�ٱ��8%�;��2ս<}��6��EPj~v��?�U����D~�R=:���Ш����+ϛ䴍��nC#<���U���|U���K�ט��ب��Fx�a�����T,۶��OXy��E������\t����;�V������fKY�X:��� [�H�Ҍ�e�ȯ��o.��9����K�o)�%V$>���cfo�9Av��L^�!��/;v�B�{[S�m��
}�4!�Ӈ����z��3}���F�>���M����}�y�d��B� �D��z�,y�k���ǔ�E0�*����M�o���i��ƚ�`e^���t}�3�޴ܪ>�KQ��]������A$�*�c%�A�Ϯ&����@X͊���t�Qp=sA�&���5[�������f�&e��c��q�Hs1�S�e�=%�/ϙ��`R�P���h�r��]f~��\2,f3~ɓ����uH��55�ћ��� }�,
�(1����
Mz"�bNT<�c�p��L�Ù!��e��/�|�Ml1e��������?[� Nb �h)�{�3�6���+l2
y0%�W0'^�뿕�^i��M��[8	B���_�s�˛�N��<�p��a6��"YUP��,�7�M����D��Q�q3+��$����U�^�Q�V�H��=��M�9�"d�0�f=׌NK�W�.��:�A<���7����+Zb��0�Y�/�'�e��0p�3=fN�O�d��k���y /�$:��Ac>�Bt�i,���G�ù=G�Ĉ��_2p��!�j�z�,��N@W�ם�|O��@1�)�^ο��2Z�3���i�E�S#U��|l���N5޶ڎ��&�s�ܑҳ�ҟDs��D|��2%=��#�K����c��˅�ph5�ɍ����7 A��Y�IQ�G�'d_�]���5C4����ʹ���%���E�u4�^o1I�9^�����e���G)~�������F��j��!���^�֘��={�#�d}���^8����%�u�R]�9�i:��X�JGfL�?0��N�{����q-��mt�UK����-U�q������U%6n�vI�X�,�o7��>���[Ā�T5B�T�����@�:Z[�5�S�(�ai���}�r�E��C6�&z4�21��dq���n(̓��&���A�Bj��O�9�ӽ��q�p�Ҡa�n���g`�J��{��$�C�>�[�W����_}%��S"��A�l�M�{��@���B��n�2?��й �"��W������1���|L�Pú0Y&�����;��<^�;��(0��ʭ	hn58�Y���P� �h;�a��P��ާ�8���l�w)K��y��|}WHMCQ3�""�W�R����{�4{<�!Ļ�F�7��`����E�l�Ώ����Y|���
3��^��(G�Mu���1�!QB\�)Z.�\U�W��і"4���nҘ�H��p`����/;|�lهܾz�]	�����%ʍy��
��vJʐ:y�"��[�&ܜ�����Q�n��a�<�m:d"�������c��f��^٣d9AA��A�w�D5��ނ�����Yp��B�X*"'�P��`�zX���� �_���s�w�*z����K��9j�
Թ�Z�uvBj�y��v>�RUvԟ.���
W���^�y���938[z��x��-m���B�9�5v��R�_y|Ɠ2^����/��n&/tL�g���e��q��S�#01���Q�TBȃX�>j� �'�0�'`��;H����ٖ�7�������8���H!u8?J�9����D�|<)�iA���ø���|�b�q�h�H%��l�� 
�r�6�D\�ɋ\�|bý	]�Y�p�)o<S��9Ox�6_�
T|����	�M��¥��b�)�2��`GD:����+�7��|�lA�����0��dh���"8�>�D t_��)�����۪�dh�6�WD�J3��7#�$\��[g��s������@���y)���?��#�NgZ��	]�| L��Y`�fw
|��#�~n�S����(h?TWg�P����t�9����Fw^�����)]�R���$%,P*���Xت�������A���H���%'ht�4!���9"$�pR�/H�|����J�[]J�H�
��r�L|��B�)1��z6�$'����U�M�*��K,6 ���G�a9���j3��.f�[�������P��$"�P��(s�j\=�gFv�^�l�G�;��1�kw7��OD��VI�͗���+��Z.Q�8r�"v�-���c%~g����G��Zv��z����iK�y���-����V�*�E��I�I�y�w�����}i��R~�(����d����ڬ�G���|1S7�{���6�2_Y<��▂������a&�=�u�����? 	\�������.C�������#��{�5ƴ�C�����u�2>Սs�WCn9���O�ɓ�	�"^�!&����^�BehmJ}6���w�߬�h~>��o-�c�A�3bn��9���(��i<"dt��3�&�}�L��0l���f]e�dby��~^t��.��?�WK���P�5=3�:�Y���kv�^�
K�D����t�m�2��������}_	+&YY:�q~��ݟ�W��0.�Z}G���<��I���@@}��w��7bH���'���L6uf�♽�Qw��%u%�Q��k��v��J��nF�X�N��џi�c��n���++��Cs��A!lK���c��|	]A�����E�ic �I�m�l�?��-Ev=����,H����S�|	����w���@��s:�1�����3w;�m�F���#fbIdբTgQtT���p\&)�kj�-�v�7�%M�@R���.F���KJ�����aGtLx3f�D�;�d1H��Z�Fz�V=s����7=�ž_S|�����5�?����������'z�hRɃj���`�j�و��/x��-�E+����ȵR���>y�i�6$_Nǫ�s(�����/� <v���Mõ��vy���9%J�J ��I
*���s���^-�%�nq��,;��-Ƭي*=R��y����o�I��	�2��Z�����c�E������{P:�� �p���M8 X�q3q�Q!�{�>�k�h��p6�,�!�3n�(�6`�>�j�;���)Lᅱ��ܫz4lY��_��|��t,�^�:��`���D���ȀCka�'NN��� �?���S��͈�C�՗m�i��%�>^���w��*��,�/��xw�N�;u<���n�t]�i|���S�v�8��1���i��@�tUs�Ó�?�X��:A�rH�(d��o�m�*x��w5t�>���~���q���]ג���8���đ�s�VK��F8Q�N����8�V�5�n4��u�`��}�*^r�ns����^������V3�C}�G�T_M
�ҿWj���8U�Z�%�D�V�(i��P'��\w%�
[����Z7S_��=�?��	�v��dj�D�*� |!�eN���_���W*�t�7�Aǽ�8ʙ�����ĕ?b�T<�VZ�����1��]A��/=cw4-�jR���n�;��W��p���Ѳ��Ϛ�Oi�*UӤ5��r��{���
s�&��zNʗv9����=�X���γrfS��̌ޓ�ܰR�
T}��
[��*��M�辰 jX��a=�=0�ҥ�׹b��2C�:��g�:�I��vp/�V�%���.{�O����ǟ|���.�*L�;�!]�5<�[I3;޴~e��_*�}CT6�&@^�xب�A>&���]��s"����a� ��$�ޟ+n��ZG�Ee7��*� $��w&�_O����J����Bv�f�3������20��l���;6�8�v�v�5?ԑ��|���%�L{��g��Dd|!��D߁��&<=��<�p>²f�1K�/	݀���G'�:�G}lE>�ֱV
j��� /�DV0g�Q�����O�I�O���0�y�z�L�k��Zӏ���i*�=�Q��줲Uv����6!�1�G���`��9F��K�.g 0���p_ZC�-���$��_o���3'.l!s�^�߫�+`�9�����/˄K7\�F�'E+�d4M���W�U+^��nd�=�Ә���(�~�-�)���;���r��Z��7�������`�'�F������Av]����VKh��]=�	^ú�K������zb�o���2��gZ�7���	]������C����F���~�.���v�t�ZHkDjA=����#�dG�Ԟ�؊��u�[Y�0����4�����i���������Z����ի<y�'�����=�����V�c���dQ��3�k���Ѳg�#��ԥKb�i�����f`���V)%N.��O����Z�"����Jk���m�N�������ʤ���-|���c2��n�J� ����Kq��q��CU��k}���_0}�$���q�FP�*5��xe������8٩��|�s V�2He�|x�O�?�S��dw�ʤg7I����sa T��U΋:�Nύ�L�֖�t�P����a$hQwG�1�+t��٘�k�0������� �@������n�M����\q�H��H��m�zK�L���Hf�Bғ �\P�@+�?�v�]�����"o0�<�Ы�_b_��a���5ۈ�R�����^.%���I�,�5`w�"�>.��c,qE4_NM�'vˊ��~ν�@>�2�\[�|������_��n	wy�:Z&�s�=��\�����m׳���:@l�_��q�PMר�P�s
V	�E��^c�x�~��Ⴧ�b���?����eV �Z��`�q������*���-��%V2ǚ �G�������P�Ԙ���H�Y��!/�����,<r��<��b��q9����+����d������x�?)�)�0s��+�HO��ndUy�?��0$x��eC���q��%�D��&�P�[�+�/潕��:e#��/�񏍤+�㬄�b){��u8L{��)��	�r�	�+�6/��D���Eʢ���G~	�s���i=7�⪙�Y���� n�G����Ot6���}��5Z���D��,k��t�y�pK��h�:�mh�xO�B�v���x�-y<S�ijⶃ.67����E=�\@~���Y-�Tҭ��$��#���&��Q>D@���#��WҸ/�M�+��u�3t���\RH���� KHuÝ����	|�2���;���M8&=�?��I�u��5:�n�H���x���z*ykw~�E����ډ@ww1���PGњ����R���&�OnyAM�C���۴7}Qa������dnKV�"�
,,�X�W�1� �#e�Ko�$R5�,��z�D�v+�D��Q�~i��v�k6ҁ\ܹ��!Y7P�S�Z�޾������{Z��ŷ����8Q�\�8�EƁqQ������=c<ͼ2�!�YvG�2�[���cgy�Hb�Ѱ�7f�����^�_c�7�j��0 Y��5���j�" t��*�-���^&���i$J��/�չ�C��!��OU������R"���%l�Ϥ?| ���Bk�	��V��-h2ͤ���dN��)Xh[�７�G��z[o�0C�R�a:P�Q�YF1��N�"N��GQZ�>�� 3�	�\s��C�����'����r�Z永En�������A�:�㵅� �)4�������F�a�bncBY�� �C�)���x��pBX���H�U;��1-��Ƞ֑�ql}�L܋�<��xO{Ҽ`�L}���hD�o����y�y�\n�e1X;�A�^�;i�sQ� ��-����'j�wT��Ȱ�}�%e�fX��t��@�n� ���_f�O��|��!� "��J�����ǀ�	'�_t��@�N�hO�
�C��n8*��HG���x ץQ@��OKc?�����8�ڳ�k�g���� ��?'�<�:2G�2^$����c`qs?#����U�_w}�R$ϫ�i��9�9=!?��+��+�#��Y���&/�|vZ����J�)	���\�����%�G�p�m�`�a�P�� ����邙��fá��S�N53�[k��>?�h+%�l� �����#ə4�7��w�9oa3q�7m>q�u��°؏���ڹ�;?�kE��
	-q"����,�W�5n̈́<je�z��w���bv�rƝ���3E�gܚ�O������{#�	|�L����&����Z�����+��k�`����o��k4�Ѻ䠦�i����y��C��zvm�-Bį�'Sr��f]S�1��ǠD�0��\<��k�rr�&�	1Q�!A6bK��#�o��t��T��D\�z
O9