��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K��R�9��Y�%�itCy�k"l|�.���n�g�����P�������57`�����#K/	�����>&���$���;j����Z�4���.S-���8/xa�Pw���1)~���l�O�hqO�y�2��=w�'���$�j5~O��#��rMGeXG�NN뭣�M�Nu^��k͐��}����%t%���8�g��p0�g�DDXirPNv��G��U}*�Ǿ��b[GSg��f��3+����^Xs���a͓s�55�[�j��5Q����d��~ц
[�]���e������&#9ۊ��g�7uЦ�׸�!Gr��Uh�كϏ��9�m0Lŕ8��[�D��D�u�h�ۺ=�YF��s�=C����h�����<���U���	 ���au G�'C$������*YD����� �re9�ia&��*�U�1mbʰ�q�^��8łE	��-��Q���:G�}��(*�
�9�><�`>A���"��2f�����o��
q� &`7���n�h�i�ک��Xa_������#��0�����I�� �y�H�[��}�e|T���Y@O9!8r��g
D`�K��^/`͟�g�ݽ�rZ��p/�H���5X@v�Zpqfo��W�M ���	$����:Ǒ�EP�S���^�8��I�wz׏=s��
}�Q]��̮�$�+T�����դ/�G#���$Z�2��d�'�G}&�RK�a����FF��u���kK\�ZSa>�;: Lq��_h\OբX+vc(��Sm�Y�9�o���z�!ʹ�ͪ�p}�OCC ��yJ6.�D%zM��������
�{{��ӓ.�"c@P���Iy�-�N.E3�	U����'�E�9��mp�g楉?�a�$(��c�Eo��!�OVٺ>�a��.�~�F�QӞ.@z"�K��~����[Ǹ�9��Tu9&n��M`epׄg(A���:wK��W��5k��#�\��IʭTD;� ��Zu����Z��q�Sg{.��qj��K �cǩ�Z�O���/x_E(X`t��p-�D�=�nT�1D���*-�4A5�+�s���6j�U"a���A4�w鑅�f����xB-��+X�D��,�5��3��;�l�rf�Ŭ�����.�� 4���[�t�0���*��i���
-��i�x��c*㾕��y�p����oL����`Ϳ̳v�nQ����-�$AX�{FCW0�:$����@%z:��0~)K�ݯhw����
S��'�T^� -z�0��Z�uXWW%"��_��;1VO���� �ݤ�t#'�@[a�ŗ��܅�d4�<$��~�_�aҕ���@��n}`}l���[��O{<�*i�8�AS��<}���7.(��\�J�Y.�V��Z��@'_Nw��e�<r�V�I���~�~ѳ31�T�h]���Q:��p��U�m����R�y�����C:icPKŀ�;��l�|�nͼQ�rV��S�Kn@��Fzha�Ǡ�	�so�˼�!�L���z�а�;ذ����?
}�ge��&m^xx�)8~O���ا��T���<ϫ�w�cOd�ž�s��gKY��{Ԓc�l��M�f�2T��0����
$�IP��iv�c�1ūA�2�Oeq����՞Z�A���5�����O;	)J�*��7޼o<5�����O41oC��H��X�n1��̭(m4���I�y���A�ەС��雽pPK��YA�3m{A!{S](��rN���*��0BQ��bg
�l���b�׾�W� �A�9���T��~�p'ԓ$��OMe���,�UJx��- ��g_�󅓔F�4sF̗l���ED�zUT�o��t�xLǡ������33��N)�	�+�����s� ��6�v��v�W�O���KuQ!���}]�¿��ny�A/}*N.�3���I�Q�G�3��;�&�[��A �'g��>YG�W++���=h"ZU��zɂ�<��L�$��-~�P9�(���!kTj��)��Epj�V{J�?��]�����Y-b);�
]"�n��[9��>l���gL��א ��]|+N�/���Q�,�i9�ME~�#�\zYͬ.
�q�����ŢW;B��C�*.�ۦB� ���W�g�`�ƭ?��'J�F��5�!>Qd5����n�&�.࡭��V�£\?+ ���nlǏX���]0d����2񐣹m�g���UL���2��p�'�* ���녈D���ۀ����.�A=��1�g�s�{DF�@�y�@~�0�0es2ػf:%"S�i8u��k%ۼ��5"\`����_+���_���I���I����!|��r��q�qN�Û/��F������
���'���q�����
�4|(8�a7%W���K�U�b�@�k�MP��r�Y�󿝁_#c�o��ߴ�Z�b���AA��\��揦�Z�s���U��~�XB�ˏL��m^d�`�kL��-Qq��d�}8r�Z�c�Ɓ��*�M�\��f�=�G�����'/�ɨ�Pw L�jF�I�
��u3 ����8��-���ś~��p}؊���S�I�v�œ��6�> /�r/�8�J1䘃h��Xb󽮥�d�X�����]ó���� ����	Iؗ�)I����`P��C-]��w�f-��{������L+�3����NX�NwI��QH���[֐�n�M&�ɰ��s��V��h������>{�>���^�P�!���U�����]E��I����W�����w�ېt[jV������2�@�s�N��v2IV'ǿ���#���Bct���",FZ��u�dC`W�|Ͼ�Q�tRr1if�<�O���>8� �K�)���M�=\�atټ��,����m{��[x�ڞ����ɿ%a�SA5<dو?9���H}�W�c������j^ ��%ą����ʋ]��$��b[�`��W��"3M��j�����@��L���n@�������L�m�������H��^<�s󻪂��@��f�1Z������z�`�n�}vkfއ�Ҋ�����fBG_4�@�z�����BTk��v���AiG�D�@YN�l�.�G~P��*6�ɾ�͐�fg�@U'���z�R~dF�C�s�Y����|ޏo����@�(�F���,3�b�X6�3(J<��E;_��Y�{�k�bF�ܺ���;s����uSJ�$&<���{�g
��B4q��F���z����6��+݄r>�V��7GX�� �s?��8ځ����"�\"��JZ_�'d�e3����zK" 9o'�lU��M8N��֦	��-����.��*5���ڸ:븙IɁ��M��.
,}&衇ۂP��1+��;�X�T�����wm��L�p���9l~�6��E_5~d�(��S�w�,n����3�k;yV�ri��N,��G�&Ԗ�.�źZ�?���{Z/ǶA�T_��y��"�gi������Y�*�^Q���qۤz4��2lqs�.�<�,���_l��E�w맂NAͥ\6g��	0��B!j��K~�����yQ�Aqi�į,u�G�$��@�vص�*�g����ud7�����"�u�'`���#7�@�XQѹ� #�G98��'"0���nc���tΠ-3�+S���w���Y�`�Ѥ��L���bJn1�8b�	���(m�[1q�L+�`o��x�
2��aǈ�j���Y56���`#���1�3 ����	��j�+M�ȭ�� 0���qI��]��%��A�3b�����@ti�Y�y2�ڑ�+�%�1�x˃��;>�b�a6y�6���"���nn|�����k/���F۲���}ɴ�3��[!/��(���U��n��G��k�Ȟ�M�Ca�-m� ���n�������8�A�j��Η���/�=�cH���<�"�+�7J��6#>�`k*�(Ax�Y�|�\+���$>1������/������S��&����{;%��Y�!b�� y�1�(���si ��N/��ӷ@L�j����*1l��^��z�s/����F~��a�6aL�Z��`�w-�mc�U��� 鳻tĉ�7ra�\��eۘ��_�����)z�ܟs�LBD{VW��N}�q�ȹ�+�r4ʏ���8�4���h���`�_	��Lv��;��^��� ���^�`~ ;�ޱ�D$;E]U�?����/��u��8ӌ�:`҈"��{�!o_��ob�o�Y��wI^�X�ېO8�a`���i�hR��7��
.�(W�߄B�&cOCq� a;}����2JK��?lBjA���ʲ&s���4;4r��t�S���8d��U��B�Zq�P /����	<x�a�UE�<C�,�����I!dNq�\�-��𶩞��Ǜ|���6���{Pu�AX��l
 .7�=񰆣k*�*E�)��|vGϓjS!ґ�w��q���!cB��w��� mّ�W(H� 	/�Ǿ���F�U'�w0|��n�!�o~�Q�D��O�-M��h�H�J)���)�V�E7�3�H�T@��r8�n��:�!K���͹�a2՝�j�[��3���Mao{�h�|�$*sHEa�u���`,��lq~x�(u�������ʥ��*:���Cdo?HF�y�5�݅@�h�(`���&[q�k�]tlS�Ā��bw�8���P+�D�S'�pR�0���HҥI���;8��?��CgP?�S ¦�_-H*��5��gh�d?^�w\Da�k�����*�&w���M� �#mi?H^�D��گ	�@3�Y���:�
�L#$�L�x*NY������E�}��l\7Eb���?W�8��J����֗-�l6#E]u"FCae�=���>�:������c�GHAm�-^
zq޶�q�8�����Q�m�H h���-�;S*#�ѨH+$�]u��\�{�����|
�'���|D<<R�{ak���'���%�CR�<�~
ȁ���6���m<�
g�_j0|��iĄ�A&�~�~GQ1��#�k�)��,�lC`�\�����K��>,��~�����a#q�#��Ad�/O�؇�o<~��W�41�����Y-�K�j�V
����n���._��E�9 [-��]җ[P���ꚢ�o����y��,�v�X�^֗��-�7��wT��B