��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_��~�og��B-��e�g[���$�Ԃ���#֩�&l��=�̣
����^�����l�l�>������q�9�J�1��u��t�l1OV�kQ�`w�!�"@F�]Z�/rf,��l �[�~ĳ�&
��e-��/�S�¢}�/Xq��I������Y����K܋RH�LF�GZ�9X^V̋A��N: �\F�?�'e��jK0B�·I�q����~/��WuŮ	�L�M�}\�@�9�!Xe��|b�7)t@@�s�+2�d����^�����
-F�й#S&��Y�5|E�;���|W�8/D���4v������X��!a��J .�ym+�3��wM�PD;����k���O�2��z��-��r���Ά«���<����� �Vos�QG"�%q��W}��%΋q1"]��,	qbg���.��zw���C]�YMΎA^@��N�ٸ���r�8��v^�'dݮ��e�Az����S}R��tܫ-X�r�ň\!+�j[+=���톸��45�^%��c�7ZW���dӟ�;}�t�B&!A�˘^`"R�̈́�S��u�>%ȿ��b��l�J݈�e�HI��.������o�m#v�͓���i�&^y�c@�FO�e�Ѹ����BG��=F7�7��.W�F�?Z�(s��=��Y�ȣ<Er��tP�b��4��t>���3ҭK��&�*�.x����$���&!��A����� f�z�c��D�{�ɕm�;;����}���C�`2�G���W�	펝�A��������Ȩ�VR�<립�J�����u��:�6��x�فaQ`��ؔ�b��&�v����lC�{�����1q�5�G%u����D����\f.���W�r��H���+8�,V9�^B�Ï�	��-��?��6�+S����k�
��a��Ć1��l{˭з�l�UG�TuM_�'��O>K�`�+B���Ml��W��º5�i�QPT�t��z}\μ�����d��ᙳS��ɭtr�qc7����C�}�e~�r1��%�*���
�d@U{~��C�swLaXP�̩�@*�����`����*�O���0���)K�(��-++)9�>���wH�ˊ���J5�r}���ⷢ�}`��m�ăR�����,�k&��y��"�x��/-60eT�Ci���]�-ʖ��Z�&?�eTSy��QD^�a��M��a����I�������;��6� �/7TjTv�B��	o���-Tp+h�"k���pwv/�C��{��8�
�V���<O,'���Y�Mj��硶�/�hy9�[j�pǞ���an����P���>�=�(��s2��A�y;�Ir <��d��<�}�|*=�hr�n�n�.5�5���04<~ٳ�>tֳ����ʼa�՗&P�I�*ou�z@v^��}^��T/�Xc6�@G�ө5��t�G;�����.zś��E�S��W#�X���Naw��Z�[*R�ǜ�����/����1�K(�����l�:j��۬몒��%#�8�Awʈ��z-�Y!WJ�D]6�kz��'�SLnݤ��o/��/���89��J�6�6�`��]#GY;1u�H�|�k���3LQ�M��D�U���a�wT�C�uPq��Y\.�':��eہ(��0]&���3Rp���]�m���	���Z�j=n;<���&������`����Q0��%��$�n%Z�d���	�YN�_)7h�|���V��f�I^��RVѶ�Eh C��3Z�w�Dr_zՆ�	��E�o 8Ũ[�⥑�+�	�	T������s����H���$�,o7,���]a�68nJ��l�oUi
2�I��:?<�G�c�v��VܲhǊ��>o�I.�R��Sd�>������f�{�@�1�Y�������%�y��,�*�P*���nF����N�6��y07E���� \;Ɣ�,����� �W �l�)y�9�z�AZ�L�5��ԯEe�~�*'.;rL������J�$�Iib�b��5΢-�4���@�4��j�{X��4`}n�~�@�h��uM���|��YRf�w,.�!��S�:A�:µn:uU�80�I�(C�[�	���))��o�n"��m�#����~��4wP��W�w�%$��N��Km��gz���0?2Xάݥ��>�y�o�_�2B��x�����fj%D �I0���Q��V<�!�e�C��7��Q�|�'`s��Q��pǺއ�i�s�Aƶ�5�������[�
����^&j���[,��u3n�D�|r}8�y���P����K��p�d�-t����>~6��["y_�z�X���]���
�P%5�>7B��zͣ�û�����' �z�]o/⸜i�������]l?nѤ�H��G��`�l��1:?���i�!��2�o��^ݒ�B0$1|ea|Cā:b ������h�s��~�LJ(��RS	���hB�?� �����M�^E�heh�<�A�����)?"��6n�|o��X���t���
�C��$_GIWiUK׌�'\.!iA����S�tH$g�>�ֺ�˽���g}}��XL�bՑT��*%�$|S��tSC5�.�-��̟|=�jb{���?^��0~�i�#�4@vd�X��&?�>Z�l��K�C �*���.NN0kY����zȗӨh�E6`���f��i�����]�餻��S�i��zH`�S�<Db��U7��T�Gh�i��lf��׶<�����\�R�􂥷�f���[ft�:�;lo͠^�K���/l@�؅u���!�m��y{����w�����
P�o�vB�5H	�#ՠj";���å�a6�U�B(��d�Ri���V�Zp�Z10�n�rQI��biהּ�(?�Ԃ;����' /��4HD��x���5�}5lL�e4��J��´T�M�vôbwR��=���fw������]�2^=-t���=���K��DIӶ6GԝP$����t�ц�@ ��>�E���h|�9����t>S�-n�i���j���,;��.��<�[њ��D��:~�GM�@z �/��4�p���\׷k3��t��#/cjs^�c��l�.�4b�B�!j4��̢K����Q!' I���W��)��Y�
>��Y�}=�R͊�Q,�Ǹ	����3_۸p��F����I�s��O#0�Qz�U�x���Q���$hdZhS�u�&u�V����Ŀ]w������r܊	�p�"k�Q4���ηKL���<�Z2A [��V5���e���R�`�&�X�D�8L���e����R��o��5��Ɍ8�#�ʄ�ؑ�]
�"s���j�p��ED3R@K?s�������h��
%"e _��I�$���Nu-Do"�n���:�?)��^N�����݌yj�1pRG�*�P�ӏ�7�9U}�T�v�}Bq����	�ڸa}??Db�nBu��{���'���0p���O���}�4��|�P'a\>�D�Ja?إ��h ��%`:3L��/+w!"��q$���Z����n.L.@��T�Xq]��~�������ѝ��k�h�(̓���=}��#�r��Q�E�~�]E�$5�J�A���*��ӥ��z�b�GƂ��՘����1�kک�=�CYS�$4k"��*_�R�hH��%;���O���V�M.GP�@K����eݽ���	Z�w$��b}�	kv����5�ѧx�kp�,�|�)��]���e��խi�t� �V�b�S�*���ک��cU���-J�.f��#���V� �l��j�^J�����HJHO<�����������j&�b��R�ս�5pAD�G�8ix{�̫�A
��<	�,�To�/��o򬧐�p{R�d`�'��H2ŗ�&'��v ,�����?Y�Ϩ	 �Rt�z��&>�&$����f� ���j�wTn�;�9��<� �L<���=Np�$j�f�U#�:m>Y>]���/"�a�H���U�B�}]��	F@����r�ֺ������9\���E�j�|>���!�v��>)}B��ś���(rhu�p�O��S� ���go�?{Q�(]�i:�X\�&�x�W���
�.�%F�{$$��]7ٛ3�zB�'� r}-_IK��	�" 4F�`x~�7�B�;��=~���9��;�!/��)��u�`Iɣ@K�x�O�O���7S�Qr���k7��y C��Γ54X�ꝳ_q�CYZ8�ϥP�,��7X�����Yq_�{s��g�v���)7_�9#=�ؚ�kI�]������U�B�n�����LCS�ϳ4�Zƌ�^��7�[��LVҰ</��F���snG�޴��O��yu��꿤Z{�m�sz~�,fj:�-W��@ӑ�b�m7D�ӓ�k��m���Bΐ��B�[�.j{�j-����|�7(�%�t2ȎKv0����BΣV��,���iͻ�Y�����..�N�� ЎPC�N�iHen�)a)+sa��J��CO�]`a)�Z�g���vC�b���Z�a�?������Vmk b�o��cr	���Î�E�@�.	Cpn�#f�.�:�\QA�'�^@S����|���g|�	�Ys�n�i��H��.7H@�Z�%fmV�z��{�����p�e�#D�}�kC��mJ���,٧���T^���$ ���j�?:����ш�T��ܺ��*��/ͫD�w=��~͑IQ�'QXO3������]�
�1|�$n+�`֊=���#��O�,��@�,=ҫ�	��L�)�ha��ܜ��*�O؂Ooy���Bt͐U
ӡϞ)Ufl�G!��JI�D˺ePܪ��=�XGr�E�&tz�7�T�{,m�
��q��*��2�6CqU;u�R�ſ//~����Q�#�E���oY �1I'M+.ֲׁ�?���-��^!,$oqC�%�C9�%m`�}�n3��������l�����ϊ�U�ݢ�v���L@$�6���;��J9Ni��RV[U��2����h,bNwj͚�W��S��/�[-b�U���o�LX����Ra6��We�Ċ�!M[��S՞�%�;4v���Ӿy��{t�/-��,���>�@��^ֽ�u��'s�+�~�>#����0?�8���T(�D�ʌHjy���۞ώ��~R�����R��2�
C�?�{���"�629��{�~�p.�&���,Ad�Ȁ�!�)��Ҩ$H�(�9|�����,�R]��Z�PVH^��c�A�fO�F�Y�s�iж��tٲͤ )�%�f;����(�%�JR_��e�����XM �cBL�D>ߺ7�(��v��{��N4ż�x��(�+��8?]G��Mf��_Y������o�{��K{�5������'�=�ҿ <�U3�p H��D�L��_R<ʮ�D��(R'J���=׺��B�X�#�����O4�
`�	-���h-��������y��"Ŧ|#�=�IԔ�ز۾4���z{90;DVS�{ջ�T@�-S�y�C
���#�µM<�:��{���(zz*j�f;wn"�1]l&��XT��������%"6�ᨍ��K?����b�M�G-ͧ�񃔷)m$B�'�CeX]�4l��G��B�<(N	���j|�m�3���C��*�mڹ���s}+Ч>\�v�!�ئ���M�Q����7��:Ot�0(������6,��A�{�|N���d�7�FSQ���h����``��R�'��trx#&I�!z�'��ޅ��T�����9������ؖ\/���.��ea6.��Ի��.��3Sb�.B�>������8�L�LR�����e�2���/2r�n|7��Y�g��Ry�����ܔ�/^r�$LH�D�鏂)�F-�� ��AL�!]�#/��Ui/jҰ��(^jU�Ư3Ct�`�u�FZ����	�4F7Ǭ�@=&�|ˢЩ��n�f�Leþt1�'��)�`�����9��[$��[��� c�E:�4Ե�P�PT}�hq�|t]��~;+�q���i^{,�F�������nˌ���r���D�{Ꟗ��B
��c�_ZOmn�� C��1@��3������5�0��K�����}i���A-Ea_juccԾ�K(�-61��O��!|G d���ifx�֣�	ӧ<�+	�L�)�'�.|h�W<'uS��ڙ̒�
;Q\�\#�ux��X�dq��N�{�"EЫ� �A��� ��ߌN����[�XJ2���\�r���$\�9s0}x)B�RF��j�H9� �G�%��\��܁�e���p���b��[�AF���ˏ��",�K�^)��
�}+���c����JO>�(Q��>n�{`�4Ő�!�9��B�@�K�̕�hyN��@��=E��_�8)C��hT�8��~9�q�6�g�|?Ҧ?��� �@��w�}���x��8�є��t�(��W��ī��(f/�(��#�l�4�i\8e&��R���:�Ѣm�$�>�5��p��D�,� ���,h8P��c�+d�L���A�t��_S����G �"�ʇ�f�Xj
�A9�MD��"D���H$�Li�Rf ��k$&w��Ԗ�:b��/^�'[l"S0�%7o��!�h>�-9�0*��(��9zyi�S	�J?��Z>J�'��w��Ғ�u�2F��DQ�$a�6���YF3C�Xλë��b�V����wG��R��}i9*Dt��	��8ò��ժ�q�c8T+^0���T#!C���'?�7��J8v�(Y�����ډ՝b����pQ0���U{�!�RŊ%�^k-io��ջI+���i�3�j=��ӯ-:�胙���i�?�%�bv��\�/))&�&��#3v(@�z�A�Ztl�Q7Ӎ�MN��N�U�W��;�Lz�^��I	��i�NY��س��|l*ɻ35����.���q� ��í�g{?"7V1a�^�q�ܡ�C�zS�����t�lzy���0��;������J������z���ٲ 5��G���-��Y�����&����Wg�����/��|Bl�U���b6����k�xRQS�޹/��2y�8�_�:�+�8c@�m)��Ga��ou*Eu(Z�tMa���yS7�sr�9�b�+l�Il�3��S=��'�
�[l��;�8i�s�YD�����㉭Z���� ��x�J^�n��C��Ӂ�x:�OU���5���6��=��xY</3-K���wدh@k��F d|�Q�ؕ��i�}���vk(��9����m`䩟 �,H�����;.2����i�$v�@��5٭N�*�o�N>)O����c�(Ɍ	�ç��4��~���h�^y��\��<I]�E�%�Dz�\8�x���P�r��I�E&�{�,��E���[61�&u�x���Z����,��w�%K]�����ך�M+_%k�z��#��$e�d"N����\���c�Ȣ����8� cM�d��c��( U'���3���T��-�xpP9�kM������N
�L��*_�$b�!3Z�6����`쇑<i�O�h�-��o�q彠ĨM�l?NԽj�L����r�_a��?�Ʌ�$>� |�����Y��MלnШ�M�Y,D���T6�F�h��w-��ؓI��ck�Jl��k����u�t���L\u���@�)���U�� H���V���mD�E�f�}@���f���;��3��U�Q�&����L��G�z-8mrl.��H��);r�S(���i��a������f9N�4�8��'�u���B�9��`�8�X�oi�0�}�C�1B��,�.trR�q4�)��/l��ޤ�|���(���S����^AZ�	�����ed
�!������l7�[��G�:ˋ�5���,��Į��$�;�r+�f�����_�� ��ס]��o���<@��Z�����"�]�1�i	d��R@ׂ���v��������JO���W5�!��j2���}�X2����W�7c�Ρej=RVݞ`Qwo9�\��q�"�6e��ưTY%�l�~|�o����r��n)�h(�k�MJ�薺�f���T%<������nWu��m��98���"�Vz=%�ڕ�4��:O��^t�6n&#݆�ҵ(��'P~+X��㢖j��Ҥ��a�6�*���ʇ��2&wRQE�#�ڧ��J>��7��T8(y���iL�z~�B;�_˿��{�w�*��o-���F���a	�s^�ߔ�v�F�"h��[���\t�4?�3�C(����IY�;y�a~W�@!ƈ% =@����^��/�(~\
�oT2	��?�	f�K{bց��@.R����C��oL��n]�cZ����φI���.�HX_yz��w]�c7K���9��Tm�޸d����&�U�rv,�-�v���X-����]n�Nף�}�3���0�~a�l�UڛdJ���>f;d�������"���R_ĩI�//Bc�_ְmoK�x(P#7c�R��xj��{c�lO��-�N�A*���6$�8�W}��"�54����퓊���,���:X�4��؋M�����W
�4�R�N�B_Ѯ����$����6�p�{a�N���B05V;��I#��%01^���`�����1O?lci�1��K�O��~�l	 8k�d��(��Es�?7����:��K4�1�G
�A�~G�*%�d��@.�'��b��[���L{�_������uS_yzP�ʢXr�����N���nY�YD�І}&)�Q��#-*,�{�]�8M D�����n��v����e�4���+��N�j���uÁʝ=`��&W�Rp|�	)<7�2Ls!��A���
�6J�qK��������^^�#\�I���m*?7{�m�,�S�w�	�
�7��GvSy
r/����.��v��d�Ś�qS�O�{	s�>����H�{���mGZG6~����n��X	rJ�u�?�V�U&��m�ҍ�z;sؐ��zFN�1G��gv곔`>��"؉�}5�4"~MeN:'菷�a;1��G�]�(d�yzW:���������+�A���$��Gi��y��Jr%���駻oe�9���4�>I�b�6��jN_>_j��w���h���\c}����V�.'_E1���Zyb�TD��j��j���C`�ͨ(���2�W�!�%��f}CUC���5Lj�m�qʷ��VU�K�����6Ȣ�<��	1��&�U��j�p��D�yS�Wh:�����^?��J�/���¶�h�}2�}�UC$���=	��u��q�0a�!/�R
�E�����C�"��!�1�y���>�)>�d�X�S�	H�~��H}g�z{[K���F
����M���.2"L�jTJ�TSN7��E#��<�(Zu����s��LFdn�	�� 9B<i���
����
�3��ȏ�LǗ�G�B?5�j�˷�A-qXS���unV�;*���*�"`�ґŴN�L���A��܊�B?�SԪr�ۣ�R��� �j����L���wEGq���<հQ|��q[f�W0hx�y3�b?�D�ֆj DtqK,G&9)�N��ZZ-������MA'i�h�z
<�2R��EA�k\s�W�	��v��1��u�B���Jw�On�9-T�>�_�0,��� ���2�)�r{��z�"Z#Hd�}K�2���x!N84�zړfBK�g�j
��wI��,��@q���c�A`J+����~H8�k�<N���[�B+rZ縺K���E$n4����M��ld�܏���1U79 P�D��<=m�1�>Z�w�d~�0f�u���#�r���\Y�瓫D����=�P8Rz��n���G�^,���t���/��Ҟ�F�(����f7�@q���F'�=�꣓<�V �;o��O�	�I�}u�����C��2,���d��c�Q����;��}O2����s����]q�$К�{P���$لz��,*~E-ù4�s���]/�x;!e0�M��*t�
b~QD��]�$6���j�p=W�����t�!�f8q���`j�N+�|��0�}�}6"f���5��pz �i�l=����R�ك;C���2��j��J�uV#�|Ky�3�ν����+�$>�$���Ͱ�h����SQ���~>�;��D���N
F��qj;��@�LQ�0A;�C���؍���,�N6���+(���lǈ8��b�ڨ�P|�`�c�R�o2����A��[k�гԼo��p�� i�!�-�]�4�����LM�44f�XYjX�����a�}f������`�C��~��|����m��DE*c��PF\xбk�����-���<k_����kʺݬ���To'=,c  ���-��n,��NK��x,]{H���>��5��dm�C|��ߤ#�ƣ����#�`Uj��W�K
�%�f����^Ɔ���=%�+�r�������ыx;�[a!��}P����f�b��r�9X��(��<��}�A�y�M�4\���^w�i���z���l~����ev�б(�4\P��x@I���^\� �q︻8�d�V9�{d���{�L�ə��3���)5P2��iz��N�:[��	u;m���P
E6��M��	�܃=�q@�>o����e�����GTD�BrL5]e)�8<G��@	!����=�(�ގ�Ʊ��-?��%�a[�k�Ϥ���t�+���=:fr���7�<Xh�YH��w6\4��)��n��hx�w��^v�F�.��A��oګo����|�p�V8���3���j�q�؁�Y�J6�s���e�^��	FR�o)�^�*���f"����M��M���{7�[�V�T#VBd�2���[��߽����K��� ��	�7�-rJ��E���8���z;[�s3{��]�EB��u��'�pbL"����;+�9��ҦP�i�A,��?����8�t�p��˜�j�9@��ާ[T�Ao��3�=�N�T�<��'��8Im�(R���w��ސ��q�/�
K�zVÖ��2=$\�%Xhyo��Үf9,*�EBIgHl��b1�mk$la$v�
n�bD$`Z��z.�;cX��@��|�j�L�j۸��ndL;g��ma�i����7�4Sj�L_�@�v��}((�<���\���՛�Bf∌ǟEl�"�u!�I$q�n.�l5�j���r�����J;��o������}�c��s9q���ZS��zT6l��4�^�/�ƌ�� ��l����*�P�šX�S��
�4�I)�8n�W�ƺ<����ŎH��Y˓QĞ-[^�}o$���7�}TB��񫄶V#&Ѐ�!;u69��^Ө����bW5R�G.dw/�*���Ƣ�`X�}�BTڟA}���xO{��;���z��j��t��p���[bZ��&�ў�{��s1�InW�7G`�O?0����F�V��/Q�8E [�Dxh K��p_?*xYƫ*�x�k�\�1c��;�q��1��$m�c����*��X���P���Z�8��i!b�-Y.�e���I�A:����d���i#Y�E��~g���GQ���& �p�`��h��������W r�v�P�*>�#���}ҙ��@[���v�C�6܇M~�7��/ס�Snhs*���a �������N�%4��v��k���h>���7�mY�s�^��9x��$@j�&ǽ�`��֤��MMP����֕�n��a]9hT�hG��o;�e�)��U)^'f�ibb>�mu�����xa�X��	f�d��F��91wh�BǱ2����=Ȑ��Q��4"H�����_(7d���<�X^ݬ��M�Rv�/~����"T�ȍ��kMd�}C�mFk#�SB����@���%B��J��r
��Q������N�9�x���3�"�h�<7ÝY�)?	ԇɼ����o�`,�J$V�/�d,�:-��}	fL�)�h0��2u�q�	t/,q@x���~K#��N���{F��ʑ���(�:6�y��j����k���abt������E��~��7 ��U�t�Y���Z�M6*�5�>�u@^|��[�a�Vڊi`�G/�	���,��+3�⵺�u���6�Pp��>�ݣX���!����R�����P�W��&��A&+Hf\�y�e@c�D=V_�3������~�+�`g{��h�7|sI�*,e���-�<�^�\pj\2��<�y���f�[49����6��0�
�7!����>���Ƚ�͇��c��k�A%kkއ�c���+�8�����nI\"�Zًn8ct�����.�t`���d��ɨ�A�!�ɮ�5�1T�v i�g_v6d����9̂p����L���.��8�8�4�k��R�kD: ��C�0v=����+cQ�C��� sz`p{�J(����o�0��L���<���S�2\��V����J
Y��q���(Ǧ���ά�U���R:����a�I�4-A��tFt����Z�ge�@O��)��F���}���6�<���7~yÑB��ل��;�ت�>��զ���˚p�=yA�/w�z��dr鎝|\5	=g(ܺ⬎�r�B�����>$~.�`j�v�A�ʠ"z����B_o�����������8Cw��l���Ay1"�}2�mR��+�	���#�.��Q)��Rn�˄���5���"��Z��P��2����St��2']�J{2J��v~EU��y�0\����Mcj!���}�_3䯡+���m6XOOT�]�	Z����]v��m�K����@�| �ꈸ�<��ce��"��F��X�Z$��;zE1ո��d����������.�'䍇�l"�y������,�,��@1}M�!ޝGh>��KA7�qM���o��<~}6���X��3>Y4-�~��KfSƫ&��C��=Tzn���nԄ��#������ ���@��c�	�*;e_�˼�p�T3v�B!GJe!;�sIv��ũ�Ό�P88����!���[������� �H����o��9�w2:�6�-��[�{��1��b�@��/�݁��4~�;���*�������e	�x����O?��Z���r�"3/���:��9?;T�֌��z���#�\�S�_�Y�q�x�q��nǑ"~R��
;�w��6@��dT7���y%�)�Q9+�l�������J��u�!�9Ku�bN&��
��IS�����4�,�pJ�`�>�B��P��A�V�)��Ͼ�X�L>u�`�l;A�Ji �H_�Wh��O{���zDU��A7j^�Z��Қ`�GxQʚ�����+��d���uT�X��kO���}+76j��e!R����6�"�PB���pkD-V�0tn�~��;EJ
�9������N�x��e������V����
�^�j�y���c��J�nR�2Qk�T�
(�U{l D].\���S 2o~�nl�[P��R���@�/��hYvY��7B&�w�����@N�)�s�8�� �)����[$�M-9QȦO���̡tB�-���"��#���Ibab�焔�CI�5��qx%Հ�҅���ض,]�@n����N�d?0[�b�E��ҨS�;G �Hċi�VV���a��^ }��k\�~ bsլ�W�顒�]Q�H6�]�'�m�؆���O�19GG_h��o�a��E+S��m�2�b���:��;c�<O	�5�S=]���(B=�
~t�N?�?,� Ia�8�2��]	��$�`,g�m*���\�((� 7|���kUq�Vv���.	�c�0���j�e3xt_"�n�vC�[&��d�����`o#���V��7-WL�@뤑7�rΠԳ���\f��B�2�
����	5��s�`n�{n��wsd'U�(�T�vo�Wy̫R���̤f#��]wDI��f���:yV"04D�2;e)Q�3�� YA���Bm�5��Q6�,i��ok�W�_lp-Ve9�b�Q�qD�y	�wcDM/�4w�\TVSZ��-(z�5�XG�Ė���<��{�#{�&�<n�E�� �Z��/No��܊&i�
20�������	;Ŵ�Ҭ14��GT��z0�G/�}*�숈�|�d�
\�)��G�@&l�g�o\���ܶW2�ܚ~�Dz��OA����'纚�	�Bq���b*2�TS�z�6eW�6� %dɕnP<����K'6�l-��Q�D��{�c�Q@�Rp��>���Ӛ��lk�9�4�Y O]D@.ѥfݍ��u뒤��B҄�
��w��ʒ�D�
9J��~Z*$}P�[�ՈM+$Yt�$�]2���ݡ����y#�H]d����M�[W�9���L\��u%�[p�������9���A�Xe|CI����@�8�w�|����<"mse�R赗vjX���Vb��7�?���d�dx˵ Z �����{��+���]����*���Ż���f�LZ����H��AF����A����{:��3��
�;� �9�zh�������m�Fl��1`x'>ҼV��,�����i�V��~=P4�;l7� w���*A�k��O��u����{�OG	��:�����(9OL'������쬊�e�_�mwe�6��,�L� 6�s��s��fh�Ӱ��=l�m�����?(�B�M)�-�����?�Jx��3M%f�<�+�8��R�kAɿI�h�B�4ଆDrB�|�_����?�W^����X;➱�{�ԙW�Blm�7EP�8:B�g�b��T���+�f��S��sb��ȗ�ia}�:�$��G��eOZ���)��.k�~z8����}w��rC���M���q���պH�B�yefX�d]�B��"E[i>�V��S�f�KZ*��O�	�Kx(gP��졓�L��V�V�߼��q����TfkT����y�p��K-_ �H��=��
�2#�|ur�Ϧ��p���0Aؑ����I�g@�
c�k#�3�Ͷ����0�W���mo��e ��⼉�B�LO2�Xv�{t�Y�Ŏ"�4���_`*��i���s��6�M�.û��vf�tdg� >g���d�KTq�t�Ң��@�B�e3oZ�:i.��-����`�So6��ا0i]@���]�l�!*��o��k]�*���h�D�	R7����4y
���-��]�U���^A������\���a	�bk��,�V�r�-���X[OD��d�/�k-W^��>3��E*���b����G� ���w]p"(c���(�ϰ�-@F6��Pq�����ż�qH�[D c`��|v-8+��-�KZ2�Qi�����9z��)g�9���8��$�u�BU�D߸��3�O�X��ho\�a�W�'�<$ru�Vgv�%�Yθ;=M��cd�5�H��J���)��������Ʋ6��M��ԉM"���^���xl�^���+��7g�pt�M3�e4����7�C���ԋ�d�́�
Y�9g��t���T��% ��u��qA��7�a�ˬ�<�5\��� �&�����EQ��X�cS�����:Pj��ڔ"�2����_`-���ݺ���p�'t�������8MT������g���L]HȂ ?�����!d~Jm���lm�9`/@�!\&ޛױ1޸���.��=���ZJ�0":����=��V�˱�����f%.�	�JK�����2�%�&��Vs�$��_��{�E��U��g8�׋��Z�e��g�^8N�d%�'��f�ȩ8�O/y��!��e�=�8�Q:-9�6t�q�!�(5���w����M�7�?<8�7�υ���>-gH�i<)l�]8���]�����ʲ��6R��iq1��D DT�ʾ��r�y�4�9I�����NFb�B��\�@��6�Ez�"4��7V~Y/=ˆ�	Qvb6 j���-�j˦M��;�X�<�-E�:y�r��e?#6](%��B�ڇ=&��w�}�fй"H��H��c
X�S-He�9%��;���/���MG�� �YC��}���δ���ˮ`�"��������wMǘ�'6�� ��/��� �	*�S��<�=`KPHym���rX�$�_"aTCb:RZPԳ�I�;��k��3E�F�s�K6�I��o�F0q{1Q֔����=a�v�:�����x��|
��ŰN���	C���,�֡�z����@nJ��7US��e�8$\Q5��\d�;�Q�5��c�>��ھa���(�7���O����o1{�G��ԽnZ����G#��I�BCD��v�j���}e���Dzp\q�h2�38�:��'�G��Һ�s���}2��~��o�Oh*�V<��a0��/����N��} �3c8��������P.�ɺ�3��?��&�n�����=����/�<jI�o��tw�ŧh�M�����rB0��.HP���R/����y�j�uס�$��#��N���mֺ������
�c��Z#��� ��c6i�r?A�: �F��]6z&ȍ�M�l��P��;�(�C<��G��dX���4��O�PWUޕ1�k��t0�O��濟A�_Ǯ�����*���o�I��G-;�C7Hm�^�]������[}R�v��e���k`�^:�ɨfs�+јCs�Gj`��;�C~åbŞ�3y�V��.�Ɍ�X���h�'���e�߆�c�u�[��P��ց�ȀH��D���趾@Y��0�Ք��\렮,׈j��(pv�|�(#X����+�JD�7)49�Iߝj>�_.��A��ʼT=�m^ ln�k�l��!����t���`���[��{&�b<�_���ĩE>�TZ�)3k����Ǧj�	`R���4M�7�RܹT���O�dx�U ��^h��ɖU�m����T+�y���ǜ֐VzF䤭J��cg��E�����76�1�,N��9���1yPLF��J= �>�;4F���6�X��S�@���Q�~A�SÞ��`�:!c�k�i�J� �!�D���o���L��s�}�@����!��0�V>���:�����n��N\l�D5�۽�en`c�ou�53$�e6�_"���d�~�ϣ��`W�U�5up~�1D��I������7�YP�ɷF��3B{��?6+�~�σ"�0FQ,�c�.�!�آ�U�˙}v�o���ڍ1Ms҄�R�Dv�@7�w� ��hCER��y������w�}���(Џ���Y٘��hǝ)�kw���3��]D}��o#�� � �fD���/�ֹ�l�����&H����G�v{���`�y�U����������!����ւe� ��5�+8�5&C���0�~%SG��ZiP��	�^xBR�.��4�7��v��${�����C�jJ#���)N�K�_-��lҔTɬ��4���=0���`)EmyQ7��R����B[��v��3�(τ2�X��A�[��M�������
����+�1q�//��W�(���H"��k��3v�E�!T�4'&���M;�]뇍5�0~W ��.���{��Ğ��/������&d�{��f�·!b���3�,_xc_H9x����uܫ����կ)_Ý����lm��PݸM<�=cED�:^q¼���	pE����o�ׅ���L�3��$���(���Ђ�eLc�E
m'B��;G .��������4Aś��hE�6�,Mᮕ�QAtA�N��9g��3|���@%ǺP�~��9���O��<���b5\I�kZ���~
h���}�f&��e��)Xc������;7�>�0���s��
@8="(r�~���'3[Ӊ���ZB?Fvg_�+Y^@2��U<�K�к���G�X	�����@&�ʋ�[RV�����ڜ���%����HK#��Y1vm��H�s�?��Z��������2CL��A�J>w���v�8	H�W5����~�!VR ��	�1��8��᙮�)d�V��~=<GNE��Sr�3�C��"e��J�%+F��$�������u�NB�O�ԅq�,7�b�p�&�r�����F�I1}���S�2���)�k"��l�}[�nR9�x�"��21�>���,6�v��"�x�⮑��?3��&lB�	�E���?yMiA�"�]�<�b#�$���#A�?���CX�F�hT�&1>(��#c[����DH�G��v�4vew}�ˆ��֨'��7?gs���v˞����^}Z���-%Q�XSRK��P����Q��(��ɕ�qi��>|�.'d�N���q{UMan�����.Fnd��� 8-���y�vk!m����"@{N#�M;�BY�i2�:���[l����y�g@\e���.FR�I#r���T��1&��5�N�7��j_h*��g��{����r�e��8_!�6G��2�D�(�@������]����Sm���6�����-��D^����"��PٺW��[�U�*r����D�Y��z�o%�1!���^��orJ�����Q2�[�
�Éu�W�KD7q�vl������?���L:�h�RЕ#�����:�k��P��h�*j�J��<�u�գ8���E@'K(����]�7���[K��Z�J��d�-e���Ra/+���%{�̟Bxf̢��u�k0�A�)�������v�\2��u!��8=X<�X�B|;�9�.�Pڜs�B������L͢��s<��:�[��&R�O^Vͫ!����Ր�AbA��@
���憻!�#��P�7[4��G�')s!5;�F66��z��W7T����B��HQ��
~��#���y�.�����Н�v�za%�U^����#]�͇b�7�W��ɸ6��|%�7���N	Ƌ�cڇ� ���m3D5��mk��~ �S�6�S�W�����y�G+h��ֲ��;����[�S<ur�xy4�6-�_��ܿ)�ʘ��$3m<��Ag�@(4v {���/
�~ra$%�Wt�����s՛�dH[��G��8S���z}:&!�����S�T������A���;X�j��-���0���#jwva�.`����b��I��:�ns�6����7�oR��g�;�st�/K��77�q��+҉q�Ig�2|w"�
����g��~sHHZ�Y�)�/��5Y�t���Er8�?�vo��i�զd�Wu @6��[�5!��J�^5٠=e��?z`��a~�v<�g�k�������R�or�}�U��8�-��\�|JA��⌮R��=���`��;���9Я�@����0�g���<��`�<}�S(����n|�VĚqcm�c��y<G�鮉�n���^\�Fe
��
x��oy�tcU�|/�}�}8##h�[ڱyG(qgj�`�����Fl4�sױ��_������`�Ͷ�,��<�uD�C��������xtY�Iب�ٓ�he�a#�ع�m4��M�,�,;�pX�6|a4�F�<���p�%XW&�b �����)�����<d�y����$�qĢ���c���3%�b(5�>m�Id]��&��s}~�����w��i�D�j�#p��9��v�T�M������~�MN�B����Qzy�E�����z[��C�E�8�[iӁ	�RՒF!Mx���yB�_��>y��u�4AH���si���M_^D�U��!̍��4��8aG!�h�xOq��O�۬�w�9�CI$4������h�Pi_m�dC��J�7�|��.�:��ε�͎��Ki;��Q�${���З���D�&���ѷZ`Q��і���Qe���358�yC����_��m`C��QyT�J'�$?K�19�Bq��Pʏv�����^&�P !�5���!}����I�~ఴc���?m�:���:�W��ߕKEk��#�KO���3?q� ���n�B�ÙFg;���5�%y�]TR�k	�~�I�le� >S�Y6�F��]C��5�$�Z^LSq��\�A���̋̏r�jS��~UK��]
o�,p�v>���DMR HY�����[��]��_�ЂϚ�N�X�L��d띲�誌r�x~����kʢ�Ó������8��J�%y^(xC�P��4��A��Tm��t������3c!]{��e{U~�M�t���f v��2EU,�+u[�Y��$>l�\~Ǒ�G*Er���k����+湆��ww���?��?�= ҅6U�Q��qǱ���H���p�Tox�q�t�a�N!�j��� �r���i<���w��F<L�{}�I�%��B�pA�d��@�;ϒ�2[.=d��9'�<�����|�tTA������*��,�{��8g�6�!kcI��ȣ�s��}IA�Si%?"��oTҢ{��hDKf������.3��x�hn|I}��t�[�p�5��<�~Gkm�!>3BmI�՟�#���g���H�BZ��E��~���
J����a>��w�+HyKB/����Ѐ�y���K�)�ۯį �՞=D{>��]�vz�O�*�F�4��}t,�	���x�{ �e�-4�~A�nR ���hI����Q�6:&�i�[��c��ҍ��h��>�j��#PQ�@m�,�����{��*����2)4�Tᶤ��:7��A6� �]2�h@�Q4o�oͯ�VP��¢
]�@�G/�y2�n��g�?����j���=�Ae�6����T-\CYwT���-ϗ&fЀ������m�*d4���ː�h^��E6d����k`�K�|݋�R,i1��8$>�N:,���VNCL�1�a�ߩ�{�>��0�s(�6����tg��V7?���*U_O��<�l�?����v� fq��"�֞	��)��҆���	ϕ�+ �A�_���|�.Sw�:�^���2/���%�̘��:�ն�o���7Q����7m��z����-42L�['�!�������`ƭ>�A5lP�LT.y���5���4�������ܢ{�ZC��l�}��� ���k�˱�=�+�F�YՈ�:0	E��.ϛ�/�g�PN�?�d�㉸�/Ч �$�7*`�4�;�����	+���iC��!/$[蚯K�]"f-��6'Q�%iH�as�F>u|N���ڪ��N5J�)�m ��U�Y2��//h,��H{�i�M��lg�m-W�;�`�'*�{D5-�t�*@ޡ����4�l���������.�V� �%D��t���G�q��;�x+p�F7^���z�)�Si���oS�j�9��f ������ i�:�ʫ .��ɓ�ƻvd�o���~NS��	Zmw�ܢ�lю�A�	u�s��Ū�T�n���պ����u�Ż*�[�����"���XOg4 �y�gi�J�J�q�z�
va���G�f�j����cւp�2�K�j3K_�0ꊌ=�,?W�ջ��B)ý?�〩
M1�&%�)�	�� �_S%.���k�^��]��#����y~���Z����FZh�۵������������������~f���UVD���4�L,Ka@[Hc)�o}A�`w+{F˚����6��bFX�E=����qc`�hx���*�FP���W&������S���o����ٖ��X �ȷ�5�T��)�$���V�����d�R�7}I�__{ε�� Q �C���|Y�X��Ğ�si�1����������b���~�%:�̡�3u��oQr�Ȥ�/3��L�� 6��XA!��Ko�1s�w���6@�L���<R?'��	!���tc��Lj�h��d��a���PpV�F��٫�� �אJ�'f�C<���jٍ]��E;fߝok��p���#m��D����=�ɼi}l^������qsWù��F%��ʐX���T��`Sˤh/�r���v��7$pի�!��ӏ6��M O6�	��e�A�N,x1MZ��´�a�Ƒ<�#�E7���wV�j���q���/-X������gA���� y����� ۲#�?o(���y���/�tmd��Z�sfZP^�}�#;��1St��Bn�J�#"�ڸ=4�R(���$D��'��Xy�BIQ�2�EH����,̣I��ij�393�	��Io����a��O���Ͱ�j�M	0r:s�/DIlX� E�8��3��g�Fk�M��i��v��rئ�������w�H�а�M�~f;�{�6 ���l�xO|K{�'#����@T
�߫����p^D7�q�O�j�������_��y`��fm�����w6z�C�#��l�1���!������<g�VR����s��4�P&�"��xo^>��\���S�>�vr�)��ţcC�ߠLN"M����H1d����4 �А�[[
X��-��:��5j[5��#05E��P�1>�P�Ş�ƣ�nc�)+a})5�n�WP����L�����i�o�f���������>�5O��ؙ/��ݐr�,�R�ҶhtpZ��}��q�ea�ߗb�F[,l��3���u��sx`(F�z���'f����J�����Dgj!� ����܁�j��j�	űn!���z7���23Y��=��}IZM䩴�O s�ܼ6O�������s����M�}�A�-o;D:���4l�{8T_�`�HQ���Z����A�G��J�&�̲�N����������)�	��w���o��;�m6�����g�����g"r>��,��ŝ�m����҈�P�%����t�/��$�f�{ݳk��)A%��p$�����b��^LUCae�yk�1��X:�#syg�+���s�a�9�H
�&���~"��'����_�}�S�*g[KJ�ب�ƙ���k��̽{�d�-������;��2o����~�����!�܍�nP���H���㹈�=�	=�9�4Z'E�s�+(y�R�M�� 7�U2�U9O�ֶ������^��<�5K���-iq�
Rzc��IPx��p����� �(O�[u}�x��I����S<������9,�Ƴ�"K	�Η�����������VV�����(݀���i`��F���蟵f��.��q�?�&FnlE7�|�ũ�c����ɹ-%�1�	�u��x��T����G��Wț�Q{i�m{���%8��mDI~R�O9���Pv꩙]�V�5����vD��u^��!%�zK���\�)��*��U��ʖQ�K����$�5�Ϡ�|Cyy�8<�
�x��I�V��ܴ�Q��L��h��+�ę!�"_X���<��5���|�O���������a��1`�u䂈h
ٔ�f&p�͆�_�|O�̕]�R.i[%��.�� I
H�˹D���m>DjPq
�J{*'�%��L]�\K���9�r5�X�HYQU�y	$��[����Qlð�R��i�/�s~S�D���/�d�����,�+`�ad�Kc/�W�ʔ�F��T�f�%��{ �������ژ�c*v�V�O�y�=���?�R�8V��V����6;aj�7�]d���p���Zc!��i82:��O�����[�RC)��O�;�<���&ݡ�XɃ��F�QʊsaR`^�y���;Ɉ���D�Ӷ2��6�ʧ�E�!��{ҩ�6��� a��Y�Y ��P�So		�;��,�*	z����%v�
/:����������Y.��0��M�{������l�{Hia��:��l��Pf���(Xk�F����x�a���� ܲИ�ts��]�'�E�������C���i/!�L��{��
�N�&{U�r9?.퍏x@�IP;�!��_��+1��t9�J92����
k,���+#x7���ٔ�Ze��D��-����PL�.��KR���K����D�L�O���K���=�6�K���.����5���@�1�4'��	xo�%`�i���m��(�~>cu�B�f3[G:X�s(�Ѐ>���{�3�\����,�)�}���5��� �p*2P��z^ ��p�����V\+ {Ь�]�e���@�Lg��	A�dU�W�W��զ(�c�������u�B"��+�S��uKş�<�����iD0��̮��-^	,$��R@M�΁K��a��3^��@�����Fަ��Jٛ�A��$�+�$P;v�E�!��t�^��0t;g4��M�2����/���S�Ȑ*,�Q�0����������	a)+�;$)l��I�.���	Ht+)s�����1�z�	[1@+�%�����������:)W���3��ҙ�����c�<~�rH�N�X��6r��Ԃ�۬RH�A�(2]�K#>f��+B>��I��֯.����F�·�)��|�`���!K�#0�Hq�a��'�����+�����
��Ȇ!T��A;G�:���ݛn��a�K�	w*�i?O��2���Y39A!g�H�j��閁�΄*�i��'	���@# ���hVc^��)�B@_�T��W�,��a��׃�p.rT�'�!���o^�h�8����8��QpH3w��Jv^y�ᛛ�{����ps[�W�2��n�J�ߞy�((�w��hmi�9��F���?2R9�\z�R]�}��XYcG�p:�(��UI���]�qYrlA����k�+xq���g5.�T��^��Ti���%`Q�1��阵�F�ЪCSyX@��ɽ���}!C�w�������ݏq�.��^#�><�+qw'c���陰"�q�)j��m'2�*��ު�v������6\U�*&�Zm�-T������}L��`��&�[�V/5�]-�w��*���X��WZz(�]�`^K�Iܩ=���J�T^���y@�je�t�!�-2o! ��\�tt���]��	)dTٚr���oƊ�ׂ�m'e"����R%�����	[d����URf��
�o<�G��NZ�4B��0N��;��+�w� ��9�����KX���%@��(�X����5������~�< �J�]�DD�ix���\|����݉P{-����$ڷ�"�ꘒ��c!�q��w��*�c��}P<uZX�����0�(1�v������4%ۘrx��M���UY"���ѢJ��k��ozه�	s�ڤ��X+��%f�4 Ғ��TTE�k��J�L7Q����|����8���(KEU'<�
�OS���:�2J�'-lF������Q3���iih��#(��&(���7_T���p���=��j�H&�ݯ��MnU�J^�2��c���B��=��,��[�N�d�Ec����uK�l�5��!���C��*k<��6�韃���u&��mn�����a�]am�^����Zy���U�Ue�lt��h�сs���������ta.bcP9d�h���|���5��
p�7l�\�V�жo~�ΰ]�\��%R��t���} ״�L�Ҙ�j���""�,��K��Ɓ�I<r�M{���*���i^`7Zu�v�s�+O�+���h�D��ҽ[eW<��Vi��=8�������T����-J�k�Y��z��g}\c6__�,-T�����=Xr��"��2�e��A��7�x^��ƍ%��k�<0ۺX�^y�.b��g�B �:t��~z�W�x�����F�x1�D�.���m��� �%9?�Z��ߝ�,������b��R<n�ү�Y��\��n�1�r�O�����qMĉ骔�5.8g�//�/��Q�w5qY����NKH�f�X�
�;`��Qr��uV��"�&�z3���U��X���y�;���6�@�E��V^����9�~m�����F;0w����~{"���q,k;c�Q���ҘFq���ռ��,*�Z|����C4�JŽM��-:�f�(�5w�iP�X�����U֥v���<3,�op>x0���v/��j��o����B	$��퀿�22.$
p��F�\�XD1�$H��T�1qZ�%�B���yh��V�������Ռ�
{,+�|�U��`l����;�W�m̆�����A,Lj�vfpe3Mh0��Ý1.��1B�%�19#��uz���8�W���`�S�K�lc�M�5�0;'_������i�-dr-F�$:K+h�4a�C5y@�}7H�TF�Hr�Y��늮,���IC��ɺ�rG�(cU۞I��߻�"��~���;ܮ���)�8=��+G�f���|��IJ�kRX�`���r�!�giF�3a#�<�{)[�&�`FA�p6�|���.Q�i�E¾��UvFj)��\����� ˅g+����	F�;pvp�
ll����u���o)�e�@�񤟞U{q2�L.6g� �rȧ��z�x�&��)��8���q�^UH���15)����{�鋀s~aے�0
rz�����׺ 5���l��kz�������L������TmV9j���CejS�H�n� 
�<�� �T)�o��;%���Qa뷦�(���7��:W+�%�'���F�ӷ�c��B|ґߚ���#MaEÛx^��3�0E�,ՁI��y!m�eg����8��:.:������W�1��	q4	@. Zmi�GH��*& ����	 ���V�������^���+Q*Ȭ�2-��3��iju�6f���ƌ8��R��Z�L�"�xw��#�δJ--,\��}un�^<"���;�72������(j���x���M�Iy(81�9�:for/�?�d��f�����٩���NC,��<=~7��xB�v��d�i�1�5��ܲ��HzTV���S�f�F�Z��g ��{ث�g�|�'��~�
�ѧa��G[3�ɚ�u��ua�4�J7�d0&��V��p�6v�(}� ��3r�n�����R�zj%ԝ�sV%wr�B��x��E��գb�\�~�"��ag��l��{JzmXOk�e1�V��PtA�U�ZH�)Ke$�Q�8̣#(���7R�<�����n�����x�0h�	Vt����"$�d�a����$I�T]܆x"�_��2RI��}�(v_�B8���O���͙w�	ٶ�v�'��9ƺjL����A�����~G3�7nw�S-���op�}M�0��Qd�ȶ����%�=������τ���j;�����צ+&�/E�cB����"�<�"	�-�o79�W�V�x)��1��3�\�}�6Y��Bb�rS�ۋ������~����jcpq.���z��r�1�*�HMmӞ��ws�JhM�m�>�|���*q���;/;>]����Ƈ�S���01�\��
cH7M)���8e[��Q�(U�,P�_�m s�x�����X���,�����V|��~��hx0�r��n[��>Ա��7���OI�ݲ�C�"����C8uy�QX�~��l�x=Qe�DHS�Q�x=�0�0[^���ݿY��H���|���j�2�c3�ڲ!�JS(<��~!ݮ�Ĥ�^=�-;�-���A?�g�TO��4wh���}e��r�Ϭ[�e؛��Z��)�-����dT+�xXZ<l@y/�Q�zrI�"�#�o�	nAs���N�)7�o����X�$��WH���G���B���Z�S�Y���y����4�wx���P__���~#E��5�����tr�ֱ� ޏ�M��/��yAjJ�k�%%ޮL�ab������<ʈD(E	��b�'�l�R�����G�N��7A��nt:t�<�kr�T2��37�3���#��{�6m�ŢF��q�����&r>��N�0��L�'0��ۥ=��~�e�L�.�Lu�8Lm����u�䕇:����P� �q��%GDh��f�<���[��N	N�ܲɯ���k��*����`(����P�M����q��c������2�A1�CV5M��.-t-�F�Y�0냊tEL��ЈļQ�2'�CO���F0����ROJ���v�a�P,�����)B�M鉠���{A�Zfj���M=Q���0�^�t�$W��>���KW�� �s�1�ksࣿ���98��Ck��<A�~�� J����Q�rc��	����]�
.��(W4�7eW�6ܥmn�����ǒep���Bz6R����TG�Ac$)Ǳ�	Q��x�}�ٌ�l瀕F�;�㫍a�F�|%�5��S� �Z��^�<&�ų^现����"���%F�9���gq��H�m���@�`����OČ�,ؗ[�<Jk�T�	ҁuDE���_�1w�:�0e-y@�8��#��F�W�#	��o�����[]��7���ޠ,+���]�2�>��f�xY���W�W�u���:h��N�����d5�[�=��b��^���u�b�e,Z�zbK�����h�d1p�~�����=eje=�ך� �cM�����5vM��f�Vn��oa�f�W|É��<��
�Eu�,�w0H\Š�f��t��_#j��<6���{dˁsV����T�P��61�x �Ё8���ޞ��h�o঍��xJ��v����K��Ɓ�أ!��a����lt6&	t6ޜ���ȯ���X� ��U�+o��h��� u�
@�V���6�����^|���O�f(���^���
u�}؍!�h��Uij��kS`s��k�w����~�&���<��EZ���ʉ�/�ڌ�>x7�/I��Ӛ��"��3[�z���2��Ǖy�ѭ�&�ĺ*Ak��� Z"�e��`�T�����?��Nry�]:7���Y�a�z���xGg��S!�*
��QJus��*w��p�������H=4�b�(���\����o8mٚ{�\-,���s��L�ɒW+��~���L�܋d�fͧ�3m�&ڕ`*�:E�?cN��j�����ūJ�ة������n��>Y�R��&h�Ш�A&�� �4�nZ�?�6�ǒ�N��$\�%��R;�#�{	e� �y?c����7�����
�Sp=�V�L�L�;x3
�a5�E:�/BF(���� ����['L�����_�G��/���ՙ�s�p�q/����A�{�jkkE�a�gD�e��6����z���R�QC¦����㍍��`�}B�j��F������M+āj�,���Ȧ���{�-YH'i̠4�@���knU5�X��rP֍��U���)�B��[��~�T>�.HT��]���J붨�j�����0ؗ���#H�p��L' UN�	��^���t�U�����8;�-p����>�᫘w!+�hÖ��jVS<F���Z�v�v_1lуU��,w�}u�?b!X������X�_���&�?����
vZ��e;4Dh��mz9�t��SL��3�Xx$��C�JA���0�Z��pa��