��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG��_ �9FL#�>�5NAd_�9`�Z{{ۈ�{H���q�'N�3�j����/�@�>r�9�3�AV���FNU?U��9:%�<�����4sT4l)@��Hcɑ��i34��P�ȷ�&��i�zI�L�)9���k�	��C��c���m<P�������7&F�]X��1��a�Բ����`���*>���,��#��<���bg���_ڂ��hd��6w=��&'�kM5X�VHo����1�EVxfcG�U��ǅ��g��ױ��"��\ `L� Ȭ�:F=7�A�]��)y���>^A��܋h	��y�I8�H�ıɋ�F�+�h��O��D��@Щ&�a�V�G�V,/:�tF�nd��m_�[+���(�1�ѯ0��嶥��,��c�ߵA�+@�|Y=ѫ@�T���Rb�-n�Ϲ<D߭8'��W�dǣwxb��o�j�x�E�6-�|"�|.�;ID�5�&{�"���A$��j��Ks������F!�e|3B!�,c��@��n���5����8��=��+�q�즟���x���f��'������:�ge묀e��o�h�{��A��@M�2���I'"e�a����_$W��V�K;۫ɚ��x�~���3xW��h~E���md���I��775���+���"�����W����P?��8��iϼ��ޓ)�C�h�lџ�Ԫ�I�@�B1�&N��c��{��᭢]z���w=9>�-��l4("Hʾ ��2`4��6�u�U���^$!�-�L(Jt�����R퀬���ڹ|'�\����JeJQA��6H됦�����^P�hX�v��l%�ڴKO�#RU��vc�����|ܱ�Z�@����Y��|�����$��&b�!;���`5���ɰ(�������MӏU�ؾ'�/���_���c�_Ȣ