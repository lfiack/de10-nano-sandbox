��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG�V������ܴV�������`��m<�#n
y#�r@���
�y2��D�L�;�Z׮I�� Hq� ���6��m�]1Z5�m�-H�8�4d��W
��h�u�]$�*��d��lLqa�/R��B��2C҇�z�bm�S�'r�Z��M_�/���f�l��C`�/ҁ�Q�\�a��uWE 	�k��F�a�P�>�S{׀(�⹣�zR�h���*�DC��[�I���Q<��g5꨾��ىi�;��	�1�1Uз+���]4��kٟf5�G#�2V��)$D�0�.�-����r�}��.�m1<T>gR̳|%�Z�Ń���U���7G��~�V�Q����qׯz~���̫_�щ�?��Q�J�I+[�����i��'X��b��1�8I�y6oc�p��y���#�@ne��Y�R��{|��2|;r����ej�f��K�ν���+k����~����x
�k`T
U���k
eBS%�~y\��^4g��� {/�i�t����-�n�5��7���ZV�}I@Ė��$4���_W �~��������+�%n�  *�^A)։��h�`j=�LC�"���#�r[�%p�����M��T@������*w����W]q����郟�yEԡl�g�숛ϧ��ɑ���o;� ��F���V�0�8�ه}�!B�2��[	�ܖ�kw���3Vk�i�p	��V�ǉ�ulG��3�ԓ���.͢E3- iF�����s��N�.�#?�!�E����_�q�dCw�����dNn��	������[�v�y}�fx4�`�O��W�qf|�T^gP�Z���\� H�U��F�foN�I���0 �{�{��@m���*��e{!�)�h���!ߎ�,(6	2�wUٕ9�H�Pz�|��i]���>3���p(��M�4W�':=����7���$�6����#%j�$�5F�(9����}4|Z��Ĭ�>?tZ��'���ꁔ���N�,5EPӂz���q�l����� "�gԏB��鶷�-.�+$eX
Ņ�6�p!�v�3�y����>ZT�B��do��?ڀ(��(�G$�8�Н�z���;�,?P������q�[J�.��R��gP����i��!/����F�~�rU/�#���#0	��C�z��}�.n�<7[�do�jy#U>�����j|�S�u�La� v��}�x� �L���P�7�7��� ۄZ��
Z�:���RBBK` sXm�멺�U����k��b���)����.b閑���d��&�"?��Տ}2�� 4���ĳ�>�g�k;.aw|���=���|�Y-�'~�TM8r�/���ed<�dT�<u���Ny<M^�V�<�Z ���ޝ�;E=�7��4��2�	�Ѿ�G�_y �� @XJ�g_�@VJ�ږ�Sc�2( #$"d;}rV�G��h��,�@uq�zc�~�����z_��G@z4ԡ��PU�GO������
�Z�����_��BT�j.p_/���vZ֭���C�R���/7L�F��X܊E2���G�jÈn��jL�/T���Ę����Ą���0���:n���5S��2E!�8;_�XsRr�Pv|��z�����>*H��x�e��A&����2�{��jsչ�'dzt]l�$�����PkU�J�a����?�Qb5��m�1���1�P�y1w��K�\����yj��Ŷ�<O1�����c�1��q��C����b�En��7����@�w�$�Z\��Ɠb�W��K����(
\���ʓT4{"��d�e5��1��yM}qv�@R{�g�j_��Yp)�xqUO���¼���B8{
���A�͈����*ѻ��(�'ʝ?���nꕪ��C=$h��ԑ���]X���Bo�>�0V��p�yTX�״0�_`?VE/9�:�_��F���H��F1�����ȥ�H�ӝŞL��z!��=��͑������2�h�|�]��S24閧��g���l��G3p�}�Z�I*{#�v�{3�w,���1���M�a6��R�叓�6o%n,��DO�:�Ǵ%!eoGUj��;
��,.T<]!<WK�����Ye�Y�;V+�V��A��n�s��ƺ�k�oh�����V��f���~���84<i��?d�Y��	��%��d��>i��gi����j2�����o%�����/����][�@uw$��kx����ϕ=Ѿ`�I#x>�(�`��_��%W���/���2�V|���>	��GH� ������?~��3P��;��5�Νu�-&Y<�
��M���5�:D�A�7R�Qy��%o�i�N��|��
�"�����[D��a���2�l�,�x��"��/Q�㖔ٱ��k�r��@1�O �p���7(�*� p��T�k�� ���}��[��X;q>ྊ�qsqz`C-#���]n}�S�x�ju��}�D�wH�����
�Dl��rlr�l� �5!X�:��J���T�5z���2���z�0��qt�{���<f�N�9�)V�*���zrr��vR���
Pm1���d*�#�=n/����^.�s�J��l߭�Դt����Hp+&�1���I���ݝ/�(��m�3%��kd���!(�ݞv�(^W�lG���	��n��WoY���D�Q��4�`-�&'�
.�+I����ѡ�^�{�P�k
؜-�8�^$_.#�2��{���DiQ�����7Lșϕ�b��_���R붙��3&��9���"���Z��'uh~	�?�z6Ġ-�e밊c��	���7�Rj�T�G<�%>��WqG$r�p�`���_n,�Ȍ냧�,��H-i����O���
��<�7W3L�#�^Qޒ|Qf���l�>A�Q]n����C~���Hl�s%�á��ɨ�������v2���l�"�soCU���w�$���4���z�37��ũ��o;O�Ig	0Rֲ?��rC�0��/,*�^ISZ:����%���,�Q��EcF��I��\�r��^H�^P�m\��"�N;�t����\�.=��c.�e8|k.���`���28N�
&4�ث�,���:��M���"a{�)%�W}�I�P87��fȹ��=�	�ଝ�yw53pV��Rc��`�L6�׌�MG=N�^I-�"�o"-Yv�����ф�zkq�^�Δy��RiД��B�܍���Z��(�M-#�H���m!�	!+��+�����ڜ��@�$��	avg�?5��d�Lx=;���Ȱ"�g�� <�q����e�C+ڶ�����Qa���<�t��"��Vv�X�}�͗p�9��2��|(l7��D1rG	�=P��\��M}#����xfF�R�� F�ш:y}��1����Wֻ��>-��p���J�t�G���sr��� ��~�M�j:�3��٪_�V���>s�Ԩ��3�Mo�|��)B��_���?�N����M�02#Hwn�6�M� �P� �W�6�'{i.�0_S°���u�g#��d��6�	u��Mu_��p��z� ��`q�\^cs��_�M=�5����a����X�x�J!�6H���Y��m���$�`�� qL:�A�ֽ����:+j�.�JM�m9�ĢM��1: N4ca��{n^)��\�N%�q7��#�n׎�7�lg�.�?���3��O~1ea�\�4�5�8r���5¯�Ɍk�`pG���o�R�S�:�4��y��zNX>#����,�(A�mW�΄�3�@�2��-g�m;iv8�M~�嵱Y��oF�u��7�@�������|�0N}@��_��(�c�{填�y�����{TF ���N�UJ$��%�M
Wu|��S=�����l�����0]R}y\�|2tW����#\��_������p��r��eJN�'���������,��,w@s�� j�y%j����q-y��c���ve���ps��M͕��Z���~z��6YGR��}�`�
"g�����V #���� ���U��L��C�`�(T��M>���69(O+QI�����F�"��;�B;E��}Q�������楁+혼?"|-��WPT+��3Kaaf\���rvJMS��=ԥ�Ew��c�}�(;��/��,� ����yUՒ�	Zw�C�z���Q��5�0���2�����С�G��
�ƿY����K�P����B�o�Diw<�����S��6Z`+��A���S�wg6c!v�O���k�IL��i8�v�f����q~?dh��ڳ�!��Ih�q`����'=[��i�rMi�sƺ7@9���D@1��;�	#��W���-#6�	�Π�����Z1�K䯄k���:'���@�**]�+7�c�2�1{q��亷MM�R�ύ��̩���;���כQ*���Z)�S�ݽ�XOl~�������d�(�J+ģ��]ͤ�4�h�h��:"�h�k�8>�a�[�%��e���9ո�%�x*c��T�-1H=xSPiZ3��\ўt'�����Ӣ(^;5>QE���;�<�)�Ky�'�&�.*�4�'���0�|�O��Z"쟡�$����Qigw�d®�Ľ�D,��\��\_��X�cyc���:�z���FԠ��l$��(������Y�n����1q���~��r�hN����|B����5�ݍ]|{�.u��-�:��5�گ���v�S�o"iҠ��������߃	�w8����.�2���]X�D�$��#wn֢�ԘFݥC�tH�f�$�U*�Ks-��?�dRA*:~YeG.�k�����5{ee?�aamY,���7mF딗-V�Ϧ�+^��lA@�w¿\�1n�X�ss`��>���CP��U�`&{��΍~�!��&���%C@E(B^�t4���"^�Y޿Z8l��)�C<N��fs.��,�n�q��	�bˑ�m��C���3����+&��!�md9=���Z!�T^{�UNN�,ٚ������8�x�r�%���0p�0~Fp�Y��ؖ������`(���W���E�Z[)�����F�p�����(\�4M��D?��JK�c�r��������s�\�����?�ĔLy����]p�W����ؘO�|��q̱��̺K��PV��6�*}�Sw��