// ============================================================================
// Copyright (c) 2015 by Terasic Technologies Inc.
// ============================================================================
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altera Development
//   Kits made by Terasic.  Other use of this code, including the selling
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL/Verilog or C/C++ source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use
//   or functionality of this code.
//
// ============================================================================
//
//  Terasic Technologies Inc
//  9F., No.176, Sec.2, Gongdao 5th Rd, East Dist, Hsinchu City, 30070. Taiwan
//
//
//                     web: http://www.terasic.com/
//                     email: support@terasic.com
//
// ============================================================================
//Date:  Tue Mar  3 15:11:40 2015
// ============================================================================

//`define ENABLE_HPS

module DE10_Nano_HDMI_TX(

      ///////// ADC /////////
      output             ADC_CONVST,
      output             ADC_SCK,
      output             ADC_SDI,
      input              ADC_SDO,

      ///////// ARDUINO /////////
      inout       [15:0] ARDUINO_IO,
      inout              ARDUINO_RESET_N,

      ///////// FPGA /////////
      input              FPGA_CLK1_50,
      input              FPGA_CLK2_50,
      input              FPGA_CLK3_50,

      ///////// GPIO /////////
      inout       [35:0] GPIO_0,
      inout       [35:0] GPIO_1,

      ///////// HDMI /////////
      inout              HDMI_I2C_SCL,
      inout              HDMI_I2C_SDA,
      inout              HDMI_I2S,
      inout              HDMI_LRCLK,
      inout              HDMI_MCLK,
      inout              HDMI_SCLK,
      output             HDMI_TX_CLK,
      output      [23:0] HDMI_TX_D,
      output             HDMI_TX_DE,
      output             HDMI_TX_HS,
      input              HDMI_TX_INT,
      output             HDMI_TX_VS,

`ifdef ENABLE_HPS
      ///////// HPS /////////
      inout              HPS_CONV_USB_N,
      output      [14:0] HPS_DDR3_ADDR,
      output      [2:0]  HPS_DDR3_BA,
      output             HPS_DDR3_CAS_N,
      output             HPS_DDR3_CKE,
      output             HPS_DDR3_CK_N,
      output             HPS_DDR3_CK_P,
      output             HPS_DDR3_CS_N,
      output      [3:0]  HPS_DDR3_DM,
      inout       [31:0] HPS_DDR3_DQ,
      inout       [3:0]  HPS_DDR3_DQS_N,
      inout       [3:0]  HPS_DDR3_DQS_P,
      output             HPS_DDR3_ODT,
      output             HPS_DDR3_RAS_N,
      output             HPS_DDR3_RESET_N,
      input              HPS_DDR3_RZQ,
      output             HPS_DDR3_WE_N,
      output             HPS_ENET_GTX_CLK,
      inout              HPS_ENET_INT_N,
      output             HPS_ENET_MDC,
      inout              HPS_ENET_MDIO,
      input              HPS_ENET_RX_CLK,
      input       [3:0]  HPS_ENET_RX_DATA,
      input              HPS_ENET_RX_DV,
      output      [3:0]  HPS_ENET_TX_DATA,
      output             HPS_ENET_TX_EN,
      inout              HPS_GSENSOR_INT,
      inout              HPS_I2C0_SCLK,
      inout              HPS_I2C0_SDAT,
      inout              HPS_I2C1_SCLK,
      inout              HPS_I2C1_SDAT,
      inout              HPS_KEY,
      inout              HPS_LED,
      inout              HPS_LTC_GPIO,
      output             HPS_SD_CLK,
      inout              HPS_SD_CMD,
      inout       [3:0]  HPS_SD_DATA,
      output             HPS_SPIM_CLK,
      input              HPS_SPIM_MISO,
      output             HPS_SPIM_MOSI,
      inout              HPS_SPIM_SS,
      input              HPS_UART_RX,
      output             HPS_UART_TX,
      input              HPS_USB_CLKOUT,
      inout       [7:0]  HPS_USB_DATA,
      input              HPS_USB_DIR,
      input              HPS_USB_NXT,
      output             HPS_USB_STP,
`endif /*ENABLE_HPS*/

      ///////// KEY /////////
      input       [1:0]  KEY,

      ///////// LED /////////
      output      [7:0]  LED,

      ///////// SW /////////
      input       [3:0]  SW
);



//=======================================================
//  REG/WIRE declarations
//=======================================================
wire				reset_n;
//wire				pll_1200k;
//reg	[12:0]	counter_1200k;
//reg				en_150;
//wire				vpg_mode_change;
//wire	[3:0]		vpg_mode;
//wire 			   AUD_CTRL_CLK;
//Video Pattern Generator
//wire	[3:0]		vpg_disp_mode;
wire				vpg_pclk;
//wire				vpg_de, vpg_hs, vpg_vs;
//wire	[23:0]	vpg_data;

//=======================================================
//  Structural coding
//=======================================================
//assign LED[3:0] = vpg_mode;
//assign reset_n = 1'b1;
//assign LED[7] = counter_1200k[12];
//system clock
//sys_pll u_sys_pll (
//	.refclk(FPGA_CLK1_50),
//	.rst(!KEY[0]),
//	.outclk_0(pll_1200k),		// 1.2M Hz
//	.outclk_1(AUD_CTRL_CLK),	// 1.536M Hz
//	.locked(reset_n) );
assign reset_n = KEY[0];

////video pattern resolution select
//vpg_mode u_vpg_mode (
//	.reset_n(reset_n),
//	.clk(pll_1200k),
//	.clk_en(en_150),
//	.mode_button(KEY[1]),
//	.vpg_mode_change(vpg_mode_change),
//	.vpg_mode(vpg_mode) );

//assign vpg_mode = 1;
//assign vpg_mode_change = 0;

wire        gen_clk_locked;
assign HDMI_TX_CLK = vpg_pclk;

//pattern generator
//vpg u_vpg (
//	.clk_50(FPGA_CLK2_50),
//	.reset_n(reset_n),
//	.mode(vpg_mode),
//	.mode_change(vpg_mode_change),
//	.vpg_pclk(HDMI_TX_CLK),
//	.vpg_de(HDMI_TX_DE),
//	.vpg_hs(HDMI_TX_HS),
//	.vpg_vs(HDMI_TX_VS),
//	.vpg_r(HDMI_TX_D[23:16]),
//	.vpg_g(HDMI_TX_D[15:8]),
//	.vpg_b(HDMI_TX_D[7:0]) );
	
pll u_pll (
	.refclk(FPGA_CLK2_50),           
	.rst(!reset_n),              
	.outclk_0(vpg_pclk), 
	.locked(gen_clk_locked),     
	);
	
//vga_generator u_vga_generator (                                    
//	.clk(vpg_pclk),                
//	.reset_n(gen_clk_locked),                                                
//	.vga_hs(HDMI_TX_HS),
//	.vga_vs(HDMI_TX_VS),           
//	.vga_de(HDMI_TX_DE),
//	.vga_r(HDMI_TX_D[23:16]),
//	.vga_g(HDMI_TX_D[15:8]),
//	.vga_b(HDMI_TX_D[7:0])
//	);

HDMI_Generator u_HDMI_Generator (                                    
	.clk(vpg_pclk),                
	.reset_n(gen_clk_locked),                                                
	.hdmi_hs(HDMI_TX_HS),
	.hdmi_vs(HDMI_TX_VS),           
	.hdmi_de(HDMI_TX_DE),
	.hdmi_r(HDMI_TX_D[23:16]),
	.hdmi_g(HDMI_TX_D[15:8]),
	.hdmi_b(HDMI_TX_D[7:0])
	);

//HDMI I2C
I2C_HDMI_Config u_I2C_HDMI_Config (
	.iCLK(FPGA_CLK1_50),
	.iRST_N(reset_n),
	.I2C_SCLK(HDMI_I2C_SCL),
	.I2C_SDAT(HDMI_I2C_SDA),
	.HDMI_TX_INT(HDMI_TX_INT)
	 );

//	//Audio
//AUDIO_IF u_AVG(
//	.clk(AUD_CTRL_CLK),
//	.reset_n(SW[0]),
//	.sclk(HDMI_SCLK),
//	.lrclk(HDMI_LRCLK),
//	.i2s(HDMI_I2S)
//);

//always@(posedge pll_1200k or negedge reset_n)
//begin
//	if (!reset_n)
//	begin
//		counter_1200k <= 13'b0;
//		en_150 <= 1'b0;				//frequency divider
//	end
//	else
//	begin
//		counter_1200k <= counter_1200k + 13'b1;
//		en_150 <= &counter_1200k;
//	end
//end


endmodule
