��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_A?N��Y�jo���e�YI��#~B�t��@E����2u�@��G^��8�=�Q�Ps�t�N����ꈱX^�1��Fȑt��X���ސ�t\J���6����9*���$�L[P��#L�pfR������N�Gm�IGlr�FUx��盆(0�ܥ�!٨Im]�>��r�J������<{��	,�Y x{��a���T���9P7	����p��(p>��7YN����aD��Z�<�ѭu�W�B#�X�fn�ٿ��f����x�ڦ9B��B߳&B�24��f�����˹'qF�R��nE'��r=	���Tf0��6,p���g&O>Z���^y0�S.��RF����v�����CG<����G}J����y�'b���Q�;�K����ɘ>��سP�̫�Tہ����`J�� ]u�"��Mҧ��Mx�(�Hw�g��qV��8E!/=Н�-�9�E"M�3�n�o�b���� �P�Lc�! n���v�c�>��n�a}���D���(��G���'D�i����}�U��3��;K������Q�&�3����aLxmEQT義46��W������N`�hl���\ �ew!�L1���a���g�]��)<�cG��Ħaý��)�t2��a��_��t�D.���Q6�����̕&H#F�^�(��:��i*F�Y�n�����?������c�E�	Կ\�cb��z:��W,L8����o~��@�F��r�iAds�U	��̺���<�ʹ�m3V3=TH��n��@W	��#���B-�8C�S��nU�H���|����=�,t7s�c�f�4#U�^ :�)�C�+�2�(��a,��:Q�� ����_2�����c�2�U��zMjhHGd@f"jV��:��� �l�Rb���K�#�ƽ���"�}q�D	� ��=D���K�ߊ��3�j�����Z���:�I/s���e@i 5�0��}���Or�Z*���u待%��ia|?E�9?7���v����ƺ�A=uC�����`� 7�n��	��U$!	<D��:�vG�,..����K�.�2[o+����x�͞][�SNb?6��b��R'���w[7*����oh$���V�{��\o�'�A����em�J�ݰ�t���x��,�ͬp��D8�����Y�AP�ߋңi�e=���[�:��*gJ�
Gz�<MT_D�¬hb�qvf�qvJ���$��K�1�	�c��R�����; �����kN��X��YX"�w/��o�3��~A}�Y*�\TM�va1��e�H6�����������u/��Ѝ�ar�f
sQ�VW|�nSQ�V�5aK���+>���a�Y�����Tf!�����o���gQ8hk'Hk����i��Ij�}ó�ۆl%GN6Y�cyt���(QV=���-}�Z$���P�#t4�qLKY"UO��#��q^܉>��
��!o�K{�]�7�1�pHޱ6U�>lj��r�l��s���#����]D��4<&�h_�����Z-��z�ƪ(A�2��dPč��5�g+5�Td��b�����7 2�[N9�.�=�0�JO�q�vЧn���<l(������Wnj��_��_F�}��6�4\�Z���jKǶY�V�޲z�8v�L�w�;/�Z�ܒ<��g���-^k�+��n���*)X�+�}{E�i�a�8��I�0�&�Μ0W��,����6����)o���u� �7"
�_u�ÅbB��b��x��W]߸���j�����>#�}a_��շ���Ŋ���: -�D��AQ��bYh�/0�E#�6n��MZ�P�����oIL�[��4��"i0
+�k��E�N{�7��w�(�V3�.Ij)a 0Gջ>N�2J��^F��e�:DݤaW�+pc[�9���Fr�0�Z]���Y�z��nƸ!���
-�0ʦ�(��P�t1�4&���a_��������exp"v
@�A�}�qW˓����%�(�Z��F�c[<8"	��쪨��4C�����w�6�:�5���_�D�[5)�ڗ��U��ȃtyo�%�����WR���r2�6K�x1Y\�2�()���c��V��ۆ�&�y��i;�i�n��P�\]� H��n�e����z�q�ҙw���Ah��-�o�����^���#�?֯�W 30g�9�4���/�U�Vz�����s�L/$ y��RL��PR�R&��X�Kz�!���-���
�����K�y�`�2�N�� �*�������K�b����7~FL@ =����.C�m�F�2��x���x��T&:��x>Et�wY��S7]��fqv�y�U��"�>/ū���R��_�Jb@�Ϯ�Q{�GT[�ܫ���$l��kI��y�����+����N�prl�EX͓\����q�p�l=��-o���V�
,w%F����0�c�vg9|�J��(�0]�-=���L?Y|Ce7�餙3���m�m����.�=�G^|��.Ԋn�]u�JR�F)٨h*�K��V�8����VRB��΁�N-`^y�!�.���u����fd\a<�;1���y�W �uI�r��O��ǖ��������/]T�����1�LݞMn*S�+�P�����dD]x���zB�x�- ���3�4h[��T�ذA��2�4fc���@z��%�)��SÈh"��/(�Ys��t`��s�����%d�u&�^�b�D�&��'�h�=g~g�n�Yz+���J�|Ve:���л��+)�J�B���X�jP K�E6T��Qy(E�ٞ��!�1���!Gg��`��We�
~��~Ң�f����N���}M��uǬ��4�#��7U�����@qF�*��<�f|f��ipjf'1����u6�ʶvz3N�ߩW����|N��D ��_�V�_5������ke׉�:;��4MF��rLj �AJ(*�lW@J����ecW���M�/�euU
�����f�s�X!�?���[����qY�Nm��ǀD��:1��8����2�i|����g�̜n��Ԍ7�b�~�r�Q�'~��^��}[�������|��S��cn�YZ4�a����wĩ1=�`%�|�S͹Su}Z2#�8:(\�4�������WV����@��Q�5 r|�&� ���}$N�i�˔���dL386|���{�U�=�-�����mx�Qtt�.WIY`�����R|�H [K`�䫕��\R��]Y��?�@u���ã[l�y� 8���hE�X݀j�=�x��nu�?�,�]�f2�NT���t�>���0���ۉ����/�r����e�}�T9���h�OuV��5,C�2B��wr�q�bR{���X�-Q�OPu���֟@>?<�{;�L:��"�sJ����"hJ� �^So��Ax%�9��j�l,����6���;NǶ�za�8^��s�ʸ�Y�ݾ�&���N���LM Ȍn����e-�M3����;�w,�d�A���4��w��8�K��u�%�9kŚ�g�k�����F����,���㝓�0y�0�q����G��5o|���~Om�&�[�Q���*�Q`����(Ǒ5�Uj{������>~ۡb	t.R�@Aj���~};�1.���)ZL�9n"�f
�/9��N���c��&�BL�����E�s� �W��~X�y�Z�ҳ��tEBO%l��A�ׅ�~/�q7�YL~�{1��rO	I�(i	�ن�i�&���"�=���{��y���y(Y4��3��!ٵ��!�L��]��m9A3�jG�91�gҊ�d����+���Ӣ��]�.�w�ꨫ����_���ʸ'#�vAg��J���Tt����X����W���Y��en�aݝT@k��'����,�M��K6u�@�� rP0 G٧L��J6MRy�Sw��)�d��ohmMG�Nw6 �Y���)u��?,��2M[<rQ�kx��쥾�~Dа�b�C��[�@��z��G�0���ͩ�����)Ih$t��Y;*�?�\!prTF.Bʭf�Nf4��>L7��d���_7�p@�5oJ��!*b�`�Gaח$�f� ��̍��.��*1V	�|�^�?a�����=��G��=���̲_Z���d���8�����5V�(��2��x,��'V�b�<(ʃ�Ţ�&e�;�>��uj��"���6R絢H���n�X�RZ'�	٣S��~��ͦ�侷G�jN���8%�k�P�fx���G�m�	�}��>���+�v�Cf�m��؂ړӋt$��\Zm^�=���l�A"p�o/������5�pO�1M��7�,����v���|�K���1g�e�_��r�լ�oO-D�F�ND�U�O��Ծ��d��|��tE��ۄ;�Ppo���ȯb��0W8S/Ϛ�'y�y��
'�9���"o��Ϳ%φ�"�8�XG)�K��1r�5���S-}���;��2�*�`;�U���^�+�<Ǐ���y7-�P ���1��ɰ��8Ѡ���Ǳ���Wݲ�_����u���ɐ�4j�W��{�6�)��:��JrI�8v{?L~H��|X��~�ЉJ0[�ŷ�zi��F��@r��=뇒'������5��U��X���˖=���X�6Q�L�?ֳa;3���2m*EK��Y�^��&��o��k��LK~1�)��R�O�1B�^�a��t '��:3���nu�";�*�g��?�)�����s���B�)�Cӑ��a�oӮ�n���\2{��"K��V�3!�te�S�����6X����"W,�8�`Ik�M>lg\����m��a�����x��i��g�M4� {�ǹ�;�٧0�}x$��Z��	�G9�m���׏�Hx�C�Е;���)��_�%?|��n�݅��J
��դP��EB���ӴYb���=���|�5�6��	PH���03�h�p6\#�_�^_,�H�%�K��=+�(!�;��q�G�8�o�rm c�[+rE<���'�6&E�z�Ƃ��v���Ivf��Eժ�_j[R^~e�;{�E�7�����������2��V��4�������k-��t9Y�n��b�h>c}������;��3�����c8�r4V��	K��J����4<}��j�d���噒Y?U/�ߡ?O�XuFL��kJ�~������$UcO�S�(+�2�h�gC\������^�d.OaQv���<r�gi2<4X��&����"���.r=R���1
O��O��k��l�~%��Uu�Mk�ޝ>U���q�h	*p�y+��]��;Wݷ�
��������L9�������Vhe/j�vDf�wj�V	��:pC�w����������Fʭ���F���
�jE�ɥ;
��d0��pɡ��v�N�B�f�SS�E��m�8�|�Ai:��^�S؈j�@~OHk���g�P��.�HA(���#�zn�u�P?��;�ɲÊHDyi�zK�3�`e=�� Qt�Ʉy[�������~�-]:b���v�1����T�9l�l�,�?RG����)��},y`2��!��U?��<�Up`�e����:
.t�F��Һz�hWb��ɛ��b��{�_O�4�Im�E}���;�w��E��q���^Ɛ��A"=�.丯.�=X��rs��.���BOc�ӀU���+U^���Enq��;�@I���l@IAu�C���u��{@kM���
��0�*�8nf_֛e#
�%��"����P���`�h,h�C�@�P�]�/����*=|��&b�ȳ�a�R�X���_x�	��*&����ȸl�j��mS>7��� Y���h�i�H��됲r"M�h|�<U�j��|i��rx���"�\V�^���s=��ㆬ�p���#�O:a�5�K��5�Q�Ꮩ9����^�p�ɟ#�� �\��L2�n�=�iG�a�b��jb>��UH��,d����\�����;e)�tVS����E7|mNd�J���⛟���������et��J��YDV�����oًʤ�^%��y��7��te#iFK���X��FO.O����~g�I&Eխe��`�#�|�-����NK%@��i��w��dl����	��a�f�ۊ���� ��$���(��:Y-�ֳSP,K���e���kV�N,({�3��F������������f}�6��f%Y�B�U���7��\\���zS�ێْ�����3�ڎ�ĹM��05�JOt��#��X���#�T�d�P�Q`�G���{�	bd䮌���� ��ك����}S��/FJa�ַ�e�E����mZ�I�v9@N��
���O��_u�y��t�M֖%��[_B� @��v��I��r\��Ȝ{��ʽt���}wS�f�9pS�^ar$������K0��`Ow*�ߤf����r���g�M[WS��g��	����]jE8c��T�v�L	�0�A��^5Bg��53Rv-��d��XM��-�3Έ8�+`�~e�]��-�+��.L�P9���	hZ?�P��pyt��f�)U�rF:�����^�^:gG���q[Aa-,hC�}�����,s6#�=����E�U(�x#y�\P!3��L/�D?�U����V��肒�����H�Ǳ��6K�6P�m��rW�NX�
���3�s�9����� g�hX��ͳ��(�~<D�R�����;g ��xf�ʩ2��m���:��q�Ȋ_~fE�Pg	M=�[���W��J}F���9J5,�ӈ����ز���4jP a�`{���.��X4g]�-*�(�Q
؏�I�Uw���yQ}CVO����=-��,-lH)�#8`����T/u�fI���P�����2�_�;�O��	x�$��$�K�3�sT��9�7��-�_bu*�������\6?�D"8�*�+�|,d�����M2|6#���h����k�'�C�Ϗ���{x�_�4;-�g���K���w����R���lq{H���dz���3X�Č-7��s(	�{��	="������G-�YB�(�K 5����Cപ%���e���[���Џz͵Uý�CJ�9�
�'u���/��g�����U�}�Ҋ�+�o��,�U��MG0�DV[�0CQ��9	v�g�p[d���嫢�CQ��	=�4��iI���`�O��(���D��
.���I�t��mW(�����^�o�����������[]�~��L"Bwq� �@L�ɓ$Kb`�[2��hq6�vlq��OL�u�iYD�T��r �Bo�V�X��7tm"I��v�p���cj
 '�ܳ�T}A��_��k�'���d%�c�K�B�a�!���/؋�F�k�~�R�G����@]E�d�!v�J�,��rf�F������]���4�]h.*��+�n�4P��jq̱�D���,kC���%��i�Ś3�M���xb�rƈ���j���Ab�8���q�A4�Nrxak,wa�zCK�c��<����>��A���>ͳ���;cv�k���.j�{�aqF�ٌ��<Q��>����4���U�����6%�\Yxmֶ`�n	�aq១��!T��+*�fu��s��p8���Q�t�,�uD��|;�U��#l3C}%~�\R3BU��P_Ls�hi�<�零���t��r^�cơ!y'c���|����$�[P��ߞ/$Eڠ���l����3��7�a��qvbQ�i�j'*�O���"^���ԁ�Uv��-�᱓މ���/�1�
A�/���S��У���Eh���(b�.p�I'1����\�ZȺ�s����a@(W%P(��Ȓ�� ��`�AMg� K�����Eb�a#�4,r�ޚ��h�׷��$�O(�]
n%{