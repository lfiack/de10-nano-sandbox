��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�APq�lG!7s�H=s,,R!���#���$aFoU����s�^�&����w����e���c��l;?y���0�Sb)5���kk�h=<*Ã	���_E��sS1綌]b/�Q� ����5�1�é��\"x�U	��L�]�<��l@A�oz'�������\�׿j�2�-��'��	�nI�_^ MKVHG!)���7��Ur�`.xʨ��o����t?���r\��V�`�5c��x���Y檹*N��ΐ8��㰅r���vi�-gc;��k_�t�r"����b����y-9M�ǧ���;r̩��0G�%�|��pj�%ՒB������0��_�_
�I6�&�f0	C4u��W��!@�Ժ��t1��^�lvK2�I���;��<���W��7���V���:�_j(���,�sw�D�|����X�I��ˈ�QF�jgIOz�,%�:ň?���d6�b�s����ᬀC#�G�8@��h�'���A͠[,�z��ˆ�/���d�3�۳\53KC7(kd`�Z٧>n>h6�r��bc!��'9�b|G�s���_���ɏW�SL��� e���(�xm�����'�6�܀4`�)��s��>�/��ܢ�C�a�^/$A5�~N+��K�2���5�ǒJ������=Kjd�RN�g����������4�,H�=�>=\Ψ��C������C�0�9*$�6����5����p� _(��g�i��r�F�g[�T�����ʭ@g{[�t�x�Pƹ�t�sB��9�Fѥ�l��f+�^�Z��Pj����P������F�n;6����-�}��6/{�JL�7��p��o�_�)jx�O��.�7��KZ����n�o1ݼ	}���<�<���S�ﺛ:�I���:�H8��ՏE�4|�1��=�m���Yωɲ��P$�r$�0mެ�7q��ZН�<��ʜ`�p�>Wք����V�&6Ng:�,�j�t ��jsv��ud���a�8� �*մ`���^|��4>�e�*����[�O�I��~��7��.�芚/��\:�k��1@@�6�we2?%B������j(c���/�DS�{�/���h�5@`��"��Dqw���!o���=������G�)��>W>��R�L8�YF8���Tm<�x�_ ���ksaw1�(�#�[�/�
e�SE����LN|ԋ�M���Wc������@2�� ;p=����եx�_F)�R�U8M�Z�"%7���YO�{8�ʱlL�,��X�g���]��cC6��9���{ax�G}5��=O�P�[�x�5�;�x��gW��x�nZ��wzz��YAt�l`~XT�*��ijh�l��=���MCJ��~�@)�sU�"k�A��5����S���﨟ʎG��~�I$~�N�<\�W�l��RDS��C�n�͘)D@�<&�<nEn�e&��0�8Z�i����$d�rP�9
����J	��o2�S���<��+�&�~gj��,$�X��(��ܮZ��7��k�`E����rD4���_*aLpp���h(r�;! �������_)�Ճ����վN����Z��u�1B4rux5l�r#M��wq������~��	��=T#0�J��w�v�g,�$W�bH����;C�ǲ�Y��g��çn{�Uf�G|���z�s$b�A<r0"Y�>̕atb�<��0eܔ3p�M�ݒnQ���Fπo,
X�[����i�͗n�K:c� �}aS�����rl�EW�:�2KDOR�,�Ա��b��pj�V�(��4�[�U�ԯ�Gਨ��ٽX������R; z �+��bi�f�Q�b�ک�o�V�.$Mx�_���x��IQ�G��[��AZ���ɲLդl�*�4Q�/RH��bQ������Qĵ �i&_��J���{mR'D&��V��`[@y�N�Q-8��M���=+OIm�,��3s\�*T��i�Q~6܃8�b�_3���c[čV�l����W Ǡ��v�al�Mۉj9dH=���7���}���]�M�&��ӚU�
މ�2�����6I��3���aR�a��"g?y�HIf�
��M��m���{��'�3j�{������}�W��Q#���GŃi�x��{�C��� 6�I��=񺳘��̸�����C���1�sɂ����~VC�B3��-I���a/L-m�
g�; G}Q��)2��4u�T�-�H�u4�)*�t��9��X$�?>GϞo��Bzs�l����B�C?�x���.Ό���� �¯&�Vzҡ�޵�w�� ����E�P���,�/�@S뇀��vLAA)����e+SV��; :�᱾��ln?��suڵ���}�^�}�wJ��.ਕdj��;.����l<����'�!�-\*�爏�e%�j���h�#5�Ä�������\mcɦ��z�ퟎ���7��C8�� )Za���D�x�O�bU��W�#R�9�LTyK����5p���Zz�w��YLyl7^��	���*�yѾ�%��呶�(��+~3��-T2O`��^ H>(>9o�04�B��b:��Aq��`N�D��^���*i��6U�tCTR�Fj ?��j�����&��k�FG�4G]ۈ�%��N�`�H��k�T����O�`�L�N�pq���ja;vn�c�)�#�����emA@�ZT�6;�3N���9,|��b��/��hVK�QϠd�R���$6+�O���1�Iޝt4օ:c�\���;�߽��ڊ��nv=�]��n[�k��|Vr8{ӵW�L�'�Ϲ�O'`F�ڽ�Ƶm2��9{�L*�e��{�kҫP�I�t � � ��.�K��������f�?��"�r)�8�/��8�ko⯡�^�n����- p+ 5pتŖB�z!"b'��I"L�;U����Y=�����ߩ�'���Q�����.�kΜ��|���[���(�R8O�9�G����cj(r�P�f�"����@[J�ԇ��k5\	���`��q��8�m�J#�er�u���&�a6�S���N /j��x~��)z�xU&R���I���Է��Y�W��	��Ϥi&ُb�n�a1r�3��sv�1��.M���ɋ(���q�,V��=jB�E��|g�ݩ�)�e�K�l�Z���~C=P����b�OŇC$�Id����Y�sGs�k��[Fҵ�=���l 8��äRp�X3��|��*�!	ҏ�� `D${x�꼆��=1\�z�6+k�}�f��a��f���h�(SL���7c���3���T��� L-���.�J ���B��)#���� c�6�d5��-|ᄙ�ё>�G �'����ˀ�O�R�,/4��&T�vl���;���%�؜!�{I�5q�{i����U�� [���e�{g<EM�Z�͹��U�}����<(Q�+�7����h��-��������X��7~T�\���H���j�ۼ���i̒��R���9�<��Ґ��⎒.�,a�"ܖ,��$v(�]6�ͨ'f<y� y8�F@�ܳ���y��b���F�'�GR��Rn����`{��5b��k�E����Rvo_H�=�>ZV�ق�7���Uʱ�\��>�Ŵ�2�v.��]��')n�;����<��}��q���_? �
x'Q5Y0$�(i�k�E�7S�`��T+����'�:�J���f��|�z��k��P�6�p�	7���5�$l����Ą\nv�'h"-{�W��Z�OCL[��s��'�81m�j�'���H��`u\R˙��Թ�Ө��o���p�VVnK���M�xޙ�ͻW���e��iv_�`�v{6Q��~ŕN�;���L �-L])
!���u��%-s������pH��f����(�/#O�%��nm��.��`�p�����\~>���:�����(��>�"a>P�C����5ǁ³11�����,ȘF�TE�R��_�:Q�6	���;r@��I� �
�2�� �)��2z�$�������9$G4*���h���x�&2V���ǚ�9�2OJ4���]y��Ixپ�#�����镁 �����}4��1\�n/��"�훣�x���aV�H:�B�S�>&��Y=��v�˄��!is�@�:c ��z?92%�UH�}��}�x4%���>��p�7���9J�x�l�c'�A��	�j�ǀ�-q��sK06����J)���X���˫�jv�>��4�ra^
�q)�1��B��ڹC�6��F���샅"�o�\jb��W����ׂI�۸�Ju�V+���5���(���"3�>\>�U���q;1��}�Z{y��*�T>d�8N3��C1��2+ӑg�qW�x���"61&~���9�Q+;�Y*S���D�B������5^�c7�����N���ye"��������N���z��u���H��IFJ�T�pq���+���BQ��w�gNr,��VG�����;k|���i�n9N���^G�9��<*�����m�ʬ�3t�b�2��b��%�Һ�����m��E�a��|�OL��|��i*j]� �:ڬ_�$P̓Wި>`�Y+u��'wS�I�g�x҈�/����������.������L*Ӣ���� %f_������4��ˇ�?��{=�����a[�h�2��B9��5&V�cz?��Y���?=&��t�)
Ss`�>!��w8�ݠ�eF}B�'�<��8�t$[oU�yO��>NPl��a�8�5��'D�@��B�I97����/���U)j��CzC���~���F�e��=:|�u����20�Q�7�^`%��d�K���8ܻL͘(`�M���A���Gn�ܭ4�P��E�@��LM��W(��,�K���=f�rEx_6��ή7���O\�,�iax(/�g7Z��LNV�����D�'N�z惧�s"�4�K8l���=u{��(��bO�+�'��s.uk�՘���Q���0�}����b������T\��LsY���c�deI���E��tQ�p/�PP�@Ķ�����r<^;;��-�����8Zs!n��9�yq㇛���θ�Z�P���F��J�j��\��	pxj@h���G�8���A`(i����)�i���C��{,�/;W���~����Nҩ+?�k6�c�q�Z,�O�9/MQ�R���ҧ��̃aR�(ʡ�����3Ev�b٧:�������V�=)��/q?[d�x�.j��N���W���@��#B�!��;��ȋ�IA���H~�1ΦU���^	Ӯ�yq9�F�~ G���4�,AJ��|,M�a�X2��8�%%�[qK��n��W�֛`?�K�-�ΰ�m�ڠ����)�dyL�[�`��*1Ql�����Z�ĺ
ܻtl����a<��[W���W�F�y\����0o?ln�ͿL��$7����aTlV�"�\u ^O����R%Ŵ;����?���H��|e�.3�A�Ig�ѳmf];�r�u{V����}�}x�{��c�9n�ک�e5��<��&֥1� qM�P2d�{��b"|��3���.<
3����jb	��k\��Ma����q��ʨi�m@w\��&� &lT3H�RTE�#%��7����Lx.4�m�%�)L�3�@g.�c/��~[B�cKi��Iɗ��.��L�T��e�	�}B�!/P}���9��@%޼M���<}R��I�	��^.�EHF#�!�ׅ��O���ٺ�Ʃ�\ʍ*��QPd"�,l��ء��A���-K�u���~y��"����x���� ��˳��W<#����z��F�d��d�,�a��"`�e��f��d^�԰��E�'���ʑ�Ƿ�o�&��y��DED)�CA|⚺$�v�j �t>]ʋ�����
ʚi:_��J��VbWhsl�P�\��ɲ����n�d ��Fg�:�_z��Dp���>��3��Ȝ�S����B�b�@��Xf���_E���`n��W4$�ԲI^��!��*I�) >Ú��s;�&?S�����*p[�܊��iW�JkeVT+ج#�"��i8��o1��]z7V�f��!/[�4}��$��L ����+�D{���y��"��9ʂ�ݖ>���$}����V
� (6