��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_}���l�'���(p��9��^P�m$n��B�`~�^�%�L˲�|���P�G |9k�?�{;]n.�V[��CG�32�E��2��%���4�T����u'�c�}��>�)iXf��#O�Ⱥ}�R�m�4�4��zm�3����������F�yn5�Fo�Ұ��k<�ml::S�~�~�;���P��V�we�3����`���0�A�"أ����I�1�FL��^<�ͱ�n�-�3�O�Qb�J�����6���I8@W�>�`�ܭ�fƊ��ח'[�L�p$�s�ĸL�ě�
=" ����3F��E��q_�:�����̳���
b��#�?�:��I��z����l��8V�������n4���G1��+��C=:+ �K�$��Y�rs+{�U������v����?szۼl� ���-��i�������`*�R�K4�㼨����_
lGJI�׸���Z��|F�M�3�.�������(�ėl��	�D�L�X��"Q��M,sJ�J��=+���e�sn������|�jo����KE�dP�q� -��a�9c8�|�2-��蝡����D�vo�@5HN�[�����È��+ˡz�+���Ic�-w�f��]�^Tѳ���z�HQ�y����JO8��Md�r��
�s��(�W,ǜ4AZ��Oh�Ky���~��x%b��VލJT�N�����/�֣��O|E�p�;�<}=&�ǳ��2Q��ChX��>�$?x���8h>�)�GON�k��b�6'RvH|s��*L��$)���ؑ ����^�pQ��YVp�z;������j��;t���� �����(4�}@�{�� VC�Q`)ۻ�' �I\;��F���g�2�%�f*��g�����T�
�8�m��`]�O ��jX�6ae�E�)2�����\IȀtgî퐦��}H�q�R�M�����,�k��
��'SŚ����U�*?,�Wj�i9���tN%� ɥ�{��;��EL�f��) 3��`��x�\r���� ���$B�3�h�O��I��	w�����Yci4%<`<���E�vY+1��`#��YA���4����ࠚ"�u �xp��2�]��R�D�W�o\�ȁ&t��ݶ~��n��=�!iD��Ζߎ���_���M����fz��QO�-���ƹ�·�3ۊ�ܵh���c�8w�Ѓ��_���N�m�t`'�H�Hޠ�?jVo-�Z�n.���r�gt�l�+�>���=�)�p`@&\Я���-&��9q�K��p3���ס���Qc�����1��W�v��?��[�/M�Y���ۆ��9�q�h6�2��e�uY����c����i4Arݬ�ޘ�fÌPZ���H�N:�����n�5�	�wG
_����\f��_��:��%��Dz#1vd���e-�?���T�J���Z�ֵ�&�]��nח4����
�դP%���7�2��?�=��n#,��Ό1Da��M���ܔi�Ռ*;~v�X2k��s#�$\#��Ծ�Q���� 2G�DvL��������~��2n��t�͉(]�wm����<A���������h�g���`�\\`?6\xx- +�/:���a�x*�����7�Ѥ�4��w�"c��kG������e��	���-k�	6+`�q�+G���΅�I�0x�g�C�D(YN�r�i�i��9Iҹu��$i�+���۷���RPx�$�mh�g�5=w�xSg��ŏ^���:�cޟ��Y�吕���%��w��d]�)�=X�9��X�y���9��`����zy5�&��*0{%qt�2j���w�i���
����F���B]p͓�P(��:����~٭�꭯fɬڃ�R�Gő�(��}�5�xl�t��ju#L+�KL-�.��޼�}�>���e=$��^�*��& �s]ͅ4.���r�S�M��Zm��	�ð#c�ېA��U�j���L
��q�9��gBل���? 8�CJ������(��:�M��:7gw@��w��/�`��EC�O�`���Q���	��R��'Nu-e�ͻ��!�_Ix�#ᛪ,��=M"��+A��&���:�o��c��m�h3wK�w��P(�����̨f������0.������1�W)�b�`e��F�}M|8��v95A�B�/*�Z)�ћ_���Lpӈ�ڀ ǥf%�3|��[n#&��R���ZX�.b�����B5&�zHib�F`.A�6f�8+(p��[s��U'u�D�l����z4��/x/�8z�*���{���uz��;>�����
�B*�aUD��rO�V˨p6����OP���|>��&7��Ac��R���	C���2Kc��̬�:���)B�1���1�aU�^�Ψe@g_�` ������TH���a�7�f�R�lG�;���Ӕ`E�H��,�����b�d'���8j��i�e�G�(Upܖd�{>|�sN�ESF7��C���A�w����hǯ'��r+x��Hݹ�o��,W܍�D-�����M�60#��߹�X ���_��4��uY�}���X����/����1O�7>�k��d`� t�w��A#������f��x��8���p����Έ��/�g��z�.��桚^�&��cNܐ�4S�QD�a[�*�[�8ʉW�p*Y*PGu$���o֜mD����6jh�����{)Y*dT�Qu�f��a������"e�6`�$1xAd����<�B�-����������E��(��&�򿪵/�������G�V���C*�х�|�u���H;�D��B	܉� �}	eLa�f��s�/	H�~AxAb6箷u�kc�;��O�&��<@��s����v�����i9���	�'e��h������t��� 
vD��KqWeG1�Y�[��2Z�x���L�̪~+�8N񛀈#�����.�I0��A,<A�y+�Z�_a{�z"�_m53RٟA��x*?x��]r��0R��Y�EfC�,�u�x��=oT��dV�)$�$W��ۙ�?����LN61s��Dsr����N����q�Y����d��Rr67���ȕ�9~�'м~O�xW�
t�X�Q��__.a��0�2G{�������9L	4�K�c��J�����ס@AFf����d����j����2_qz��aǭ	�
o��l��*f�'������(�q���ފ�ݧ)�e��f2�{斍�W_�s�Wط����r�v�'�&�UӍG��q;{��O�G[��3^��
�&�FAJu�c/z4�N�i>��a�����:i�����,tA�����Ja�0T��-;*�&xY�k�
�X�z�д����_ڳ,�;�|j��dK�=⫯�<I?~�7��y�1R&{�-���ޡ�6SW����/[��E�,�w�@ b�I�Sb����8q�Eo�:stA�sX���	�����>�Z�怪����c4Y���0|T4椠�ui~w�d�B�A�����Z��t��`cc�;{��G^���h�o�4tg"�\��A�ka	�un����lbW��?�gg��o����p��]�=�����TU�M(o�Ġ���g��#���w�o��W߈��8ݘ#�L<ƻ�"��!"9��>��:T+�[!�%�9q7���f��۾�*a��.s�L=���y�x̀q\5F�4�qYf�Y����7���}V�r�O.!:��L�|��9gU�4���Wl�fG���+��!�������$�"~SY}��T��@��pg�6��3�uI���*���zN��D|��Qt^o�p����6r���v���0	6����İ���)Ϩ2pL�L�ʳ�O�������sd�U����}|]t�l�����J�hD����V���K��J;��1"-t�sy�Z�$\#������+�"oڜ3���	�\N��k���y'+=ҳ�4����|4k�W�}�)6cT��|T���ΞЩ�?�JG�x���p�{V{F�����V~�H�
5ё r��p�V��O�����Ӈ���n�S4�)d��S��Xi���^����!s)��^�o�0��qS��*0���(m�>u��|;�n#G�F0�-_i��ċ�4.�#w��O���c㥿"ӌ�I5v���\�f&��;+x�������O�<�J�#{�o�Oh�&�
����}r��P���g( ��?>��PĲ� ��N��j(R��(gO� ˧e���Ļ&+n�n�Q�+�?�B�g��N%=���l���X�<�����S�Z�w�����%�9t��ޫR��Z���⍊�[�~!�6h�C)	W�m�0�	bo7�U���^�����!�oz�'-'�X���hCO���d2���Jn�d: Q0�r�������B,1��φ�+2���I}?���+bS��C m�O�<ة����$JӢ������u�� =�5򭫡�^�����%�*�*����BO,��E>K�˦e5p�4U4�.�o��8I�g6*3���M"���O7�S���F7ӛ��}�n�.�\�o}-3q9�s�����Vi�������)F}��Aj �㤃�5ITZ�q�]�IN���H3�
�n�e���!d����n����<�}I=�
�2'�g5 �:N*+�(��4�*#��r�U)"��Y���d�c�u�3�
�X�&�����fU�%�#dv9TA�h�����p6�wC��C"9~��k�(�&Y ��&#Hb��Iٴd<��\0�\�`0���c/_�u�؇l2��$���f(�.�-�ث�K	//��'���UN�-9 ��vfvTv4����:��	��2�0D*�5�3�����
4��/�0R�\)
Pq}N�&CZ-�Y����` �_��Q��e��������G{@[	��H���(��b[`�U-�H�tq�ì ���G�AD�v�-0�5;���G