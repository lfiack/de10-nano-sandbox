library ieee;
use ieee.std_logic_1164.all;

entity dpram is
    generic
    (
        mem_size    : natural := 720 * 480;
        data_width  : natural := 8
    );
   port 
   (   
        i_clk_a        : in std_logic;
        i_clk_b        : in std_logic;

       i_data_a    : in std_logic_vector(data_width-1 downto 0);
       i_data_b    : in std_logic_vector(data_width-1 downto 0);
       i_addr_a    : in natural range 0 to mem_size-1;
       i_addr_b    : in natural range 0 to mem_size-1;
       i_we_a      : in std_logic := '1';
       i_we_b      : in std_logic := '1';
       o_q_a       : out std_logic_vector(data_width-1 downto 0);
       o_q_b       : out std_logic_vector(data_width-1 downto 0)
   );
   
end dpram;

architecture rtl of dpram is
    -- Build a 2-D array type for the RAM
    subtype word_t is std_logic_vector(data_width-1 downto 0);
    type memory_t is array(0 to mem_size-1) of word_t;
    
    -- Declare the RAM
    shared variable ram : memory_t := (
        x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"60", x"5f", x"5f", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"61", 
        x"61", x"61", x"62", x"62", x"61", x"61", x"62", x"62", x"61", x"60", x"60", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"61", 
        x"61", x"61", x"60", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"63", x"63", x"62", 
        x"62", x"62", x"61", x"60", x"61", x"61", x"61", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"61", x"61", 
        x"62", x"63", x"64", x"64", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"61", x"63", x"65", x"62", 
        x"60", x"63", x"61", x"62", x"61", x"60", x"61", x"63", x"63", x"63", x"63", x"64", x"63", x"63", x"63", 
        x"62", x"63", x"63", x"64", x"64", x"63", x"63", x"62", x"63", x"62", x"62", x"62", x"63", x"62", x"62", 
        x"63", x"64", x"62", x"63", x"64", x"65", x"64", x"63", x"63", x"64", x"64", x"64", x"64", x"65", x"65", 
        x"64", x"64", x"64", x"65", x"65", x"65", x"65", x"64", x"63", x"64", x"64", x"64", x"64", x"64", x"64", 
        x"62", x"62", x"64", x"66", x"66", x"64", x"62", x"61", x"61", x"65", x"64", x"63", x"64", x"62", x"63", 
        x"62", x"62", x"65", x"65", x"62", x"64", x"65", x"64", x"63", x"63", x"64", x"64", x"64", x"66", x"67", 
        x"66", x"65", x"67", x"6a", x"6b", x"68", x"64", x"65", x"67", x"66", x"64", x"64", x"68", x"66", x"64", 
        x"64", x"66", x"66", x"64", x"64", x"66", x"69", x"67", x"64", x"64", x"66", x"66", x"66", x"66", x"64", 
        x"63", x"64", x"65", x"68", x"65", x"66", x"67", x"67", x"68", x"68", x"65", x"65", x"66", x"66", x"65", 
        x"66", x"66", x"66", x"66", x"67", x"67", x"67", x"67", x"66", x"65", x"65", x"68", x"67", x"65", x"65", 
        x"67", x"68", x"66", x"65", x"63", x"64", x"66", x"65", x"65", x"66", x"66", x"66", x"66", x"66", x"65", 
        x"66", x"66", x"69", x"69", x"67", x"66", x"68", x"6a", x"68", x"66", x"66", x"67", x"67", x"65", x"64", 
        x"64", x"65", x"67", x"6a", x"6a", x"67", x"67", x"67", x"69", x"66", x"66", x"66", x"68", x"67", x"67", 
        x"6a", x"6a", x"68", x"6a", x"6b", x"67", x"68", x"6a", x"6a", x"67", x"68", x"66", x"64", x"66", x"66", 
        x"65", x"66", x"67", x"67", x"66", x"68", x"68", x"67", x"69", x"69", x"67", x"65", x"64", x"68", x"69", 
        x"64", x"62", x"65", x"66", x"66", x"68", x"68", x"66", x"65", x"65", x"67", x"69", x"69", x"68", x"67", 
        x"66", x"66", x"67", x"65", x"64", x"63", x"67", x"67", x"65", x"65", x"66", x"64", x"64", x"66", x"65", 
        x"65", x"66", x"66", x"65", x"65", x"67", x"69", x"67", x"66", x"66", x"66", x"65", x"66", x"67", x"64", 
        x"67", x"66", x"67", x"68", x"67", x"64", x"64", x"65", x"66", x"66", x"65", x"64", x"67", x"65", x"67", 
        x"67", x"66", x"66", x"66", x"69", x"69", x"68", x"67", x"66", x"66", x"69", x"68", x"63", x"64", x"68", 
        x"67", x"66", x"67", x"65", x"64", x"64", x"64", x"64", x"64", x"64", x"65", x"64", x"63", x"63", x"64", 
        x"66", x"67", x"66", x"66", x"67", x"67", x"66", x"67", x"69", x"69", x"6a", x"66", x"65", x"67", x"66", 
        x"66", x"66", x"67", x"68", x"66", x"65", x"65", x"65", x"66", x"67", x"66", x"62", x"61", x"64", x"65", 
        x"64", x"66", x"67", x"67", x"66", x"66", x"66", x"66", x"66", x"66", x"62", x"63", x"66", x"66", x"66", 
        x"64", x"65", x"64", x"67", x"66", x"64", x"65", x"64", x"63", x"64", x"69", x"6a", x"67", x"64", x"65", 
        x"64", x"61", x"62", x"62", x"61", x"61", x"62", x"63", x"62", x"62", x"63", x"63", x"63", x"64", x"64", 
        x"62", x"65", x"66", x"65", x"62", x"61", x"62", x"65", x"62", x"61", x"63", x"65", x"65", x"68", x"65", 
        x"63", x"62", x"62", x"64", x"64", x"65", x"65", x"65", x"65", x"66", x"64", x"62", x"62", x"62", x"64", 
        x"64", x"62", x"63", x"64", x"64", x"62", x"63", x"63", x"60", x"64", x"66", x"64", x"63", x"64", x"65", 
        x"65", x"64", x"62", x"62", x"62", x"62", x"64", x"62", x"63", x"64", x"64", x"63", x"62", x"65", x"65", 
        x"62", x"61", x"62", x"64", x"64", x"64", x"64", x"64", x"62", x"61", x"61", x"61", x"63", x"63", x"61", 
        x"61", x"61", x"63", x"64", x"63", x"61", x"61", x"61", x"62", x"61", x"61", x"62", x"62", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"63", x"62", x"61", x"61", x"61", x"61", x"62", x"63", x"62", x"61", x"61", 
        x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"62", x"62", x"62", x"61", x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"60", x"60", x"60", x"61", x"61", x"5f", x"5f", x"5f", x"60", x"60", x"61", x"61", 
        x"60", x"60", x"60", x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5f", x"5f", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", 
        x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", 
        x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"60", x"5f", x"5f", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"60", x"60", x"5f", 
        x"5f", x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"62", x"62", x"62", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"62", 
        x"62", x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"61", 
        x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"62", x"64", x"64", x"64", x"63", x"62", x"61", x"61", x"61", x"61", x"62", x"62", x"64", x"65", x"62", 
        x"60", x"62", x"62", x"61", x"61", x"60", x"61", x"62", x"63", x"64", x"64", x"64", x"63", x"62", x"61", 
        x"61", x"62", x"63", x"64", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"64", x"63", x"63", 
        x"63", x"63", x"62", x"62", x"63", x"64", x"64", x"63", x"64", x"64", x"64", x"65", x"65", x"66", x"66", 
        x"66", x"65", x"65", x"64", x"64", x"63", x"63", x"62", x"63", x"64", x"64", x"64", x"64", x"65", x"65", 
        x"63", x"63", x"63", x"65", x"66", x"65", x"64", x"63", x"63", x"66", x"65", x"64", x"63", x"61", x"64", 
        x"63", x"63", x"64", x"63", x"63", x"64", x"65", x"63", x"62", x"62", x"65", x"66", x"66", x"67", x"68", 
        x"66", x"63", x"65", x"68", x"68", x"66", x"66", x"66", x"68", x"67", x"65", x"66", x"69", x"68", x"66", 
        x"65", x"66", x"67", x"65", x"63", x"65", x"69", x"68", x"65", x"65", x"66", x"65", x"65", x"65", x"65", 
        x"65", x"65", x"66", x"67", x"65", x"66", x"68", x"66", x"66", x"66", x"63", x"64", x"66", x"66", x"66", 
        x"66", x"66", x"66", x"65", x"64", x"65", x"65", x"65", x"65", x"65", x"64", x"66", x"66", x"64", x"64", 
        x"67", x"69", x"67", x"67", x"65", x"65", x"67", x"66", x"65", x"68", x"67", x"67", x"67", x"67", x"67", 
        x"68", x"68", x"68", x"68", x"67", x"66", x"67", x"68", x"6a", x"68", x"65", x"67", x"67", x"66", x"65", 
        x"65", x"66", x"67", x"6a", x"6a", x"68", x"67", x"68", x"69", x"68", x"66", x"67", x"68", x"66", x"66", 
        x"69", x"68", x"66", x"6a", x"69", x"66", x"69", x"69", x"67", x"66", x"68", x"67", x"67", x"68", x"68", 
        x"68", x"68", x"67", x"65", x"66", x"69", x"68", x"66", x"68", x"67", x"66", x"66", x"66", x"66", x"66", 
        x"65", x"64", x"67", x"69", x"67", x"67", x"68", x"69", x"67", x"67", x"68", x"68", x"66", x"64", x"67", 
        x"69", x"69", x"68", x"67", x"65", x"64", x"66", x"67", x"67", x"67", x"66", x"65", x"65", x"66", x"67", 
        x"67", x"67", x"66", x"66", x"65", x"65", x"67", x"66", x"66", x"67", x"68", x"67", x"67", x"67", x"67", 
        x"69", x"64", x"65", x"69", x"68", x"64", x"66", x"66", x"65", x"66", x"67", x"64", x"66", x"66", x"68", 
        x"68", x"67", x"66", x"68", x"6a", x"69", x"69", x"69", x"67", x"66", x"66", x"67", x"65", x"66", x"6a", 
        x"69", x"66", x"65", x"64", x"63", x"62", x"64", x"67", x"67", x"67", x"69", x"66", x"64", x"64", x"66", 
        x"68", x"68", x"67", x"66", x"65", x"65", x"65", x"66", x"65", x"66", x"68", x"65", x"65", x"68", x"66", 
        x"65", x"65", x"64", x"65", x"65", x"65", x"67", x"69", x"69", x"68", x"66", x"61", x"62", x"65", x"66", 
        x"65", x"65", x"66", x"66", x"65", x"65", x"65", x"65", x"65", x"64", x"62", x"61", x"64", x"67", x"67", 
        x"65", x"64", x"64", x"67", x"65", x"65", x"64", x"64", x"64", x"64", x"67", x"67", x"64", x"64", x"66", 
        x"65", x"63", x"63", x"63", x"62", x"62", x"63", x"64", x"62", x"62", x"63", x"63", x"63", x"64", x"63", 
        x"62", x"64", x"66", x"65", x"62", x"62", x"64", x"64", x"63", x"62", x"63", x"65", x"67", x"66", x"66", 
        x"64", x"61", x"61", x"65", x"65", x"63", x"62", x"63", x"62", x"62", x"62", x"63", x"64", x"65", x"64", 
        x"63", x"63", x"64", x"64", x"64", x"63", x"65", x"65", x"61", x"64", x"67", x"64", x"62", x"64", x"65", 
        x"66", x"64", x"63", x"63", x"63", x"63", x"63", x"63", x"64", x"63", x"62", x"61", x"61", x"63", x"65", 
        x"64", x"63", x"64", x"64", x"64", x"62", x"63", x"63", x"63", x"62", x"61", x"62", x"62", x"62", x"62", 
        x"62", x"61", x"63", x"63", x"62", x"61", x"61", x"61", x"62", x"61", x"60", x"61", x"61", x"62", x"63", 
        x"63", x"63", x"62", x"64", x"63", x"62", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"62", x"62", 
        x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"61", x"61", 
        x"61", x"62", x"61", x"60", x"60", x"61", x"61", x"62", x"61", x"61", x"60", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"5f", x"5f", x"5f", x"5f", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5f", x"5f", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", 
        x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", 
        x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"60", x"5f", x"5f", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"60", x"60", x"5f", 
        x"5f", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"61", x"61", x"62", 
        x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"61", x"62", 
        x"61", x"60", x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", 
        x"61", x"62", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"63", x"62", x"62", x"62", 
        x"63", x"63", x"64", x"63", x"62", x"62", x"61", x"61", x"61", x"62", x"63", x"63", x"64", x"65", x"61", 
        x"5f", x"61", x"62", x"61", x"61", x"62", x"62", x"62", x"63", x"64", x"64", x"64", x"62", x"61", x"61", 
        x"61", x"62", x"63", x"64", x"63", x"63", x"63", x"64", x"63", x"62", x"63", x"64", x"64", x"63", x"62", 
        x"62", x"64", x"62", x"61", x"62", x"64", x"64", x"64", x"64", x"63", x"63", x"65", x"66", x"66", x"65", 
        x"64", x"64", x"64", x"64", x"64", x"63", x"64", x"63", x"63", x"64", x"64", x"64", x"64", x"65", x"65", 
        x"64", x"63", x"63", x"64", x"65", x"65", x"64", x"62", x"62", x"66", x"65", x"65", x"65", x"63", x"65", 
        x"64", x"63", x"63", x"62", x"64", x"65", x"64", x"62", x"62", x"63", x"66", x"67", x"67", x"65", x"66", 
        x"65", x"64", x"66", x"69", x"68", x"66", x"67", x"66", x"67", x"66", x"66", x"68", x"68", x"66", x"65", 
        x"65", x"66", x"68", x"68", x"65", x"64", x"68", x"68", x"65", x"66", x"65", x"64", x"65", x"64", x"65", 
        x"66", x"66", x"67", x"66", x"65", x"68", x"69", x"66", x"64", x"64", x"63", x"63", x"64", x"65", x"66", 
        x"67", x"67", x"67", x"66", x"65", x"65", x"65", x"65", x"64", x"63", x"63", x"66", x"66", x"65", x"64", 
        x"66", x"66", x"65", x"68", x"67", x"66", x"66", x"65", x"66", x"68", x"65", x"64", x"65", x"66", x"66", 
        x"67", x"67", x"64", x"63", x"65", x"66", x"64", x"65", x"68", x"68", x"66", x"67", x"67", x"67", x"67", 
        x"68", x"67", x"68", x"69", x"6a", x"68", x"66", x"69", x"6a", x"6a", x"68", x"68", x"68", x"66", x"66", 
        x"67", x"67", x"68", x"69", x"68", x"68", x"6c", x"6b", x"66", x"65", x"67", x"67", x"6a", x"6a", x"68", 
        x"68", x"67", x"68", x"67", x"67", x"69", x"68", x"68", x"68", x"67", x"66", x"67", x"67", x"63", x"62", 
        x"66", x"67", x"67", x"69", x"68", x"67", x"69", x"69", x"68", x"67", x"67", x"68", x"67", x"67", x"68", 
        x"6a", x"6a", x"69", x"68", x"67", x"64", x"65", x"67", x"69", x"69", x"66", x"67", x"66", x"68", x"6a", 
        x"69", x"67", x"65", x"65", x"64", x"65", x"69", x"67", x"68", x"68", x"67", x"65", x"65", x"65", x"69", 
        x"6a", x"62", x"64", x"67", x"67", x"66", x"68", x"67", x"65", x"66", x"67", x"66", x"67", x"66", x"67", 
        x"66", x"66", x"66", x"68", x"68", x"66", x"68", x"69", x"68", x"66", x"66", x"68", x"68", x"67", x"6b", 
        x"69", x"65", x"64", x"64", x"66", x"63", x"66", x"69", x"68", x"67", x"6a", x"6b", x"69", x"67", x"69", 
        x"68", x"66", x"65", x"65", x"65", x"66", x"66", x"64", x"63", x"63", x"65", x"64", x"65", x"68", x"66", 
        x"67", x"67", x"67", x"68", x"68", x"66", x"67", x"67", x"66", x"65", x"64", x"61", x"64", x"65", x"66", 
        x"66", x"66", x"69", x"69", x"68", x"66", x"65", x"65", x"65", x"68", x"68", x"65", x"65", x"67", x"66", 
        x"64", x"63", x"64", x"67", x"65", x"65", x"65", x"64", x"66", x"66", x"64", x"62", x"61", x"64", x"66", 
        x"66", x"64", x"65", x"64", x"63", x"63", x"64", x"65", x"62", x"62", x"63", x"63", x"63", x"64", x"63", 
        x"62", x"64", x"65", x"64", x"63", x"63", x"65", x"63", x"64", x"65", x"64", x"66", x"67", x"63", x"65", 
        x"65", x"63", x"63", x"63", x"63", x"63", x"62", x"63", x"62", x"62", x"63", x"63", x"63", x"63", x"64", 
        x"62", x"63", x"65", x"65", x"64", x"64", x"65", x"64", x"61", x"63", x"65", x"62", x"61", x"63", x"65", 
        x"66", x"65", x"64", x"64", x"64", x"64", x"64", x"66", x"65", x"64", x"62", x"61", x"61", x"63", x"66", 
        x"65", x"64", x"64", x"63", x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"63", x"62", x"62", x"63", 
        x"63", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"62", x"61", x"61", x"61", x"62", x"62", x"64", 
        x"63", x"62", x"61", x"63", x"64", x"62", x"62", x"61", x"61", x"62", x"61", x"61", x"62", x"63", x"64", 
        x"63", x"62", x"62", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"62", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"62", x"62", x"62", x"61", x"61", x"60", x"60", x"62", x"62", x"61", x"61", x"61", x"61", 
        x"61", x"62", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"61", x"60", x"60", x"60", x"60", 
        x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5f", x"5f", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", 
        x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"60", x"61", x"62", 
        x"62", x"62", x"63", x"63", x"63", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"61", x"61", 
        x"61", x"60", x"60", x"5f", x"5f", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"63", x"62", x"61", 
        x"61", x"62", x"61", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"63", x"63", x"63", x"62", 
        x"63", x"63", x"62", x"62", x"61", x"61", x"62", x"63", x"63", x"63", x"63", x"62", x"63", x"64", x"61", 
        x"60", x"62", x"62", x"61", x"62", x"64", x"63", x"62", x"63", x"62", x"62", x"62", x"62", x"62", x"63", 
        x"63", x"64", x"64", x"64", x"63", x"63", x"63", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", 
        x"64", x"65", x"63", x"61", x"62", x"64", x"65", x"66", x"64", x"63", x"63", x"64", x"66", x"65", x"64", 
        x"64", x"64", x"64", x"65", x"65", x"65", x"65", x"65", x"65", x"64", x"64", x"64", x"64", x"64", x"64", 
        x"64", x"63", x"63", x"63", x"64", x"64", x"63", x"63", x"62", x"65", x"65", x"65", x"67", x"65", x"66", 
        x"63", x"64", x"63", x"63", x"65", x"64", x"64", x"64", x"64", x"64", x"64", x"66", x"66", x"69", x"69", 
        x"66", x"66", x"66", x"66", x"66", x"65", x"67", x"67", x"65", x"64", x"66", x"69", x"68", x"69", x"69", 
        x"66", x"65", x"66", x"65", x"63", x"64", x"67", x"67", x"64", x"66", x"66", x"65", x"66", x"64", x"66", 
        x"67", x"67", x"69", x"66", x"66", x"69", x"69", x"66", x"65", x"67", x"67", x"66", x"65", x"65", x"66", 
        x"67", x"67", x"65", x"65", x"68", x"68", x"68", x"68", x"67", x"67", x"66", x"66", x"67", x"68", x"67", 
        x"65", x"64", x"64", x"64", x"66", x"68", x"68", x"68", x"67", x"66", x"63", x"64", x"64", x"65", x"66", 
        x"65", x"65", x"64", x"63", x"65", x"67", x"66", x"65", x"67", x"68", x"67", x"67", x"67", x"68", x"69", 
        x"6a", x"69", x"68", x"69", x"69", x"6a", x"68", x"6c", x"6a", x"67", x"68", x"68", x"67", x"66", x"64", 
        x"64", x"69", x"6a", x"69", x"6a", x"6d", x"6d", x"6b", x"67", x"67", x"67", x"66", x"6a", x"69", x"67", 
        x"6b", x"6b", x"69", x"69", x"67", x"66", x"64", x"66", x"68", x"68", x"67", x"67", x"68", x"64", x"65", 
        x"67", x"68", x"66", x"68", x"69", x"68", x"6a", x"65", x"65", x"65", x"66", x"68", x"6a", x"6c", x"67", 
        x"68", x"69", x"67", x"67", x"66", x"63", x"66", x"66", x"67", x"6a", x"67", x"67", x"68", x"68", x"6a", 
        x"69", x"65", x"63", x"65", x"66", x"65", x"66", x"67", x"67", x"68", x"67", x"67", x"67", x"68", x"6a", 
        x"68", x"65", x"67", x"67", x"66", x"67", x"68", x"68", x"66", x"66", x"66", x"65", x"67", x"66", x"66", 
        x"64", x"66", x"67", x"67", x"68", x"67", x"67", x"67", x"67", x"66", x"68", x"6a", x"68", x"67", x"6a", 
        x"68", x"67", x"68", x"68", x"68", x"64", x"66", x"6a", x"6a", x"69", x"6d", x"6c", x"69", x"6a", x"6b", 
        x"68", x"65", x"66", x"66", x"67", x"69", x"6a", x"67", x"65", x"67", x"68", x"69", x"68", x"66", x"65", 
        x"65", x"67", x"68", x"68", x"69", x"68", x"68", x"68", x"68", x"66", x"63", x"62", x"67", x"66", x"64", 
        x"67", x"68", x"6a", x"69", x"68", x"67", x"66", x"66", x"66", x"66", x"6a", x"68", x"67", x"6a", x"69", 
        x"67", x"65", x"66", x"67", x"65", x"66", x"65", x"64", x"65", x"65", x"66", x"65", x"63", x"63", x"66", 
        x"65", x"62", x"62", x"62", x"63", x"63", x"62", x"62", x"63", x"63", x"63", x"63", x"63", x"63", x"63", 
        x"64", x"64", x"65", x"64", x"64", x"64", x"64", x"63", x"65", x"66", x"66", x"66", x"66", x"64", x"65", 
        x"64", x"64", x"64", x"62", x"63", x"63", x"64", x"66", x"65", x"64", x"64", x"63", x"61", x"62", x"65", 
        x"63", x"63", x"65", x"64", x"63", x"64", x"66", x"66", x"64", x"65", x"66", x"63", x"64", x"65", x"65", 
        x"66", x"65", x"64", x"64", x"65", x"64", x"64", x"67", x"65", x"64", x"64", x"63", x"63", x"64", x"65", 
        x"65", x"65", x"66", x"65", x"63", x"64", x"63", x"62", x"62", x"62", x"63", x"64", x"64", x"64", x"64", 
        x"63", x"62", x"62", x"63", x"63", x"62", x"62", x"62", x"61", x"61", x"61", x"62", x"62", x"63", x"65", 
        x"64", x"61", x"60", x"63", x"64", x"63", x"63", x"61", x"62", x"63", x"62", x"62", x"63", x"63", x"64", 
        x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"63", x"63", x"62", x"62", x"61", 
        x"61", x"61", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"62", x"62", x"62", x"61", x"60", x"61", x"62", x"62", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"60", x"60", x"60", 
        x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5f", x"5f", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5f", x"5f", x"5f", x"5d", x"5d", x"5e", 
        x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", x"5e", 
        x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"62", x"60", x"60", x"61", x"61", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"61", 
        x"62", x"62", x"63", x"64", x"64", x"62", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"61", 
        x"61", x"61", x"61", x"60", x"5f", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"61", 
        x"62", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"63", x"63", x"62", 
        x"62", x"61", x"61", x"61", x"60", x"61", x"63", x"65", x"65", x"62", x"61", x"60", x"62", x"64", x"62", 
        x"62", x"64", x"63", x"61", x"62", x"65", x"64", x"62", x"63", x"63", x"62", x"63", x"62", x"62", x"62", 
        x"62", x"64", x"65", x"64", x"63", x"63", x"64", x"64", x"64", x"65", x"64", x"63", x"64", x"64", x"65", 
        x"65", x"65", x"63", x"62", x"62", x"64", x"66", x"66", x"65", x"63", x"62", x"64", x"65", x"65", x"64", 
        x"66", x"67", x"67", x"66", x"66", x"65", x"65", x"66", x"66", x"64", x"64", x"65", x"65", x"64", x"63", 
        x"63", x"64", x"64", x"65", x"64", x"62", x"62", x"65", x"64", x"66", x"65", x"65", x"67", x"65", x"65", 
        x"64", x"65", x"64", x"64", x"66", x"64", x"62", x"63", x"64", x"64", x"64", x"66", x"66", x"62", x"63", 
        x"61", x"60", x"66", x"67", x"67", x"64", x"67", x"68", x"64", x"64", x"66", x"6a", x"66", x"66", x"67", 
        x"66", x"65", x"67", x"66", x"64", x"65", x"66", x"66", x"62", x"66", x"67", x"67", x"67", x"64", x"66", 
        x"67", x"67", x"69", x"67", x"68", x"6b", x"6a", x"67", x"65", x"66", x"67", x"67", x"66", x"66", x"67", 
        x"68", x"68", x"65", x"64", x"65", x"67", x"67", x"67", x"68", x"68", x"67", x"64", x"67", x"6a", x"6a", 
        x"67", x"65", x"66", x"65", x"67", x"67", x"66", x"68", x"6a", x"68", x"65", x"66", x"67", x"67", x"67", 
        x"66", x"65", x"67", x"67", x"67", x"6a", x"6b", x"69", x"69", x"69", x"67", x"66", x"67", x"69", x"6b", 
        x"6b", x"6b", x"6d", x"6b", x"6a", x"6b", x"69", x"6b", x"6a", x"6b", x"6b", x"68", x"66", x"67", x"68", 
        x"67", x"67", x"66", x"65", x"69", x"6c", x"66", x"65", x"67", x"67", x"66", x"65", x"6a", x"69", x"68", 
        x"6c", x"68", x"63", x"64", x"69", x"6a", x"6a", x"68", x"66", x"68", x"68", x"66", x"68", x"68", x"69", 
        x"68", x"6b", x"67", x"67", x"68", x"67", x"67", x"66", x"67", x"67", x"67", x"67", x"67", x"68", x"67", 
        x"69", x"6a", x"68", x"68", x"67", x"65", x"69", x"66", x"64", x"69", x"69", x"69", x"69", x"69", x"69", 
        x"67", x"64", x"62", x"65", x"67", x"66", x"67", x"67", x"67", x"66", x"67", x"67", x"68", x"6b", x"6a", 
        x"68", x"68", x"6b", x"67", x"66", x"66", x"66", x"67", x"67", x"67", x"65", x"64", x"67", x"67", x"66", 
        x"63", x"65", x"68", x"67", x"68", x"69", x"6a", x"6a", x"69", x"67", x"67", x"68", x"68", x"67", x"69", 
        x"67", x"67", x"69", x"6a", x"6c", x"67", x"66", x"69", x"68", x"68", x"6a", x"68", x"66", x"69", x"6b", 
        x"68", x"66", x"67", x"66", x"66", x"6a", x"6b", x"67", x"65", x"68", x"69", x"6b", x"6a", x"65", x"64", 
        x"65", x"68", x"69", x"69", x"6b", x"69", x"68", x"69", x"6a", x"68", x"64", x"64", x"68", x"66", x"64", 
        x"68", x"68", x"65", x"64", x"64", x"65", x"66", x"67", x"67", x"65", x"69", x"68", x"67", x"6a", x"67", 
        x"64", x"64", x"66", x"67", x"65", x"67", x"66", x"65", x"68", x"68", x"66", x"65", x"65", x"66", x"66", 
        x"66", x"63", x"64", x"64", x"65", x"65", x"64", x"63", x"63", x"64", x"64", x"63", x"64", x"63", x"64", 
        x"66", x"65", x"65", x"64", x"63", x"63", x"63", x"64", x"64", x"65", x"67", x"66", x"65", x"66", x"67", 
        x"64", x"62", x"64", x"64", x"66", x"65", x"63", x"65", x"64", x"63", x"65", x"66", x"66", x"66", x"67", 
        x"64", x"64", x"65", x"63", x"62", x"63", x"63", x"65", x"64", x"65", x"66", x"64", x"65", x"66", x"66", 
        x"66", x"66", x"64", x"63", x"64", x"64", x"62", x"66", x"64", x"63", x"64", x"64", x"64", x"63", x"63", 
        x"63", x"66", x"68", x"67", x"66", x"67", x"66", x"64", x"62", x"63", x"64", x"65", x"66", x"65", x"63", 
        x"62", x"61", x"62", x"63", x"62", x"63", x"63", x"62", x"62", x"62", x"63", x"62", x"60", x"61", x"65", 
        x"64", x"62", x"61", x"64", x"64", x"64", x"64", x"62", x"63", x"64", x"64", x"63", x"63", x"62", x"62", 
        x"62", x"63", x"63", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"63", x"63", x"63", x"62", x"62", 
        x"62", x"61", x"63", x"62", x"61", x"61", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"62", x"63", x"62", x"61", x"62", x"61", x"62", x"62", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"63", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5f", x"5f", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5d", x"5d", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", x"5d", x"5d", x"5d", x"5e", x"5f", x"5e", x"5d", 
        x"63", x"62", x"62", x"62", x"63", x"62", x"61", x"61", x"61", x"60", x"60", x"60", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"62", x"61", x"5f", x"61", x"62", x"60", 
        x"60", x"61", x"61", x"62", x"62", x"61", x"60", x"61", x"60", x"5f", x"61", x"62", x"61", x"62", x"62", 
        x"60", x"62", x"63", x"62", x"61", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"62", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"61", x"61", x"61", x"61", x"62", x"62", 
        x"61", x"61", x"62", x"62", x"61", x"61", x"60", x"61", x"64", x"64", x"62", x"63", x"63", x"62", x"61", 
        x"61", x"63", x"64", x"63", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", 
        x"62", x"63", x"63", x"61", x"61", x"61", x"61", x"62", x"62", x"63", x"62", x"63", x"64", x"64", x"63", 
        x"62", x"63", x"65", x"64", x"63", x"64", x"64", x"63", x"62", x"62", x"63", x"64", x"63", x"62", x"62", 
        x"63", x"64", x"64", x"64", x"64", x"64", x"64", x"63", x"62", x"63", x"63", x"63", x"66", x"66", x"68", 
        x"63", x"63", x"64", x"63", x"62", x"65", x"66", x"65", x"66", x"64", x"64", x"65", x"64", x"63", x"64", 
        x"64", x"64", x"66", x"65", x"65", x"65", x"66", x"67", x"67", x"65", x"64", x"64", x"65", x"66", x"65", 
        x"65", x"65", x"64", x"66", x"66", x"65", x"61", x"65", x"67", x"67", x"66", x"67", x"68", x"66", x"67", 
        x"65", x"64", x"64", x"64", x"66", x"64", x"65", x"63", x"66", x"65", x"65", x"63", x"5e", x"7e", x"9d", 
        x"82", x"5e", x"61", x"68", x"6a", x"69", x"68", x"69", x"67", x"67", x"68", x"6a", x"69", x"67", x"66", 
        x"67", x"67", x"67", x"64", x"65", x"66", x"66", x"66", x"65", x"64", x"63", x"63", x"66", x"65", x"64", 
        x"64", x"64", x"66", x"66", x"65", x"67", x"66", x"68", x"65", x"63", x"68", x"66", x"65", x"67", x"69", 
        x"69", x"69", x"68", x"66", x"65", x"6a", x"6a", x"66", x"67", x"69", x"66", x"65", x"6b", x"6a", x"69", 
        x"69", x"66", x"65", x"6a", x"67", x"67", x"68", x"69", x"68", x"68", x"65", x"66", x"67", x"66", x"66", 
        x"67", x"65", x"66", x"67", x"67", x"67", x"66", x"67", x"67", x"69", x"67", x"65", x"68", x"6a", x"68", 
        x"67", x"6a", x"6d", x"6b", x"6a", x"6a", x"6a", x"6b", x"6a", x"6a", x"69", x"69", x"69", x"6a", x"69", 
        x"68", x"69", x"67", x"67", x"6a", x"6a", x"67", x"67", x"69", x"6a", x"6a", x"69", x"6a", x"69", x"68", 
        x"69", x"69", x"69", x"68", x"67", x"68", x"6a", x"69", x"66", x"68", x"67", x"66", x"67", x"66", x"65", 
        x"68", x"6a", x"69", x"66", x"64", x"64", x"67", x"68", x"69", x"68", x"68", x"67", x"68", x"68", x"69", 
        x"69", x"69", x"6b", x"69", x"67", x"66", x"6a", x"6a", x"68", x"68", x"68", x"69", x"6a", x"69", x"67", 
        x"67", x"67", x"66", x"64", x"67", x"69", x"66", x"63", x"63", x"66", x"6c", x"6a", x"69", x"67", x"68", 
        x"67", x"65", x"66", x"65", x"63", x"65", x"66", x"66", x"67", x"68", x"69", x"6a", x"68", x"6a", x"67", 
        x"65", x"64", x"65", x"68", x"68", x"69", x"68", x"67", x"66", x"67", x"67", x"68", x"69", x"6a", x"6c", 
        x"69", x"66", x"68", x"6b", x"6a", x"67", x"66", x"68", x"6b", x"6a", x"67", x"67", x"67", x"69", x"69", 
        x"65", x"68", x"68", x"68", x"67", x"67", x"68", x"65", x"64", x"66", x"65", x"65", x"66", x"67", x"68", 
        x"68", x"66", x"69", x"69", x"68", x"6a", x"6a", x"67", x"68", x"6b", x"6a", x"68", x"67", x"67", x"66", 
        x"68", x"66", x"63", x"62", x"64", x"64", x"66", x"67", x"67", x"67", x"65", x"65", x"66", x"65", x"65", 
        x"61", x"64", x"66", x"66", x"67", x"69", x"68", x"67", x"65", x"65", x"66", x"68", x"68", x"64", x"62", 
        x"64", x"64", x"67", x"68", x"67", x"65", x"65", x"65", x"63", x"66", x"67", x"66", x"67", x"68", x"68", 
        x"66", x"64", x"66", x"65", x"62", x"65", x"66", x"66", x"66", x"64", x"66", x"69", x"67", x"64", x"66", 
        x"67", x"66", x"66", x"66", x"67", x"65", x"66", x"68", x"68", x"67", x"66", x"66", x"67", x"67", x"65", 
        x"64", x"64", x"65", x"62", x"61", x"65", x"64", x"65", x"64", x"67", x"66", x"66", x"65", x"67", x"64", 
        x"64", x"67", x"65", x"62", x"65", x"66", x"62", x"65", x"64", x"61", x"62", x"64", x"65", x"65", x"64", 
        x"63", x"63", x"64", x"66", x"66", x"66", x"68", x"65", x"62", x"63", x"65", x"65", x"64", x"63", x"64", 
        x"63", x"63", x"62", x"62", x"65", x"65", x"64", x"63", x"63", x"64", x"65", x"64", x"62", x"60", x"61", 
        x"62", x"62", x"61", x"61", x"62", x"64", x"63", x"61", x"61", x"62", x"63", x"62", x"62", x"62", x"62", 
        x"62", x"63", x"64", x"63", x"63", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"61", 
        x"61", x"61", x"63", x"62", x"62", x"61", x"61", x"62", x"63", x"62", x"61", x"62", x"63", x"62", x"61", 
        x"61", x"61", x"60", x"61", x"62", x"62", x"62", x"63", x"62", x"61", x"61", x"61", x"61", x"62", x"62", 
        x"62", x"62", x"62", x"63", x"63", x"63", x"62", x"62", x"62", x"61", x"61", x"61", x"60", x"60", x"60", 
        x"5f", x"60", x"5f", x"5e", x"5f", x"5f", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5f", x"5e", 
        x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5e", x"5e", x"5f", x"60", x"5f", x"5d", x"5d", 
        x"5d", x"5d", x"5d", x"5e", x"5e", x"5d", x"5e", x"5e", x"5d", x"5d", x"5d", x"5f", x"60", x"5f", x"5e", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"61", x"61", x"5f", x"61", x"63", x"61", 
        x"61", x"61", x"61", x"62", x"62", x"62", x"61", x"62", x"62", x"60", x"61", x"62", x"60", x"61", x"62", 
        x"61", x"62", x"62", x"62", x"61", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"63", x"62", x"62", 
        x"62", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"62", x"62", 
        x"61", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"63", x"63", x"61", x"62", x"63", x"62", x"61", 
        x"61", x"63", x"63", x"61", x"61", x"61", x"62", x"62", x"63", x"64", x"62", x"61", x"63", x"65", x"64", 
        x"63", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"63", x"62", x"62", x"63", x"63", x"63", x"62", 
        x"62", x"62", x"64", x"64", x"64", x"63", x"63", x"63", x"63", x"63", x"65", x"64", x"63", x"62", x"62", 
        x"62", x"63", x"65", x"64", x"64", x"64", x"64", x"64", x"62", x"61", x"64", x"65", x"65", x"64", x"67", 
        x"64", x"64", x"65", x"64", x"63", x"64", x"64", x"63", x"66", x"64", x"63", x"64", x"64", x"63", x"64", 
        x"64", x"62", x"61", x"63", x"65", x"65", x"63", x"63", x"65", x"65", x"65", x"65", x"66", x"67", x"65", 
        x"64", x"64", x"65", x"67", x"66", x"66", x"63", x"66", x"67", x"66", x"65", x"66", x"68", x"66", x"64", 
        x"65", x"69", x"67", x"66", x"69", x"65", x"6b", x"67", x"6c", x"69", x"5f", x"6d", x"95", x"bf", x"dc", 
        x"e1", x"be", x"8f", x"6d", x"5e", x"61", x"63", x"65", x"68", x"6c", x"6b", x"6a", x"6a", x"67", x"69", 
        x"69", x"65", x"65", x"66", x"69", x"66", x"67", x"68", x"67", x"67", x"66", x"65", x"68", x"68", x"66", 
        x"64", x"63", x"62", x"62", x"66", x"68", x"66", x"6a", x"69", x"67", x"69", x"67", x"66", x"68", x"68", 
        x"67", x"66", x"66", x"68", x"6a", x"68", x"68", x"68", x"69", x"69", x"65", x"68", x"6a", x"66", x"65", 
        x"69", x"67", x"65", x"6b", x"68", x"67", x"69", x"69", x"68", x"68", x"66", x"67", x"68", x"67", x"68", 
        x"69", x"67", x"67", x"68", x"68", x"68", x"68", x"68", x"6a", x"6a", x"6a", x"68", x"67", x"67", x"68", 
        x"67", x"67", x"6a", x"69", x"69", x"6a", x"6a", x"69", x"68", x"67", x"67", x"68", x"69", x"69", x"68", 
        x"66", x"69", x"68", x"68", x"6a", x"69", x"68", x"69", x"67", x"66", x"67", x"68", x"69", x"68", x"68", 
        x"66", x"66", x"68", x"68", x"66", x"68", x"6c", x"6c", x"6b", x"6c", x"6a", x"69", x"6a", x"6b", x"69", 
        x"68", x"69", x"69", x"67", x"65", x"65", x"67", x"65", x"69", x"6a", x"6b", x"68", x"68", x"67", x"6a", 
        x"69", x"67", x"69", x"68", x"68", x"6a", x"69", x"68", x"67", x"66", x"67", x"68", x"69", x"69", x"69", 
        x"69", x"69", x"67", x"67", x"68", x"69", x"67", x"66", x"67", x"66", x"67", x"65", x"66", x"68", x"6a", 
        x"69", x"67", x"67", x"67", x"65", x"68", x"67", x"66", x"67", x"65", x"64", x"66", x"67", x"6a", x"69", 
        x"6a", x"68", x"68", x"6c", x"6b", x"69", x"68", x"67", x"67", x"67", x"68", x"68", x"68", x"69", x"6b", 
        x"6c", x"69", x"67", x"67", x"67", x"66", x"64", x"65", x"69", x"69", x"65", x"68", x"6b", x"6a", x"6a", 
        x"6a", x"6b", x"6b", x"6b", x"68", x"67", x"68", x"66", x"66", x"68", x"67", x"65", x"64", x"67", x"6a", 
        x"6a", x"67", x"67", x"65", x"64", x"68", x"68", x"64", x"64", x"67", x"68", x"67", x"67", x"69", x"68", 
        x"69", x"66", x"66", x"65", x"65", x"66", x"66", x"66", x"66", x"66", x"65", x"67", x"67", x"65", x"68", 
        x"68", x"67", x"67", x"67", x"68", x"68", x"67", x"65", x"66", x"68", x"69", x"69", x"68", x"66", x"65", 
        x"65", x"64", x"67", x"67", x"65", x"64", x"65", x"66", x"66", x"69", x"68", x"65", x"64", x"63", x"62", 
        x"64", x"65", x"65", x"65", x"65", x"65", x"66", x"64", x"64", x"64", x"65", x"67", x"67", x"67", x"66", 
        x"65", x"67", x"68", x"68", x"67", x"67", x"67", x"67", x"66", x"65", x"63", x"63", x"63", x"63", x"62", 
        x"62", x"63", x"65", x"64", x"65", x"68", x"65", x"65", x"63", x"67", x"66", x"66", x"64", x"65", x"63", 
        x"62", x"65", x"64", x"62", x"65", x"66", x"64", x"65", x"66", x"62", x"63", x"64", x"64", x"63", x"62", 
        x"63", x"64", x"66", x"68", x"67", x"67", x"69", x"67", x"65", x"64", x"65", x"64", x"62", x"62", x"62", 
        x"63", x"63", x"62", x"62", x"64", x"65", x"65", x"65", x"64", x"64", x"64", x"64", x"63", x"62", x"62", 
        x"63", x"63", x"62", x"61", x"62", x"63", x"62", x"61", x"61", x"61", x"62", x"62", x"62", x"62", x"62", 
        x"63", x"63", x"64", x"64", x"63", x"62", x"61", x"61", x"61", x"61", x"63", x"63", x"62", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"62", x"62", x"61", 
        x"62", x"62", x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"62", x"62", x"63", 
        x"63", x"62", x"63", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"60", x"60", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5e", x"5e", x"5f", x"5f", x"5f", x"5e", x"5e", 
        x"5d", x"5d", x"5e", x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", x"5f", x"5f", 
        x"63", x"63", x"64", x"64", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"61", x"61", x"5f", x"61", x"62", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"63", x"62", x"61", x"61", x"61", x"60", x"60", x"62", 
        x"63", x"63", x"62", x"61", x"61", x"62", x"63", x"62", x"62", x"62", x"63", x"63", x"63", x"63", x"63", 
        x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"63", x"62", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"60", x"61", x"61", x"61", x"63", x"64", x"63", x"62", x"62", x"62", x"61", 
        x"62", x"62", x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"63", x"63", x"64", x"64", x"63", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"63", x"63", x"63", x"64", x"64", x"63", x"62", x"62", x"62", x"62", 
        x"62", x"61", x"63", x"64", x"65", x"64", x"63", x"64", x"64", x"64", x"64", x"63", x"63", x"63", x"63", 
        x"64", x"64", x"64", x"63", x"63", x"63", x"64", x"65", x"65", x"64", x"63", x"64", x"64", x"64", x"65", 
        x"65", x"65", x"66", x"65", x"63", x"63", x"64", x"63", x"65", x"64", x"64", x"66", x"64", x"62", x"63", 
        x"65", x"64", x"63", x"63", x"65", x"64", x"62", x"62", x"64", x"64", x"64", x"65", x"66", x"66", x"66", 
        x"66", x"64", x"65", x"67", x"65", x"66", x"64", x"63", x"64", x"64", x"65", x"67", x"69", x"69", x"66", 
        x"65", x"67", x"66", x"65", x"65", x"64", x"67", x"68", x"66", x"67", x"72", x"b0", x"ce", x"ab", x"a8", 
        x"c3", x"dc", x"e5", x"cf", x"9e", x"78", x"65", x"5a", x"63", x"6b", x"6c", x"6b", x"6b", x"69", x"69", 
        x"67", x"64", x"67", x"68", x"6b", x"6a", x"6a", x"6b", x"6a", x"69", x"67", x"66", x"65", x"65", x"65", 
        x"65", x"66", x"66", x"66", x"64", x"63", x"63", x"67", x"67", x"66", x"64", x"66", x"69", x"6a", x"6a", 
        x"69", x"68", x"69", x"6b", x"6b", x"6a", x"6b", x"68", x"67", x"69", x"6a", x"6c", x"6c", x"68", x"65", 
        x"68", x"68", x"68", x"6b", x"68", x"67", x"69", x"69", x"68", x"69", x"67", x"67", x"69", x"6b", x"6b", 
        x"69", x"69", x"68", x"67", x"66", x"67", x"68", x"6a", x"6a", x"6a", x"6b", x"6b", x"66", x"66", x"69", 
        x"68", x"66", x"69", x"69", x"6a", x"6b", x"6c", x"6b", x"69", x"67", x"67", x"68", x"69", x"6a", x"69", 
        x"68", x"6a", x"69", x"69", x"6a", x"6a", x"69", x"69", x"68", x"67", x"67", x"68", x"68", x"68", x"68", 
        x"68", x"68", x"69", x"68", x"66", x"67", x"6a", x"6a", x"69", x"6a", x"68", x"68", x"6a", x"6a", x"69", 
        x"6a", x"6a", x"69", x"68", x"67", x"67", x"67", x"69", x"6c", x"6b", x"6a", x"65", x"66", x"67", x"6a", 
        x"68", x"67", x"68", x"68", x"69", x"6c", x"6b", x"6a", x"69", x"67", x"67", x"66", x"65", x"67", x"69", 
        x"69", x"66", x"65", x"66", x"66", x"66", x"65", x"68", x"69", x"67", x"69", x"6b", x"6d", x"67", x"69", 
        x"69", x"68", x"68", x"68", x"67", x"66", x"64", x"63", x"66", x"67", x"67", x"6b", x"6a", x"6b", x"6b", 
        x"6a", x"67", x"67", x"6b", x"6a", x"6a", x"6a", x"6a", x"6a", x"69", x"68", x"69", x"69", x"67", x"69", 
        x"6b", x"6b", x"67", x"66", x"69", x"68", x"67", x"66", x"68", x"69", x"66", x"66", x"6b", x"67", x"69", 
        x"6a", x"68", x"6a", x"6b", x"68", x"66", x"68", x"69", x"69", x"6a", x"6a", x"67", x"65", x"66", x"68", 
        x"67", x"63", x"66", x"69", x"67", x"68", x"68", x"66", x"67", x"68", x"64", x"64", x"65", x"68", x"67", 
        x"68", x"65", x"66", x"67", x"67", x"66", x"65", x"65", x"65", x"64", x"65", x"68", x"68", x"65", x"67", 
        x"69", x"6b", x"6a", x"67", x"65", x"65", x"66", x"66", x"68", x"69", x"69", x"67", x"66", x"67", x"68", 
        x"66", x"65", x"66", x"66", x"64", x"64", x"66", x"66", x"66", x"69", x"68", x"66", x"65", x"66", x"65", 
        x"65", x"67", x"63", x"65", x"67", x"64", x"65", x"64", x"63", x"66", x"66", x"64", x"66", x"68", x"65", 
        x"65", x"68", x"69", x"68", x"67", x"66", x"66", x"65", x"64", x"63", x"64", x"65", x"65", x"64", x"65", 
        x"64", x"63", x"64", x"64", x"64", x"66", x"62", x"62", x"62", x"64", x"64", x"63", x"61", x"62", x"63", 
        x"63", x"63", x"63", x"63", x"63", x"65", x"66", x"66", x"66", x"63", x"64", x"64", x"62", x"63", x"63", 
        x"64", x"65", x"67", x"68", x"66", x"65", x"66", x"65", x"65", x"64", x"63", x"62", x"63", x"63", x"63", 
        x"64", x"64", x"65", x"65", x"63", x"64", x"65", x"66", x"65", x"64", x"63", x"63", x"64", x"63", x"64", 
        x"64", x"64", x"62", x"62", x"63", x"62", x"62", x"62", x"61", x"61", x"61", x"62", x"62", x"62", x"62", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"62", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"61", x"60", x"61", x"61", x"61", x"62", x"63", 
        x"64", x"62", x"61", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"60", x"60", x"60", x"60", x"5f", x"5f", x"60", x"5f", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", 
        x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", 
        x"5e", x"5e", x"5e", x"5f", x"5f", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", 
        x"63", x"64", x"65", x"64", x"62", x"62", x"63", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"62", 
        x"63", x"63", x"62", x"61", x"61", x"62", x"64", x"63", x"63", x"63", x"63", x"64", x"63", x"63", x"62", 
        x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"62", x"63", x"63", x"62", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"62", 
        x"62", x"61", x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"63", x"63", x"64", x"63", x"63", 
        x"62", x"62", x"62", x"63", x"63", x"64", x"64", x"64", x"64", x"64", x"64", x"62", x"62", x"62", x"63", 
        x"62", x"61", x"63", x"64", x"66", x"65", x"64", x"64", x"66", x"65", x"64", x"63", x"63", x"63", x"64", 
        x"65", x"64", x"63", x"63", x"63", x"63", x"64", x"65", x"66", x"67", x"62", x"63", x"65", x"64", x"63", 
        x"64", x"65", x"65", x"65", x"64", x"64", x"64", x"64", x"64", x"64", x"65", x"67", x"65", x"62", x"63", 
        x"65", x"66", x"66", x"66", x"65", x"65", x"65", x"64", x"64", x"64", x"65", x"66", x"65", x"65", x"66", 
        x"67", x"65", x"66", x"67", x"63", x"65", x"65", x"64", x"65", x"67", x"67", x"66", x"65", x"65", x"66", 
        x"67", x"6b", x"6b", x"6b", x"67", x"6b", x"6a", x"66", x"62", x"81", x"bd", x"c3", x"a4", x"9d", x"83", 
        x"72", x"94", x"bb", x"d7", x"e2", x"d2", x"ad", x"82", x"67", x"5e", x"61", x"69", x"6b", x"68", x"68", 
        x"66", x"65", x"6a", x"69", x"6a", x"6c", x"6c", x"6b", x"69", x"67", x"66", x"65", x"66", x"67", x"67", 
        x"66", x"66", x"66", x"66", x"64", x"65", x"67", x"69", x"68", x"67", x"66", x"66", x"66", x"69", x"69", 
        x"69", x"68", x"69", x"6b", x"6c", x"69", x"6a", x"6a", x"69", x"6c", x"6b", x"69", x"6c", x"69", x"65", 
        x"65", x"66", x"67", x"6b", x"68", x"67", x"6a", x"6a", x"69", x"69", x"68", x"66", x"68", x"6b", x"6b", 
        x"69", x"6a", x"69", x"68", x"68", x"69", x"6b", x"6b", x"69", x"68", x"6a", x"69", x"69", x"68", x"69", 
        x"69", x"68", x"67", x"67", x"67", x"69", x"6a", x"6a", x"69", x"6a", x"69", x"69", x"6a", x"6b", x"6b", 
        x"6a", x"6a", x"6a", x"6a", x"6b", x"6a", x"6a", x"6a", x"6a", x"6a", x"69", x"69", x"68", x"68", x"68", 
        x"69", x"6a", x"6a", x"68", x"66", x"66", x"68", x"66", x"65", x"68", x"68", x"68", x"6a", x"68", x"68", 
        x"6b", x"6a", x"69", x"69", x"69", x"68", x"66", x"65", x"69", x"6a", x"6a", x"66", x"68", x"6a", x"69", 
        x"68", x"69", x"6a", x"6a", x"69", x"68", x"69", x"6a", x"6a", x"6b", x"6a", x"69", x"68", x"69", x"6b", 
        x"6a", x"67", x"65", x"68", x"68", x"66", x"66", x"67", x"68", x"66", x"67", x"6a", x"6c", x"68", x"69", 
        x"69", x"69", x"69", x"6a", x"6a", x"6a", x"68", x"67", x"68", x"68", x"67", x"69", x"68", x"67", x"69", 
        x"67", x"65", x"66", x"69", x"6b", x"6b", x"6c", x"6c", x"6c", x"6b", x"6a", x"6a", x"6a", x"68", x"67", 
        x"68", x"69", x"68", x"68", x"6a", x"6c", x"6a", x"69", x"6a", x"69", x"67", x"66", x"68", x"65", x"66", 
        x"66", x"65", x"65", x"67", x"67", x"66", x"68", x"6a", x"6a", x"69", x"69", x"6a", x"6b", x"6a", x"6a", 
        x"68", x"66", x"6a", x"6c", x"69", x"68", x"67", x"67", x"6a", x"6b", x"69", x"69", x"6a", x"6c", x"6b", 
        x"6c", x"69", x"65", x"66", x"66", x"65", x"64", x"64", x"65", x"66", x"67", x"69", x"6a", x"69", x"69", 
        x"68", x"69", x"69", x"67", x"66", x"65", x"66", x"66", x"67", x"66", x"67", x"65", x"64", x"66", x"66", 
        x"65", x"66", x"67", x"66", x"65", x"65", x"66", x"66", x"65", x"68", x"67", x"65", x"65", x"65", x"66", 
        x"67", x"66", x"63", x"64", x"66", x"66", x"66", x"66", x"63", x"66", x"67", x"65", x"66", x"65", x"66", 
        x"67", x"67", x"67", x"68", x"67", x"65", x"65", x"66", x"64", x"64", x"66", x"68", x"68", x"66", x"64", 
        x"64", x"62", x"64", x"65", x"64", x"66", x"63", x"63", x"64", x"66", x"66", x"64", x"62", x"62", x"64", 
        x"64", x"63", x"63", x"64", x"63", x"64", x"65", x"66", x"66", x"65", x"64", x"63", x"64", x"64", x"64", 
        x"66", x"66", x"65", x"65", x"65", x"66", x"65", x"65", x"65", x"66", x"65", x"65", x"65", x"65", x"64", 
        x"64", x"64", x"65", x"65", x"64", x"63", x"64", x"65", x"65", x"64", x"64", x"63", x"63", x"64", x"64", 
        x"64", x"63", x"62", x"63", x"63", x"62", x"62", x"62", x"62", x"61", x"62", x"62", x"62", x"62", x"62", 
        x"63", x"63", x"63", x"63", x"63", x"64", x"63", x"63", x"62", x"61", x"62", x"63", x"63", x"63", x"63", 
        x"62", x"62", x"62", x"62", x"63", x"62", x"62", x"62", x"62", x"60", x"62", x"62", x"62", x"63", x"64", 
        x"62", x"61", x"62", x"63", x"63", x"62", x"61", x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"62", x"62", x"63", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"61", x"61", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", x"5e", 
        x"5f", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", 
        x"5e", x"5d", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5d", x"5c", 
        x"63", x"63", x"64", x"64", x"62", x"62", x"63", x"61", x"61", x"62", x"62", x"62", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"60", x"61", x"62", x"61", x"61", x"62", 
        x"62", x"62", x"61", x"61", x"61", x"61", x"60", x"60", x"61", x"62", x"61", x"61", x"61", x"61", x"62", 
        x"63", x"63", x"62", x"61", x"61", x"62", x"63", x"63", x"62", x"62", x"63", x"63", x"62", x"61", x"61", 
        x"62", x"62", x"62", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"62", x"61", x"62", x"62", x"62", x"62", x"63", x"61", x"61", x"61", x"62", 
        x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"62", x"63", x"64", x"62", x"61", x"63", x"65", x"65", 
        x"64", x"62", x"62", x"63", x"64", x"64", x"64", x"65", x"65", x"65", x"64", x"63", x"62", x"62", x"63", 
        x"63", x"62", x"63", x"64", x"65", x"65", x"63", x"63", x"65", x"67", x"66", x"65", x"64", x"64", x"64", 
        x"64", x"63", x"63", x"64", x"65", x"65", x"65", x"64", x"65", x"67", x"64", x"64", x"63", x"63", x"63", 
        x"66", x"64", x"64", x"64", x"65", x"65", x"65", x"66", x"66", x"64", x"64", x"65", x"63", x"63", x"65", 
        x"65", x"64", x"64", x"64", x"64", x"65", x"65", x"64", x"65", x"65", x"66", x"66", x"64", x"64", x"65", 
        x"69", x"67", x"67", x"66", x"62", x"64", x"65", x"65", x"66", x"67", x"67", x"66", x"66", x"68", x"68", 
        x"64", x"68", x"66", x"68", x"6a", x"68", x"61", x"68", x"90", x"c4", x"be", x"9c", x"a8", x"cd", x"9b", 
        x"60", x"5d", x"69", x"88", x"b3", x"db", x"ef", x"e3", x"b4", x"85", x"6a", x"5f", x"5f", x"67", x"6b", 
        x"69", x"64", x"65", x"66", x"68", x"6a", x"6a", x"68", x"67", x"67", x"67", x"67", x"67", x"67", x"67", 
        x"67", x"67", x"68", x"68", x"65", x"67", x"6c", x"6a", x"68", x"67", x"69", x"66", x"64", x"67", x"68", 
        x"67", x"64", x"64", x"68", x"69", x"64", x"66", x"69", x"6b", x"6c", x"6a", x"6c", x"6b", x"69", x"67", 
        x"67", x"68", x"67", x"6b", x"68", x"68", x"6a", x"6a", x"69", x"6a", x"68", x"67", x"68", x"6a", x"69", 
        x"68", x"69", x"6a", x"6b", x"6b", x"6c", x"6d", x"6c", x"69", x"68", x"67", x"67", x"6b", x"6c", x"69", 
        x"69", x"6c", x"6b", x"69", x"68", x"69", x"6b", x"6b", x"6b", x"6a", x"69", x"68", x"68", x"6a", x"6b", 
        x"6b", x"6a", x"6b", x"6b", x"6a", x"6a", x"6b", x"6a", x"6a", x"6a", x"69", x"68", x"68", x"68", x"69", 
        x"69", x"68", x"69", x"69", x"69", x"69", x"69", x"68", x"69", x"6b", x"6a", x"6a", x"6c", x"6b", x"6a", 
        x"6a", x"68", x"69", x"6a", x"6c", x"6b", x"69", x"66", x"6a", x"6b", x"6c", x"67", x"68", x"69", x"69", 
        x"6a", x"6a", x"6a", x"69", x"69", x"67", x"68", x"6a", x"6b", x"6b", x"6a", x"68", x"66", x"69", x"6d", 
        x"6c", x"69", x"69", x"6a", x"6a", x"69", x"68", x"69", x"6a", x"6c", x"6c", x"6c", x"6a", x"69", x"69", 
        x"6a", x"6b", x"6b", x"6c", x"6d", x"6a", x"69", x"69", x"69", x"6a", x"6a", x"6b", x"67", x"66", x"67", 
        x"66", x"66", x"69", x"6c", x"6d", x"6d", x"6e", x"6f", x"6e", x"6d", x"6b", x"6a", x"6a", x"6b", x"6a", 
        x"68", x"68", x"69", x"69", x"69", x"6c", x"6b", x"69", x"6a", x"69", x"68", x"6b", x"69", x"6a", x"69", 
        x"66", x"69", x"66", x"65", x"67", x"67", x"68", x"69", x"69", x"67", x"68", x"6a", x"6b", x"6a", x"67", 
        x"68", x"6b", x"6c", x"69", x"68", x"67", x"66", x"66", x"68", x"6a", x"6a", x"69", x"68", x"6a", x"69", 
        x"6a", x"67", x"65", x"67", x"68", x"67", x"66", x"67", x"68", x"67", x"68", x"69", x"6b", x"6f", x"6c", 
        x"69", x"65", x"65", x"67", x"69", x"68", x"67", x"66", x"65", x"65", x"68", x"67", x"65", x"67", x"67", 
        x"65", x"67", x"67", x"66", x"65", x"66", x"67", x"67", x"66", x"68", x"68", x"67", x"67", x"69", x"6a", 
        x"68", x"64", x"64", x"63", x"63", x"67", x"67", x"66", x"64", x"65", x"67", x"67", x"68", x"65", x"66", 
        x"68", x"65", x"65", x"67", x"69", x"66", x"66", x"67", x"65", x"65", x"65", x"66", x"66", x"65", x"68", 
        x"67", x"64", x"65", x"66", x"64", x"63", x"65", x"63", x"63", x"64", x"65", x"64", x"64", x"63", x"64", 
        x"65", x"65", x"65", x"65", x"63", x"64", x"65", x"64", x"65", x"66", x"65", x"64", x"63", x"64", x"64", 
        x"66", x"65", x"64", x"63", x"64", x"64", x"63", x"63", x"64", x"64", x"65", x"66", x"65", x"64", x"63", 
        x"63", x"63", x"63", x"64", x"64", x"63", x"63", x"63", x"63", x"65", x"66", x"63", x"62", x"63", x"64", 
        x"63", x"62", x"62", x"64", x"64", x"62", x"62", x"62", x"62", x"61", x"62", x"63", x"63", x"63", x"63", 
        x"64", x"63", x"63", x"62", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"62", x"63", x"64", x"63", 
        x"62", x"61", x"63", x"63", x"63", x"62", x"62", x"63", x"63", x"61", x"62", x"63", x"64", x"63", x"62", 
        x"60", x"61", x"64", x"64", x"64", x"64", x"62", x"61", x"61", x"62", x"62", x"62", x"62", x"62", x"61", 
        x"61", x"62", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"61", x"60", x"60", x"60", 
        x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5f", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", 
        x"5d", x"5d", x"5d", x"5e", x"5d", x"5d", x"5f", x"5f", x"5e", x"5d", x"5d", x"5e", x"5f", x"5d", x"5c", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"62", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"60", x"61", x"63", x"62", x"61", x"63", 
        x"63", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"61", x"62", x"62", x"62", 
        x"61", x"62", x"62", x"61", x"61", x"62", x"63", x"61", x"61", x"61", x"62", x"63", x"62", x"61", x"61", 
        x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"63", x"63", x"63", x"61", x"63", x"63", 
        x"62", x"61", x"62", x"63", x"64", x"62", x"61", x"62", x"63", x"63", x"63", x"61", x"61", x"61", x"61", 
        x"62", x"63", x"64", x"63", x"63", x"62", x"62", x"62", x"62", x"61", x"62", x"62", x"63", x"62", x"62", 
        x"63", x"64", x"64", x"63", x"63", x"63", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"63", x"63", 
        x"63", x"64", x"64", x"64", x"64", x"63", x"63", x"63", x"63", x"65", x"64", x"64", x"65", x"66", x"66", 
        x"65", x"64", x"64", x"64", x"65", x"64", x"64", x"63", x"64", x"65", x"67", x"65", x"62", x"63", x"64", 
        x"67", x"65", x"64", x"65", x"66", x"66", x"65", x"67", x"67", x"64", x"63", x"64", x"63", x"62", x"65", 
        x"64", x"64", x"63", x"64", x"64", x"64", x"64", x"64", x"65", x"65", x"66", x"66", x"65", x"65", x"64", 
        x"67", x"68", x"68", x"67", x"64", x"65", x"66", x"68", x"66", x"67", x"68", x"66", x"66", x"6a", x"6c", 
        x"64", x"68", x"69", x"69", x"63", x"5e", x"74", x"ae", x"c4", x"ac", x"9d", x"b7", x"ce", x"cb", x"99", 
        x"64", x"5e", x"5c", x"5f", x"68", x"80", x"a5", x"c8", x"e6", x"e2", x"c6", x"9d", x"74", x"5f", x"61", 
        x"65", x"67", x"69", x"66", x"66", x"66", x"66", x"67", x"67", x"68", x"68", x"69", x"69", x"68", x"67", 
        x"67", x"67", x"68", x"69", x"66", x"67", x"6b", x"68", x"67", x"69", x"69", x"69", x"69", x"6a", x"6b", 
        x"68", x"66", x"65", x"65", x"65", x"67", x"69", x"66", x"67", x"6a", x"6b", x"6d", x"67", x"66", x"68", 
        x"6a", x"6a", x"66", x"6b", x"69", x"68", x"6a", x"6a", x"69", x"6a", x"6a", x"6a", x"69", x"68", x"68", 
        x"68", x"68", x"69", x"6a", x"6a", x"6b", x"6a", x"6a", x"69", x"69", x"67", x"69", x"6c", x"6c", x"6a", 
        x"6b", x"6d", x"6b", x"69", x"69", x"69", x"6a", x"6a", x"6a", x"68", x"67", x"67", x"69", x"6a", x"6a", 
        x"69", x"69", x"6b", x"6b", x"69", x"6a", x"6b", x"6a", x"69", x"68", x"67", x"66", x"67", x"69", x"6a", 
        x"6a", x"69", x"6b", x"6c", x"6b", x"6a", x"68", x"69", x"6b", x"6c", x"6a", x"69", x"6b", x"6c", x"6a", 
        x"68", x"68", x"69", x"6a", x"6d", x"6c", x"6c", x"6d", x"6d", x"6a", x"69", x"66", x"68", x"6a", x"69", 
        x"6a", x"6a", x"67", x"68", x"69", x"68", x"69", x"68", x"68", x"68", x"68", x"68", x"68", x"6a", x"6a", 
        x"68", x"68", x"68", x"69", x"68", x"67", x"69", x"6a", x"6b", x"6e", x"6b", x"6a", x"67", x"68", x"67", 
        x"68", x"69", x"68", x"69", x"6b", x"6b", x"6d", x"6c", x"6a", x"69", x"69", x"66", x"68", x"68", x"6a", 
        x"69", x"6a", x"6c", x"6b", x"6e", x"6e", x"6f", x"70", x"70", x"6e", x"6d", x"6b", x"6b", x"6d", x"6c", 
        x"6a", x"6b", x"6a", x"69", x"69", x"6a", x"68", x"67", x"68", x"6a", x"69", x"6e", x"6c", x"6c", x"6e", 
        x"6c", x"6e", x"6b", x"68", x"69", x"69", x"67", x"68", x"69", x"68", x"6b", x"6d", x"6b", x"69", x"68", 
        x"69", x"6a", x"69", x"69", x"69", x"69", x"69", x"68", x"68", x"68", x"69", x"68", x"68", x"69", x"68", 
        x"69", x"65", x"65", x"68", x"6a", x"69", x"68", x"69", x"6b", x"66", x"66", x"65", x"68", x"6c", x"6a", 
        x"69", x"65", x"66", x"67", x"67", x"66", x"67", x"69", x"65", x"67", x"6c", x"69", x"67", x"69", x"69", 
        x"67", x"67", x"67", x"68", x"68", x"68", x"68", x"67", x"66", x"69", x"67", x"65", x"65", x"67", x"67", 
        x"66", x"64", x"65", x"64", x"63", x"66", x"67", x"66", x"66", x"66", x"68", x"68", x"67", x"66", x"66", 
        x"66", x"65", x"66", x"67", x"68", x"67", x"66", x"65", x"64", x"63", x"62", x"62", x"63", x"64", x"67", 
        x"68", x"66", x"67", x"68", x"66", x"64", x"67", x"64", x"63", x"62", x"65", x"65", x"66", x"66", x"63", 
        x"64", x"65", x"65", x"63", x"64", x"64", x"65", x"64", x"65", x"69", x"67", x"65", x"63", x"62", x"62", 
        x"63", x"64", x"64", x"64", x"64", x"65", x"65", x"65", x"64", x"62", x"64", x"67", x"64", x"63", x"63", 
        x"63", x"62", x"62", x"62", x"64", x"63", x"62", x"62", x"63", x"65", x"67", x"64", x"64", x"64", x"64", 
        x"62", x"62", x"63", x"64", x"65", x"63", x"63", x"62", x"62", x"61", x"62", x"63", x"63", x"63", x"63", 
        x"64", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"63", x"64", x"65", x"64", 
        x"62", x"61", x"63", x"63", x"63", x"62", x"62", x"63", x"64", x"62", x"61", x"62", x"63", x"62", x"61", 
        x"61", x"62", x"63", x"63", x"63", x"64", x"63", x"62", x"62", x"63", x"62", x"62", x"62", x"61", x"61", 
        x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"60", x"60", x"60", 
        x"60", x"61", x"61", x"60", x"60", x"60", x"60", x"5f", x"5d", x"5e", x"5f", x"5f", x"5f", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", 
        x"5d", x"5d", x"5d", x"5e", x"5d", x"5d", x"5f", x"5f", x"5e", x"5d", x"5d", x"5d", x"5e", x"5d", x"5c", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"60", x"61", x"63", x"62", x"61", x"64", 
        x"63", x"63", x"63", x"62", x"62", x"62", x"63", x"61", x"61", x"62", x"61", x"61", x"62", x"63", x"62", 
        x"60", x"61", x"62", x"62", x"61", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"62", x"62", x"62", 
        x"61", x"61", x"61", x"61", x"61", x"63", x"63", x"62", x"63", x"63", x"64", x"63", x"62", x"64", x"65", 
        x"62", x"61", x"62", x"64", x"65", x"62", x"61", x"62", x"63", x"63", x"63", x"61", x"61", x"61", x"61", 
        x"62", x"64", x"66", x"63", x"62", x"62", x"62", x"62", x"62", x"63", x"63", x"64", x"64", x"64", x"64", 
        x"63", x"63", x"63", x"62", x"63", x"63", x"63", x"64", x"63", x"64", x"64", x"65", x"64", x"63", x"62", 
        x"63", x"65", x"65", x"64", x"63", x"64", x"63", x"63", x"62", x"64", x"65", x"64", x"66", x"67", x"66", 
        x"65", x"65", x"65", x"64", x"64", x"63", x"63", x"63", x"64", x"66", x"66", x"64", x"62", x"66", x"65", 
        x"66", x"66", x"64", x"65", x"66", x"65", x"64", x"65", x"65", x"64", x"65", x"67", x"64", x"62", x"63", 
        x"64", x"67", x"68", x"66", x"62", x"63", x"65", x"65", x"64", x"65", x"66", x"67", x"67", x"66", x"64", 
        x"65", x"67", x"67", x"68", x"67", x"68", x"66", x"66", x"66", x"68", x"6a", x"68", x"67", x"6a", x"6a", 
        x"6b", x"6c", x"6a", x"65", x"62", x"80", x"b6", x"c3", x"a4", x"a2", x"c2", x"ce", x"cd", x"cb", x"9b", 
        x"63", x"60", x"5e", x"60", x"61", x"5c", x"68", x"78", x"9e", x"c3", x"dd", x"e3", x"ca", x"a5", x"80", 
        x"67", x"63", x"6a", x"6b", x"6b", x"66", x"67", x"68", x"69", x"69", x"68", x"68", x"6b", x"6b", x"69", 
        x"67", x"66", x"66", x"67", x"68", x"69", x"6b", x"67", x"69", x"6b", x"6a", x"68", x"69", x"6a", x"6a", 
        x"68", x"67", x"67", x"67", x"67", x"6a", x"6b", x"68", x"69", x"6b", x"69", x"6a", x"66", x"69", x"6b", 
        x"6b", x"6a", x"65", x"6b", x"69", x"68", x"6a", x"6a", x"69", x"6a", x"6c", x"6c", x"6a", x"67", x"67", 
        x"69", x"68", x"68", x"69", x"69", x"68", x"68", x"69", x"6b", x"6b", x"6a", x"6c", x"6a", x"69", x"6a", 
        x"6b", x"6c", x"6b", x"6b", x"6b", x"6c", x"6c", x"6a", x"69", x"67", x"67", x"69", x"6c", x"6d", x"6b", 
        x"69", x"69", x"6b", x"6b", x"69", x"6a", x"6b", x"6a", x"6a", x"6b", x"6a", x"68", x"68", x"6a", x"6c", 
        x"6a", x"6a", x"6c", x"6d", x"6c", x"6a", x"67", x"68", x"6d", x"6f", x"6d", x"6c", x"6d", x"6c", x"6a", 
        x"6a", x"6a", x"6a", x"6b", x"6a", x"69", x"6a", x"6c", x"6c", x"6a", x"69", x"68", x"6a", x"6a", x"68", 
        x"6a", x"6a", x"67", x"69", x"6b", x"6a", x"6b", x"6b", x"69", x"68", x"68", x"6a", x"6c", x"6c", x"68", 
        x"66", x"67", x"69", x"68", x"67", x"68", x"6b", x"6c", x"6c", x"6c", x"69", x"6c", x"6c", x"69", x"67", 
        x"68", x"69", x"68", x"68", x"6a", x"68", x"6b", x"6b", x"69", x"6a", x"6b", x"66", x"67", x"67", x"6a", 
        x"6a", x"6d", x"6e", x"6a", x"6d", x"6f", x"70", x"71", x"71", x"6f", x"6e", x"6d", x"6d", x"6e", x"6b", 
        x"69", x"6b", x"6c", x"6b", x"6b", x"6b", x"67", x"66", x"6a", x"6d", x"6c", x"6a", x"6b", x"68", x"6c", 
        x"6d", x"6c", x"6c", x"6a", x"6c", x"6a", x"67", x"67", x"69", x"6a", x"6b", x"6a", x"69", x"6a", x"6c", 
        x"6b", x"66", x"66", x"69", x"6a", x"69", x"69", x"69", x"69", x"67", x"68", x"68", x"69", x"6b", x"69", 
        x"68", x"65", x"65", x"68", x"6a", x"69", x"67", x"68", x"6a", x"67", x"69", x"67", x"67", x"68", x"67", 
        x"6a", x"66", x"66", x"67", x"67", x"66", x"66", x"68", x"65", x"67", x"6d", x"69", x"67", x"68", x"69", 
        x"68", x"67", x"68", x"69", x"69", x"68", x"67", x"67", x"66", x"68", x"67", x"65", x"65", x"67", x"67", 
        x"63", x"66", x"66", x"66", x"66", x"64", x"66", x"67", x"6a", x"69", x"68", x"66", x"63", x"66", x"66", 
        x"66", x"69", x"68", x"67", x"66", x"66", x"65", x"62", x"63", x"63", x"63", x"63", x"65", x"66", x"66", 
        x"67", x"66", x"68", x"6a", x"67", x"64", x"65", x"63", x"65", x"64", x"67", x"65", x"65", x"67", x"63", 
        x"63", x"65", x"64", x"62", x"64", x"64", x"66", x"65", x"66", x"6b", x"69", x"67", x"64", x"62", x"62", 
        x"62", x"63", x"64", x"64", x"64", x"66", x"67", x"68", x"66", x"62", x"62", x"65", x"64", x"64", x"64", 
        x"65", x"65", x"64", x"64", x"64", x"63", x"62", x"62", x"64", x"66", x"67", x"65", x"65", x"65", x"64", 
        x"63", x"63", x"65", x"65", x"65", x"65", x"63", x"63", x"62", x"61", x"62", x"63", x"63", x"63", x"63", 
        x"64", x"64", x"63", x"62", x"61", x"61", x"61", x"62", x"63", x"63", x"62", x"63", x"64", x"64", x"63", 
        x"63", x"61", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"61", x"61", x"62", x"62", x"61", 
        x"62", x"63", x"63", x"62", x"62", x"64", x"64", x"62", x"62", x"63", x"63", x"62", x"62", x"61", x"61", 
        x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"5f", x"60", x"60", x"60", x"5f", x"5e", x"5d", 
        x"5d", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", x"5d", x"5e", x"5e", x"5d", x"5d", x"5d", x"5f", x"5f", 
        x"5e", x"5e", x"5e", x"5f", x"5f", x"5e", x"5e", x"5f", x"5f", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", 
        x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"62", 
        x"60", x"62", x"63", x"60", x"61", x"62", x"61", x"62", x"61", x"60", x"60", x"61", x"62", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"62", x"61", x"61", x"62", x"64", x"63", 
        x"61", x"61", x"62", x"63", x"63", x"61", x"61", x"62", x"63", x"63", x"62", x"61", x"62", x"63", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"63", x"63", x"63", x"64", x"64", x"64", x"63", x"61", x"62", x"63", 
        x"63", x"62", x"63", x"63", x"62", x"62", x"62", x"62", x"63", x"63", x"63", x"63", x"62", x"61", x"61", 
        x"62", x"63", x"63", x"64", x"64", x"64", x"66", x"65", x"64", x"66", x"66", x"63", x"63", x"65", x"64", 
        x"64", x"64", x"61", x"62", x"62", x"63", x"64", x"64", x"65", x"64", x"62", x"63", x"62", x"62", x"62", 
        x"60", x"65", x"64", x"65", x"65", x"63", x"63", x"65", x"65", x"64", x"67", x"65", x"64", x"65", x"65", 
        x"64", x"65", x"65", x"62", x"65", x"64", x"63", x"63", x"63", x"66", x"66", x"65", x"62", x"63", x"63", 
        x"65", x"65", x"67", x"67", x"65", x"64", x"64", x"63", x"63", x"65", x"67", x"66", x"63", x"62", x"63", 
        x"62", x"67", x"67", x"65", x"61", x"63", x"67", x"66", x"64", x"66", x"66", x"68", x"66", x"65", x"64", 
        x"67", x"66", x"67", x"68", x"68", x"67", x"65", x"66", x"66", x"6b", x"6b", x"6a", x"68", x"69", x"68", 
        x"69", x"6a", x"63", x"5f", x"95", x"cb", x"c0", x"94", x"b3", x"cc", x"d1", x"cf", x"cd", x"cb", x"a1", 
        x"65", x"5e", x"5d", x"5f", x"61", x"5e", x"5c", x"5a", x"60", x"6d", x"89", x"b9", x"de", x"eb", x"de", 
        x"bc", x"8e", x"66", x"5b", x"66", x"70", x"6e", x"69", x"67", x"6b", x"68", x"6a", x"69", x"69", x"68", 
        x"66", x"69", x"6a", x"6b", x"6b", x"69", x"68", x"6a", x"6b", x"68", x"68", x"68", x"66", x"68", x"69", 
        x"6a", x"69", x"68", x"69", x"6a", x"6a", x"6b", x"6b", x"6b", x"6a", x"67", x"68", x"6a", x"6b", x"69", 
        x"68", x"6c", x"69", x"6a", x"6a", x"6a", x"6b", x"6b", x"69", x"69", x"6a", x"6a", x"6a", x"6a", x"69", 
        x"69", x"6b", x"6b", x"68", x"69", x"6b", x"6c", x"6a", x"6a", x"6b", x"6a", x"69", x"6a", x"6a", x"6a", 
        x"6b", x"6b", x"67", x"6a", x"6b", x"6c", x"6b", x"68", x"68", x"68", x"67", x"69", x"6b", x"6b", x"69", 
        x"6a", x"6a", x"67", x"68", x"6b", x"6f", x"6d", x"69", x"68", x"6a", x"6a", x"6a", x"6a", x"6a", x"69", 
        x"68", x"6b", x"6d", x"6b", x"6a", x"6b", x"6b", x"6b", x"6d", x"6c", x"6b", x"6b", x"6e", x"6e", x"6e", 
        x"6e", x"6c", x"6b", x"6a", x"67", x"66", x"67", x"69", x"69", x"68", x"68", x"6b", x"6b", x"67", x"68", 
        x"6b", x"6a", x"69", x"6c", x"6f", x"6f", x"6f", x"6b", x"69", x"6a", x"69", x"69", x"68", x"67", x"67", 
        x"68", x"68", x"67", x"69", x"6a", x"68", x"69", x"69", x"69", x"6c", x"6a", x"6c", x"6d", x"69", x"6c", 
        x"6c", x"6a", x"69", x"68", x"68", x"68", x"69", x"6a", x"6b", x"6a", x"69", x"67", x"68", x"68", x"69", 
        x"69", x"6a", x"6c", x"6d", x"6e", x"6e", x"70", x"71", x"71", x"71", x"70", x"6e", x"6e", x"6f", x"6b", 
        x"69", x"67", x"67", x"6a", x"69", x"6c", x"6a", x"67", x"69", x"6b", x"69", x"6a", x"6c", x"66", x"66", 
        x"68", x"66", x"68", x"66", x"68", x"65", x"66", x"67", x"68", x"67", x"68", x"68", x"6a", x"6a", x"6b", 
        x"68", x"65", x"66", x"68", x"67", x"6a", x"6b", x"67", x"66", x"65", x"64", x"67", x"69", x"6a", x"68", 
        x"69", x"68", x"65", x"67", x"68", x"67", x"66", x"66", x"67", x"69", x"68", x"67", x"67", x"68", x"68", 
        x"69", x"66", x"66", x"63", x"66", x"68", x"65", x"66", x"65", x"63", x"67", x"65", x"67", x"66", x"68", 
        x"69", x"66", x"66", x"68", x"69", x"67", x"66", x"66", x"67", x"68", x"68", x"68", x"66", x"68", x"68", 
        x"64", x"68", x"68", x"69", x"68", x"67", x"67", x"69", x"69", x"66", x"67", x"65", x"65", x"63", x"66", 
        x"67", x"68", x"68", x"66", x"67", x"66", x"66", x"64", x"65", x"64", x"64", x"64", x"65", x"67", x"68", 
        x"69", x"6a", x"69", x"67", x"67", x"65", x"65", x"65", x"66", x"65", x"66", x"64", x"64", x"69", x"65", 
        x"64", x"64", x"64", x"63", x"65", x"64", x"67", x"65", x"65", x"67", x"67", x"67", x"64", x"65", x"65", 
        x"66", x"65", x"64", x"64", x"63", x"64", x"64", x"64", x"66", x"63", x"63", x"68", x"63", x"62", x"64", 
        x"63", x"63", x"65", x"63", x"63", x"64", x"63", x"63", x"65", x"68", x"66", x"65", x"64", x"64", x"65", 
        x"66", x"65", x"64", x"64", x"65", x"65", x"64", x"63", x"64", x"64", x"63", x"63", x"63", x"63", x"66", 
        x"68", x"66", x"62", x"63", x"64", x"65", x"65", x"65", x"64", x"63", x"62", x"62", x"62", x"63", x"63", 
        x"62", x"62", x"65", x"62", x"61", x"62", x"63", x"64", x"64", x"63", x"62", x"63", x"65", x"62", x"63", 
        x"62", x"62", x"63", x"63", x"61", x"62", x"63", x"63", x"62", x"63", x"63", x"62", x"62", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"62", x"62", x"61", x"63", x"63", x"62", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"5e", x"5e", x"60", x"61", x"60", x"5f", x"5f", x"5f", x"5f", x"5f", x"60", x"61", x"61", 
        x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", 
        x"61", x"63", x"64", x"61", x"62", x"63", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"65", x"63", 
        x"61", x"61", x"62", x"64", x"63", x"61", x"61", x"63", x"64", x"64", x"63", x"62", x"62", x"63", x"63", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"61", x"61", 
        x"62", x"63", x"63", x"63", x"62", x"62", x"62", x"63", x"63", x"63", x"63", x"64", x"63", x"63", x"62", 
        x"63", x"63", x"62", x"64", x"63", x"62", x"64", x"64", x"62", x"63", x"66", x"63", x"62", x"64", x"62", 
        x"63", x"65", x"64", x"64", x"65", x"65", x"64", x"63", x"63", x"62", x"61", x"62", x"62", x"65", x"64", 
        x"62", x"65", x"65", x"64", x"65", x"65", x"66", x"68", x"6a", x"65", x"67", x"66", x"65", x"65", x"66", 
        x"68", x"66", x"63", x"64", x"69", x"66", x"64", x"65", x"64", x"63", x"65", x"64", x"62", x"61", x"63", 
        x"65", x"63", x"66", x"65", x"64", x"66", x"68", x"67", x"64", x"64", x"64", x"64", x"63", x"62", x"63", 
        x"65", x"6a", x"66", x"65", x"65", x"67", x"68", x"66", x"64", x"66", x"65", x"69", x"67", x"67", x"67", 
        x"69", x"68", x"68", x"67", x"65", x"65", x"67", x"6b", x"69", x"65", x"69", x"6b", x"67", x"6a", x"66", 
        x"64", x"61", x"76", x"af", x"cf", x"a8", x"7b", x"af", x"d4", x"d0", x"ce", x"cc", x"ce", x"ca", x"a4", 
        x"66", x"5d", x"5e", x"5f", x"5f", x"60", x"5f", x"5e", x"5e", x"5c", x"5d", x"67", x"7e", x"a4", x"cd", 
        x"e2", x"e1", x"ca", x"9e", x"77", x"64", x"60", x"67", x"69", x"6b", x"6a", x"6a", x"65", x"6d", x"6e", 
        x"67", x"6a", x"6c", x"68", x"66", x"69", x"6a", x"6c", x"6b", x"67", x"6b", x"6a", x"68", x"69", x"6a", 
        x"6a", x"69", x"68", x"69", x"6b", x"69", x"68", x"68", x"69", x"6a", x"69", x"68", x"6a", x"6c", x"69", 
        x"67", x"6d", x"6c", x"6c", x"6c", x"6c", x"6c", x"6a", x"68", x"66", x"69", x"69", x"6b", x"6b", x"6a", 
        x"6a", x"6c", x"6a", x"68", x"68", x"6a", x"6c", x"6a", x"69", x"68", x"68", x"69", x"68", x"68", x"6b", 
        x"6c", x"69", x"67", x"69", x"6a", x"6b", x"6b", x"69", x"6b", x"6b", x"6a", x"6b", x"6c", x"6a", x"69", 
        x"6c", x"6e", x"69", x"67", x"68", x"6a", x"6a", x"6b", x"69", x"69", x"6a", x"6a", x"69", x"67", x"65", 
        x"69", x"6c", x"6c", x"6b", x"6a", x"6a", x"6b", x"6d", x"6c", x"6b", x"6b", x"6c", x"6c", x"6c", x"6a", 
        x"69", x"69", x"6a", x"6a", x"68", x"67", x"68", x"6a", x"6b", x"69", x"67", x"69", x"6a", x"68", x"6b", 
        x"6c", x"6a", x"68", x"6a", x"6b", x"69", x"6b", x"69", x"69", x"6c", x"6b", x"69", x"68", x"68", x"6a", 
        x"6c", x"6b", x"69", x"6d", x"6e", x"6b", x"6c", x"6c", x"6a", x"6a", x"6a", x"6a", x"6b", x"6a", x"6d", 
        x"6f", x"6d", x"6c", x"6c", x"6a", x"69", x"6a", x"6c", x"6c", x"68", x"65", x"69", x"6b", x"6b", x"6a", 
        x"69", x"69", x"6b", x"6d", x"6e", x"6f", x"70", x"71", x"71", x"71", x"70", x"6f", x"71", x"71", x"6c", 
        x"6a", x"67", x"68", x"6b", x"69", x"6d", x"6b", x"68", x"69", x"6b", x"68", x"6a", x"6c", x"69", x"68", 
        x"6b", x"69", x"6a", x"66", x"67", x"65", x"67", x"68", x"67", x"67", x"67", x"66", x"66", x"66", x"66", 
        x"67", x"69", x"6a", x"68", x"66", x"6a", x"6d", x"6a", x"68", x"67", x"65", x"67", x"68", x"68", x"65", 
        x"67", x"67", x"67", x"68", x"68", x"67", x"67", x"67", x"68", x"69", x"67", x"67", x"67", x"69", x"6a", 
        x"69", x"69", x"6d", x"6b", x"6c", x"69", x"64", x"69", x"6a", x"65", x"68", x"65", x"68", x"65", x"66", 
        x"68", x"69", x"67", x"68", x"69", x"66", x"65", x"65", x"66", x"67", x"67", x"67", x"65", x"67", x"66", 
        x"67", x"6a", x"68", x"68", x"67", x"6a", x"6a", x"69", x"69", x"66", x"69", x"66", x"66", x"63", x"66", 
        x"67", x"69", x"68", x"68", x"68", x"66", x"67", x"67", x"66", x"65", x"64", x"64", x"64", x"65", x"64", 
        x"65", x"68", x"66", x"65", x"67", x"65", x"67", x"68", x"68", x"68", x"68", x"67", x"67", x"6b", x"67", 
        x"66", x"65", x"66", x"65", x"66", x"65", x"67", x"66", x"64", x"64", x"67", x"66", x"63", x"64", x"64", 
        x"65", x"66", x"64", x"64", x"63", x"67", x"65", x"62", x"66", x"67", x"65", x"65", x"63", x"63", x"64", 
        x"62", x"62", x"65", x"62", x"62", x"64", x"64", x"65", x"66", x"67", x"65", x"63", x"63", x"63", x"63", 
        x"64", x"63", x"62", x"64", x"67", x"67", x"65", x"65", x"66", x"66", x"65", x"65", x"65", x"65", x"66", 
        x"67", x"65", x"62", x"64", x"64", x"65", x"64", x"65", x"64", x"64", x"62", x"62", x"62", x"62", x"62", 
        x"62", x"62", x"64", x"61", x"61", x"62", x"63", x"66", x"65", x"64", x"62", x"63", x"65", x"62", x"63", 
        x"62", x"61", x"63", x"64", x"61", x"61", x"64", x"63", x"62", x"64", x"64", x"63", x"62", x"62", x"62", 
        x"62", x"62", x"63", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"62", x"62", x"62", x"63", x"64", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"60", x"60", x"5f", x"5f", x"60", x"61", x"61", x"61", 
        x"62", x"61", x"61", x"60", x"60", x"60", x"60", x"61", x"60", x"60", x"60", x"60", x"61", x"60", x"60", 
        x"63", x"63", x"63", x"63", x"64", x"64", x"63", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", 
        x"62", x"63", x"64", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"64", x"63", 
        x"62", x"62", x"63", x"64", x"63", x"61", x"61", x"62", x"63", x"64", x"63", x"63", x"62", x"63", x"63", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"61", x"61", x"61", x"61", x"61", 
        x"62", x"63", x"64", x"63", x"62", x"62", x"62", x"62", x"63", x"64", x"64", x"64", x"64", x"64", x"63", 
        x"62", x"62", x"63", x"64", x"63", x"61", x"62", x"63", x"61", x"61", x"66", x"65", x"61", x"64", x"62", 
        x"62", x"66", x"66", x"64", x"64", x"64", x"64", x"63", x"63", x"62", x"62", x"62", x"61", x"63", x"63", 
        x"61", x"62", x"66", x"63", x"63", x"65", x"65", x"63", x"65", x"66", x"6b", x"6c", x"69", x"65", x"65", 
        x"67", x"64", x"61", x"65", x"68", x"64", x"63", x"65", x"65", x"63", x"66", x"67", x"66", x"66", x"67", 
        x"68", x"67", x"68", x"66", x"63", x"65", x"67", x"68", x"67", x"66", x"65", x"66", x"68", x"67", x"64", 
        x"67", x"6a", x"65", x"64", x"65", x"67", x"67", x"68", x"69", x"68", x"65", x"68", x"66", x"67", x"69", 
        x"6a", x"65", x"64", x"68", x"68", x"65", x"65", x"68", x"67", x"64", x"68", x"6c", x"68", x"68", x"61", 
        x"64", x"81", x"c2", x"cc", x"93", x"84", x"b3", x"cd", x"cc", x"c9", x"cf", x"ce", x"ce", x"c9", x"a4", 
        x"66", x"5d", x"5e", x"5f", x"5f", x"5c", x"5b", x"5b", x"5d", x"60", x"62", x"5f", x"5b", x"62", x"77", 
        x"9e", x"c8", x"e6", x"e9", x"d8", x"a9", x"75", x"62", x"62", x"67", x"67", x"68", x"6a", x"68", x"68", 
        x"68", x"68", x"66", x"67", x"66", x"6a", x"6c", x"6c", x"6b", x"69", x"6b", x"6b", x"6a", x"6a", x"6a", 
        x"69", x"69", x"68", x"69", x"6b", x"69", x"68", x"68", x"6a", x"6b", x"6b", x"68", x"69", x"6d", x"6c", 
        x"69", x"6d", x"6c", x"6b", x"6c", x"6c", x"6c", x"6b", x"6a", x"69", x"69", x"6a", x"6a", x"6a", x"6b", 
        x"6c", x"6c", x"6b", x"6b", x"6a", x"6a", x"6b", x"6c", x"6c", x"6b", x"6c", x"6c", x"68", x"67", x"68", 
        x"67", x"65", x"67", x"6a", x"69", x"6b", x"6b", x"6a", x"6d", x"6d", x"6c", x"6c", x"6c", x"6c", x"6a", 
        x"6c", x"6e", x"6b", x"68", x"66", x"65", x"68", x"6d", x"69", x"68", x"69", x"69", x"69", x"69", x"69", 
        x"6c", x"6d", x"6c", x"6c", x"6a", x"68", x"69", x"6b", x"6a", x"6a", x"6b", x"6d", x"6d", x"6e", x"6a", 
        x"67", x"69", x"6b", x"6c", x"6c", x"6b", x"69", x"69", x"6c", x"6b", x"68", x"67", x"69", x"69", x"6b", 
        x"6b", x"69", x"68", x"6a", x"6b", x"68", x"69", x"6a", x"6b", x"6b", x"6a", x"6b", x"6a", x"6a", x"6c", 
        x"6d", x"6c", x"6a", x"6c", x"6d", x"6a", x"6b", x"6d", x"6a", x"67", x"69", x"6c", x"6b", x"68", x"6b", 
        x"6c", x"6b", x"6b", x"6b", x"6b", x"6a", x"6a", x"6c", x"6b", x"67", x"66", x"69", x"6e", x"6f", x"6c", 
        x"6b", x"6a", x"6a", x"6a", x"6c", x"6f", x"70", x"70", x"70", x"71", x"71", x"71", x"72", x"71", x"6d", 
        x"6c", x"6b", x"6b", x"6d", x"6b", x"6e", x"6c", x"69", x"6a", x"6c", x"6a", x"6a", x"6d", x"6b", x"69", 
        x"6b", x"6a", x"69", x"68", x"68", x"68", x"69", x"68", x"68", x"67", x"68", x"68", x"69", x"69", x"6a", 
        x"6b", x"6b", x"6b", x"69", x"67", x"68", x"69", x"68", x"65", x"65", x"69", x"6a", x"69", x"68", x"66", 
        x"67", x"67", x"6a", x"69", x"68", x"68", x"69", x"69", x"69", x"69", x"68", x"67", x"68", x"69", x"69", 
        x"69", x"66", x"6a", x"6c", x"6b", x"67", x"64", x"69", x"6b", x"67", x"6a", x"66", x"67", x"65", x"66", 
        x"66", x"69", x"67", x"69", x"69", x"67", x"66", x"66", x"65", x"65", x"65", x"65", x"64", x"66", x"67", 
        x"67", x"6a", x"69", x"68", x"68", x"6b", x"6b", x"68", x"69", x"68", x"67", x"65", x"65", x"64", x"67", 
        x"67", x"6a", x"68", x"68", x"69", x"67", x"68", x"69", x"66", x"65", x"65", x"66", x"65", x"64", x"65", 
        x"64", x"66", x"64", x"64", x"65", x"63", x"67", x"68", x"69", x"69", x"68", x"67", x"66", x"67", x"66", 
        x"66", x"66", x"69", x"6a", x"6a", x"67", x"69", x"67", x"67", x"67", x"68", x"69", x"65", x"65", x"64", 
        x"66", x"67", x"65", x"63", x"63", x"68", x"69", x"64", x"66", x"68", x"64", x"62", x"64", x"64", x"65", 
        x"63", x"63", x"65", x"62", x"62", x"64", x"66", x"66", x"65", x"65", x"63", x"64", x"64", x"65", x"65", 
        x"65", x"64", x"64", x"65", x"65", x"65", x"66", x"67", x"67", x"68", x"66", x"63", x"63", x"66", x"67", 
        x"67", x"66", x"65", x"65", x"64", x"62", x"62", x"63", x"64", x"64", x"61", x"61", x"61", x"61", x"62", 
        x"63", x"64", x"63", x"61", x"62", x"63", x"64", x"66", x"65", x"64", x"63", x"63", x"64", x"63", x"64", 
        x"63", x"62", x"64", x"64", x"61", x"61", x"64", x"64", x"63", x"64", x"64", x"64", x"63", x"63", x"62", 
        x"62", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"61", x"62", x"63", x"62", x"62", x"63", x"62", x"61", x"61", x"61", x"60", x"60", x"61", x"61", x"60", 
        x"60", x"60", x"61", x"61", x"61", x"60", x"60", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"61", 
        x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", 
        x"64", x"63", x"63", x"64", x"64", x"64", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"63", x"64", x"63", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"61", x"61", x"61", x"61", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"63", x"63", 
        x"63", x"64", x"64", x"64", x"62", x"61", x"61", x"62", x"63", x"64", x"64", x"63", x"63", x"63", x"63", 
        x"63", x"63", x"63", x"63", x"62", x"62", x"62", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"62", 
        x"62", x"63", x"64", x"63", x"63", x"62", x"62", x"62", x"63", x"64", x"65", x"63", x"64", x"65", x"64", 
        x"62", x"62", x"63", x"66", x"66", x"64", x"64", x"65", x"64", x"63", x"67", x"67", x"62", x"66", x"65", 
        x"63", x"65", x"65", x"63", x"64", x"64", x"64", x"64", x"64", x"64", x"67", x"65", x"62", x"61", x"62", 
        x"62", x"63", x"63", x"61", x"62", x"65", x"65", x"65", x"64", x"65", x"68", x"6a", x"69", x"66", x"66", 
        x"68", x"65", x"62", x"64", x"64", x"63", x"63", x"64", x"63", x"61", x"63", x"64", x"64", x"64", x"64", 
        x"65", x"66", x"67", x"65", x"64", x"65", x"6a", x"69", x"67", x"67", x"67", x"67", x"68", x"68", x"65", 
        x"66", x"69", x"67", x"64", x"65", x"67", x"67", x"67", x"66", x"66", x"65", x"69", x"68", x"6a", x"6b", 
        x"6a", x"65", x"64", x"67", x"68", x"68", x"67", x"68", x"68", x"6b", x"66", x"68", x"6b", x"65", x"69", 
        x"92", x"c8", x"be", x"8b", x"94", x"bd", x"cd", x"c4", x"cc", x"cf", x"d1", x"cb", x"ce", x"cc", x"a5", 
        x"67", x"5d", x"5e", x"5f", x"5f", x"5f", x"60", x"61", x"5d", x"5e", x"62", x"63", x"61", x"60", x"5f", 
        x"64", x"73", x"94", x"c1", x"e0", x"e8", x"db", x"b4", x"87", x"67", x"61", x"6c", x"6c", x"6d", x"6b", 
        x"68", x"68", x"6b", x"69", x"6a", x"6d", x"6b", x"6b", x"6d", x"6b", x"68", x"6a", x"6c", x"6b", x"69", 
        x"69", x"69", x"6a", x"6a", x"69", x"69", x"69", x"6a", x"6b", x"6a", x"6a", x"69", x"69", x"6d", x"6d", 
        x"6a", x"6b", x"6b", x"6d", x"6d", x"6d", x"6c", x"6b", x"69", x"67", x"69", x"6b", x"6b", x"6a", x"6c", 
        x"6e", x"6b", x"6c", x"6e", x"6d", x"6b", x"6d", x"70", x"6f", x"6d", x"6b", x"69", x"6a", x"6a", x"68", 
        x"69", x"6a", x"6a", x"6c", x"6b", x"6c", x"6c", x"6b", x"6e", x"6d", x"6c", x"6c", x"6b", x"6b", x"6a", 
        x"6a", x"6b", x"69", x"69", x"69", x"67", x"6a", x"6f", x"6d", x"6b", x"6b", x"6a", x"6a", x"69", x"69", 
        x"69", x"6a", x"69", x"6a", x"6b", x"6b", x"6e", x"6d", x"6a", x"69", x"68", x"68", x"69", x"69", x"69", 
        x"6a", x"6e", x"6e", x"6e", x"6e", x"6d", x"6b", x"6a", x"6b", x"6c", x"6c", x"6b", x"6a", x"68", x"6a", 
        x"6b", x"6a", x"6b", x"6c", x"6d", x"6c", x"6b", x"6c", x"6c", x"6a", x"69", x"6b", x"6b", x"6c", x"6c", 
        x"6c", x"6c", x"6b", x"6c", x"6c", x"69", x"6b", x"6c", x"6c", x"67", x"68", x"6c", x"6c", x"6b", x"6c", 
        x"6c", x"6b", x"6a", x"6b", x"6b", x"6a", x"68", x"68", x"69", x"6a", x"6a", x"69", x"6b", x"6a", x"6a", 
        x"6a", x"6c", x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"71", x"72", x"71", x"71", x"70", x"70", 
        x"70", x"6e", x"6d", x"6d", x"6c", x"6d", x"6c", x"6a", x"6b", x"6c", x"6a", x"69", x"6b", x"69", x"67", 
        x"69", x"69", x"67", x"6b", x"6a", x"6c", x"6c", x"6a", x"6c", x"6b", x"6c", x"6c", x"6b", x"6c", x"6c", 
        x"6a", x"69", x"6a", x"6b", x"6a", x"69", x"6b", x"6d", x"6b", x"69", x"6c", x"6b", x"69", x"69", x"68", 
        x"68", x"68", x"6b", x"69", x"69", x"6a", x"6a", x"6a", x"69", x"6a", x"68", x"68", x"68", x"6a", x"6a", 
        x"69", x"68", x"69", x"69", x"6a", x"69", x"68", x"6a", x"68", x"66", x"6a", x"65", x"67", x"67", x"67", 
        x"67", x"68", x"67", x"69", x"6a", x"67", x"66", x"67", x"66", x"67", x"66", x"67", x"67", x"6a", x"6b", 
        x"66", x"69", x"6a", x"69", x"69", x"6a", x"6a", x"6b", x"6c", x"6a", x"68", x"68", x"69", x"68", x"69", 
        x"68", x"6a", x"68", x"68", x"69", x"68", x"69", x"68", x"65", x"64", x"66", x"67", x"65", x"66", x"69", 
        x"66", x"67", x"66", x"66", x"67", x"64", x"64", x"66", x"67", x"68", x"68", x"67", x"67", x"66", x"66", 
        x"67", x"66", x"6a", x"6c", x"6a", x"69", x"6a", x"69", x"6a", x"6a", x"6a", x"6b", x"69", x"68", x"66", 
        x"67", x"69", x"69", x"66", x"63", x"68", x"6b", x"66", x"65", x"64", x"63", x"64", x"66", x"65", x"66", 
        x"64", x"64", x"64", x"63", x"63", x"66", x"66", x"65", x"63", x"64", x"64", x"64", x"64", x"66", x"65", 
        x"64", x"64", x"65", x"65", x"63", x"63", x"66", x"66", x"66", x"67", x"67", x"64", x"64", x"66", x"66", 
        x"63", x"63", x"65", x"65", x"64", x"63", x"63", x"64", x"65", x"65", x"64", x"63", x"62", x"61", x"61", 
        x"61", x"61", x"63", x"62", x"64", x"64", x"64", x"65", x"64", x"64", x"64", x"63", x"63", x"65", x"66", 
        x"64", x"63", x"64", x"64", x"61", x"61", x"64", x"65", x"64", x"65", x"65", x"65", x"65", x"64", x"63", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"61", x"61", x"61", 
        x"61", x"62", x"63", x"62", x"61", x"61", x"62", x"61", x"61", x"60", x"60", x"60", x"60", x"61", x"61", 
        x"61", x"60", x"5f", x"5f", x"5f", x"60", x"61", x"61", x"61", x"60", x"60", x"60", x"5f", x"5f", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"5f", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", 
        x"63", x"63", x"63", x"64", x"64", x"64", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", 
        x"61", x"61", x"60", x"61", x"61", x"61", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"63", 
        x"63", x"64", x"65", x"64", x"62", x"62", x"62", x"62", x"63", x"63", x"64", x"64", x"64", x"64", x"64", 
        x"64", x"64", x"64", x"64", x"63", x"63", x"63", x"63", x"64", x"64", x"64", x"64", x"64", x"63", x"63", 
        x"63", x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"63", x"64", x"65", x"63", x"64", x"65", x"65", 
        x"64", x"63", x"64", x"67", x"67", x"65", x"64", x"65", x"66", x"65", x"67", x"67", x"64", x"69", x"67", 
        x"63", x"63", x"64", x"64", x"65", x"64", x"64", x"63", x"64", x"64", x"66", x"64", x"62", x"61", x"63", 
        x"65", x"65", x"64", x"66", x"66", x"66", x"68", x"68", x"64", x"66", x"66", x"67", x"66", x"67", x"66", 
        x"66", x"68", x"68", x"65", x"63", x"65", x"66", x"65", x"65", x"65", x"66", x"66", x"66", x"66", x"65", 
        x"65", x"66", x"68", x"67", x"65", x"65", x"67", x"66", x"62", x"65", x"66", x"63", x"63", x"65", x"64", 
        x"65", x"69", x"6c", x"68", x"66", x"69", x"6b", x"6b", x"68", x"69", x"67", x"69", x"66", x"65", x"63", 
        x"67", x"6a", x"6a", x"65", x"63", x"68", x"6e", x"68", x"67", x"73", x"6c", x"60", x"63", x"72", x"b0", 
        x"d8", x"a4", x"7f", x"a6", x"cf", x"cd", x"c9", x"c4", x"cc", x"ca", x"cf", x"d3", x"d0", x"cb", x"a6", 
        x"67", x"5e", x"5e", x"5e", x"5e", x"5c", x"5c", x"5e", x"5d", x"5e", x"5f", x"5f", x"5f", x"5d", x"5c", 
        x"60", x"5d", x"57", x"69", x"8b", x"b4", x"d7", x"ec", x"ee", x"cd", x"98", x"6a", x"63", x"60", x"63", 
        x"68", x"6b", x"6e", x"6e", x"6c", x"6e", x"6c", x"69", x"6d", x"6c", x"68", x"69", x"6b", x"6a", x"69", 
        x"69", x"6a", x"6b", x"6a", x"69", x"69", x"6a", x"6b", x"6b", x"6a", x"6b", x"6a", x"6a", x"6d", x"6c", 
        x"69", x"68", x"68", x"68", x"69", x"6a", x"6c", x"6c", x"6d", x"6c", x"6b", x"6b", x"6b", x"6a", x"6c", 
        x"6e", x"6c", x"6b", x"6c", x"6b", x"69", x"6b", x"6e", x"6d", x"6c", x"6c", x"6a", x"6b", x"6b", x"6b", 
        x"6b", x"6c", x"6d", x"6f", x"6e", x"6f", x"6d", x"6b", x"6d", x"6d", x"6e", x"6d", x"6b", x"6c", x"6b", 
        x"6b", x"6d", x"6b", x"6a", x"6c", x"6c", x"6d", x"6f", x"6e", x"6e", x"6d", x"6c", x"6c", x"6b", x"6c", 
        x"6c", x"6e", x"6c", x"6a", x"69", x"6b", x"6b", x"6a", x"6b", x"6b", x"6b", x"6b", x"6b", x"6c", x"6c", 
        x"6c", x"6e", x"6d", x"6c", x"6d", x"6d", x"6c", x"6d", x"6a", x"6a", x"6c", x"6e", x"6b", x"67", x"6c", 
        x"6c", x"6b", x"6c", x"6c", x"6b", x"6a", x"6b", x"6e", x"6e", x"6c", x"6c", x"6c", x"69", x"6c", x"6d", 
        x"6b", x"6d", x"6c", x"6d", x"6d", x"6b", x"6d", x"6b", x"6d", x"6a", x"66", x"6a", x"6b", x"6c", x"6b", 
        x"69", x"69", x"68", x"68", x"69", x"68", x"68", x"68", x"68", x"6b", x"6d", x"6c", x"6c", x"6c", x"6b", 
        x"6b", x"6c", x"6d", x"6c", x"6c", x"6d", x"6d", x"6e", x"6f", x"70", x"71", x"71", x"6f", x"6f", x"71", 
        x"70", x"6f", x"6e", x"6d", x"6d", x"6c", x"6b", x"6a", x"6b", x"6c", x"6b", x"68", x"68", x"68", x"68", 
        x"69", x"6b", x"6b", x"6c", x"6b", x"6e", x"6e", x"6c", x"6e", x"6d", x"70", x"6d", x"69", x"69", x"6a", 
        x"68", x"69", x"6a", x"6a", x"69", x"67", x"68", x"6b", x"68", x"67", x"69", x"69", x"68", x"67", x"68", 
        x"67", x"67", x"69", x"68", x"69", x"6a", x"6b", x"6a", x"68", x"69", x"68", x"68", x"69", x"6b", x"6a", 
        x"69", x"6c", x"6b", x"6a", x"69", x"69", x"6b", x"67", x"67", x"68", x"6b", x"67", x"69", x"69", x"69", 
        x"69", x"6a", x"69", x"6a", x"6b", x"67", x"65", x"66", x"66", x"67", x"67", x"67", x"69", x"6b", x"6e", 
        x"67", x"68", x"69", x"67", x"68", x"69", x"68", x"69", x"6a", x"69", x"68", x"6b", x"6b", x"66", x"68", 
        x"6a", x"69", x"67", x"67", x"69", x"69", x"69", x"66", x"64", x"64", x"66", x"67", x"66", x"67", x"68", 
        x"66", x"67", x"67", x"68", x"6a", x"67", x"64", x"65", x"66", x"68", x"69", x"69", x"6a", x"69", x"68", 
        x"67", x"65", x"68", x"68", x"66", x"67", x"69", x"67", x"68", x"68", x"68", x"69", x"6a", x"69", x"67", 
        x"65", x"68", x"69", x"66", x"66", x"68", x"68", x"64", x"63", x"62", x"63", x"66", x"67", x"66", x"66", 
        x"66", x"65", x"64", x"65", x"65", x"65", x"66", x"64", x"63", x"63", x"65", x"63", x"62", x"63", x"62", 
        x"61", x"61", x"63", x"65", x"64", x"63", x"64", x"64", x"62", x"63", x"65", x"65", x"65", x"67", x"65", 
        x"63", x"64", x"66", x"65", x"65", x"66", x"66", x"66", x"65", x"64", x"62", x"61", x"61", x"62", x"62", 
        x"64", x"65", x"65", x"63", x"65", x"65", x"63", x"64", x"62", x"64", x"65", x"63", x"63", x"66", x"66", 
        x"64", x"63", x"64", x"64", x"61", x"61", x"64", x"65", x"64", x"64", x"64", x"64", x"64", x"63", x"63", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"61", x"61", 
        x"61", x"61", x"62", x"62", x"61", x"61", x"62", x"62", x"60", x"60", x"5f", x"5f", x"60", x"60", x"61", 
        x"62", x"61", x"60", x"60", x"60", x"61", x"62", x"60", x"60", x"61", x"61", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"5f", x"60", x"60", x"60", x"61", x"60", x"60", x"5f", x"5f", x"5e", 
        x"63", x"64", x"65", x"64", x"63", x"63", x"64", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"60", 
        x"61", x"61", x"60", x"62", x"61", x"62", x"63", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"63", 
        x"63", x"64", x"65", x"64", x"62", x"63", x"63", x"63", x"63", x"63", x"64", x"64", x"64", x"64", x"64", 
        x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"63", x"63", x"62", x"63", x"64", x"64", x"63", 
        x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"64", x"63", x"64", x"64", x"64", x"64", x"65", 
        x"65", x"65", x"65", x"64", x"65", x"64", x"63", x"63", x"64", x"64", x"65", x"66", x"65", x"69", x"68", 
        x"65", x"64", x"64", x"66", x"67", x"66", x"64", x"63", x"63", x"62", x"61", x"62", x"64", x"63", x"64", 
        x"67", x"64", x"65", x"66", x"65", x"63", x"64", x"66", x"64", x"66", x"64", x"66", x"66", x"66", x"65", 
        x"65", x"67", x"68", x"64", x"64", x"67", x"64", x"62", x"64", x"64", x"64", x"64", x"64", x"63", x"63", 
        x"63", x"65", x"68", x"67", x"64", x"65", x"66", x"65", x"63", x"67", x"66", x"63", x"65", x"68", x"66", 
        x"63", x"66", x"6a", x"66", x"65", x"67", x"68", x"68", x"65", x"68", x"67", x"6b", x"68", x"68", x"67", 
        x"69", x"67", x"68", x"68", x"67", x"68", x"69", x"67", x"6a", x"6d", x"63", x"61", x"8d", x"be", x"c4", 
        x"98", x"8f", x"b7", x"ce", x"ce", x"c9", x"ca", x"c5", x"d0", x"cd", x"ce", x"d0", x"d1", x"cd", x"a6", 
        x"68", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5d", x"5d", x"5e", x"5d", x"5c", x"5e", 
        x"5d", x"5c", x"5c", x"60", x"63", x"6a", x"85", x"a6", x"c7", x"e1", x"e7", x"d2", x"a5", x"81", x"69", 
        x"60", x"61", x"6a", x"6d", x"6b", x"6d", x"6c", x"68", x"6a", x"6a", x"6c", x"6c", x"6b", x"6b", x"6a", 
        x"6a", x"6a", x"6a", x"6a", x"6a", x"69", x"69", x"6a", x"6a", x"6a", x"6b", x"6b", x"6a", x"6d", x"69", 
        x"69", x"69", x"68", x"69", x"6a", x"6b", x"6b", x"6b", x"6b", x"6b", x"6b", x"6b", x"6b", x"6b", x"6c", 
        x"6c", x"6c", x"6b", x"68", x"67", x"66", x"68", x"6a", x"6a", x"6a", x"6c", x"6d", x"6a", x"6a", x"6d", 
        x"6d", x"6b", x"6d", x"6f", x"6e", x"6e", x"6d", x"6b", x"6c", x"6e", x"6f", x"6f", x"6d", x"6e", x"6e", 
        x"6d", x"6f", x"6c", x"6c", x"6d", x"6c", x"6c", x"6d", x"6d", x"6d", x"6d", x"6d", x"6c", x"6c", x"6c", 
        x"6a", x"69", x"69", x"69", x"6b", x"6e", x"6f", x"6c", x"6b", x"6d", x"6e", x"6e", x"6e", x"6d", x"6c", 
        x"6b", x"6b", x"6a", x"6a", x"6b", x"6d", x"6f", x"70", x"6b", x"69", x"6c", x"6d", x"6c", x"6b", x"6c", 
        x"6a", x"69", x"6b", x"6b", x"6a", x"6a", x"6c", x"6f", x"6e", x"6e", x"70", x"6d", x"68", x"6c", x"6b", 
        x"68", x"6b", x"6b", x"6b", x"6b", x"6a", x"6b", x"6a", x"6e", x"6c", x"69", x"6d", x"6c", x"6d", x"6a", 
        x"68", x"68", x"67", x"68", x"68", x"67", x"69", x"6a", x"6a", x"6a", x"6c", x"6b", x"6a", x"6a", x"6b", 
        x"6c", x"6c", x"6c", x"6d", x"6c", x"6d", x"6e", x"6f", x"70", x"70", x"70", x"70", x"6f", x"6f", x"71", 
        x"6e", x"6f", x"71", x"6f", x"6e", x"6c", x"6b", x"6c", x"6d", x"6c", x"6b", x"6b", x"69", x"6b", x"6c", 
        x"6b", x"6c", x"6c", x"6c", x"6b", x"6d", x"6c", x"6d", x"6c", x"6c", x"6c", x"68", x"66", x"6a", x"6d", 
        x"69", x"69", x"6a", x"6c", x"6d", x"6c", x"6b", x"6c", x"6a", x"68", x"6a", x"6b", x"6c", x"6a", x"6a", 
        x"69", x"6a", x"69", x"69", x"6a", x"6b", x"6a", x"6a", x"69", x"69", x"69", x"69", x"6a", x"6c", x"6b", 
        x"69", x"68", x"67", x"6a", x"67", x"66", x"69", x"67", x"69", x"69", x"6c", x"68", x"6a", x"69", x"68", 
        x"68", x"67", x"67", x"69", x"6b", x"69", x"68", x"69", x"67", x"68", x"68", x"67", x"69", x"69", x"6c", 
        x"69", x"6a", x"6a", x"66", x"67", x"68", x"69", x"67", x"67", x"69", x"68", x"6b", x"6a", x"63", x"66", 
        x"69", x"69", x"67", x"67", x"69", x"68", x"69", x"66", x"65", x"65", x"67", x"68", x"68", x"68", x"68", 
        x"67", x"68", x"66", x"66", x"68", x"67", x"6a", x"6a", x"69", x"68", x"68", x"68", x"68", x"69", x"67", 
        x"66", x"66", x"68", x"68", x"68", x"66", x"66", x"64", x"65", x"65", x"64", x"66", x"67", x"66", x"65", 
        x"63", x"65", x"66", x"64", x"66", x"69", x"68", x"63", x"64", x"65", x"65", x"65", x"66", x"65", x"65", 
        x"66", x"65", x"63", x"66", x"65", x"64", x"65", x"65", x"64", x"65", x"67", x"66", x"65", x"65", x"64", 
        x"64", x"65", x"65", x"65", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"66", x"66", x"66", x"65", 
        x"64", x"65", x"65", x"63", x"65", x"66", x"67", x"66", x"64", x"63", x"64", x"63", x"63", x"62", x"62", 
        x"62", x"63", x"65", x"64", x"66", x"66", x"63", x"63", x"62", x"63", x"65", x"63", x"63", x"66", x"65", 
        x"63", x"63", x"64", x"64", x"61", x"61", x"64", x"64", x"63", x"64", x"64", x"63", x"63", x"63", x"62", 
        x"62", x"62", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"61", x"61", x"61", 
        x"62", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"61", x"5f", x"5e", x"5e", x"5f", x"61", x"60", 
        x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"60", x"61", x"61", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"61", x"60", x"5f", x"5e", x"5e", 
        x"62", x"64", x"65", x"64", x"63", x"63", x"64", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"63", 
        x"65", x"64", x"61", x"63", x"61", x"61", x"62", x"61", x"61", x"62", x"62", x"61", x"61", x"61", x"62", 
        x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"62", x"63", x"64", x"64", x"62", x"63", x"64", x"63", x"63", x"63", x"64", x"64", x"64", x"64", x"63", 
        x"63", x"63", x"64", x"63", x"63", x"62", x"63", x"63", x"63", x"62", x"62", x"63", x"64", x"65", x"63", 
        x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"63", x"63", x"63", x"63", x"64", x"64", x"64", x"65", 
        x"66", x"66", x"66", x"63", x"64", x"65", x"62", x"62", x"64", x"65", x"65", x"64", x"64", x"68", x"67", 
        x"66", x"67", x"66", x"66", x"67", x"66", x"65", x"64", x"64", x"63", x"63", x"65", x"67", x"65", x"64", 
        x"67", x"63", x"66", x"66", x"64", x"63", x"63", x"65", x"69", x"66", x"62", x"66", x"66", x"66", x"65", 
        x"67", x"68", x"66", x"65", x"67", x"69", x"63", x"62", x"67", x"67", x"66", x"65", x"66", x"66", x"66", 
        x"66", x"63", x"65", x"65", x"63", x"65", x"68", x"67", x"66", x"67", x"64", x"63", x"67", x"6b", x"67", 
        x"65", x"66", x"69", x"66", x"66", x"67", x"65", x"68", x"68", x"6a", x"68", x"6b", x"68", x"68", x"69", 
        x"6b", x"66", x"66", x"6a", x"69", x"66", x"64", x"69", x"6a", x"60", x"69", x"97", x"c7", x"bd", x"8f", 
        x"93", x"c6", x"d2", x"c6", x"c9", x"c7", x"ca", x"c5", x"cd", x"ca", x"cf", x"cc", x"cc", x"cd", x"a7", 
        x"68", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"5e", x"5d", x"5f", x"5e", x"5e", x"5e", x"5d", 
        x"5e", x"60", x"5e", x"5e", x"60", x"5f", x"5b", x"62", x"7c", x"a0", x"c7", x"e1", x"ec", x"d5", x"b1", 
        x"85", x"64", x"60", x"65", x"6b", x"6e", x"6a", x"67", x"6a", x"6a", x"6b", x"6d", x"6d", x"6c", x"6b", 
        x"6a", x"69", x"69", x"69", x"6a", x"6a", x"6b", x"6b", x"6a", x"69", x"6a", x"6c", x"6b", x"6d", x"69", 
        x"6c", x"6c", x"6a", x"69", x"69", x"69", x"6a", x"6a", x"6b", x"6c", x"6b", x"6b", x"6c", x"6d", x"6c", 
        x"6b", x"6d", x"6c", x"68", x"67", x"68", x"6a", x"6a", x"6a", x"6b", x"6a", x"6b", x"6a", x"6b", x"6d", 
        x"6d", x"6c", x"6c", x"6d", x"6b", x"6c", x"6b", x"6a", x"6d", x"6c", x"6e", x"6d", x"6c", x"6e", x"6e", 
        x"6d", x"6c", x"6b", x"6d", x"6e", x"6c", x"6b", x"6d", x"6e", x"6e", x"6d", x"6c", x"6b", x"6b", x"6a", 
        x"6b", x"6b", x"69", x"6a", x"6c", x"6d", x"6d", x"6b", x"6a", x"6c", x"6d", x"6b", x"6a", x"6a", x"6b", 
        x"6b", x"6a", x"6b", x"6b", x"6b", x"6d", x"70", x"6e", x"6b", x"6b", x"6c", x"6b", x"6a", x"6c", x"6d", 
        x"6a", x"69", x"6c", x"6c", x"6c", x"6e", x"6f", x"6f", x"6c", x"6d", x"70", x"6d", x"6a", x"6d", x"6a", 
        x"68", x"6b", x"6c", x"6c", x"6c", x"6b", x"69", x"6a", x"6f", x"6c", x"6c", x"70", x"6b", x"6e", x"6a", 
        x"69", x"6a", x"6a", x"6b", x"6c", x"6a", x"6b", x"6b", x"6a", x"6c", x"6c", x"69", x"6a", x"6b", x"6c", 
        x"6c", x"6b", x"6a", x"6a", x"6b", x"6c", x"6f", x"70", x"70", x"70", x"6f", x"6f", x"6e", x"70", x"73", 
        x"71", x"71", x"72", x"70", x"6f", x"6d", x"6d", x"6f", x"6e", x"6d", x"6c", x"6b", x"67", x"6c", x"6e", 
        x"6c", x"6b", x"6b", x"6b", x"6c", x"6c", x"6a", x"6c", x"69", x"69", x"6b", x"67", x"65", x"6b", x"6f", 
        x"6b", x"69", x"69", x"69", x"6b", x"6c", x"6b", x"6a", x"6a", x"69", x"6b", x"6d", x"6e", x"6b", x"6a", 
        x"69", x"69", x"6a", x"6b", x"6b", x"6a", x"69", x"6a", x"6a", x"69", x"69", x"69", x"6a", x"6b", x"6b", 
        x"69", x"6a", x"68", x"6d", x"6a", x"68", x"6c", x"6a", x"69", x"66", x"69", x"67", x"69", x"67", x"67", 
        x"68", x"66", x"66", x"68", x"6a", x"69", x"69", x"6a", x"6a", x"6a", x"6b", x"68", x"69", x"68", x"6a", 
        x"6b", x"6d", x"6e", x"68", x"6a", x"6a", x"69", x"67", x"69", x"6c", x"67", x"6a", x"6a", x"67", x"66", 
        x"67", x"6a", x"68", x"69", x"69", x"67", x"68", x"69", x"68", x"67", x"68", x"68", x"69", x"69", x"68", 
        x"68", x"69", x"66", x"65", x"68", x"68", x"6a", x"6a", x"68", x"67", x"67", x"68", x"68", x"6b", x"68", 
        x"66", x"67", x"68", x"68", x"6a", x"68", x"67", x"65", x"67", x"67", x"65", x"67", x"67", x"65", x"66", 
        x"65", x"65", x"66", x"64", x"65", x"69", x"6d", x"66", x"65", x"67", x"66", x"64", x"65", x"65", x"64", 
        x"67", x"66", x"63", x"67", x"65", x"63", x"65", x"67", x"67", x"67", x"67", x"68", x"67", x"65", x"65", 
        x"66", x"67", x"67", x"66", x"66", x"67", x"64", x"64", x"65", x"64", x"64", x"68", x"68", x"66", x"64", 
        x"64", x"64", x"63", x"62", x"64", x"65", x"65", x"65", x"63", x"62", x"62", x"62", x"63", x"63", x"64", 
        x"64", x"64", x"65", x"64", x"66", x"66", x"63", x"64", x"64", x"63", x"66", x"64", x"64", x"66", x"64", 
        x"62", x"63", x"63", x"63", x"61", x"61", x"64", x"63", x"62", x"64", x"64", x"63", x"62", x"62", x"63", 
        x"63", x"62", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"61", x"61", x"61", x"61", x"61", 
        x"63", x"61", x"60", x"61", x"61", x"61", x"61", x"62", x"61", x"5f", x"5e", x"5e", x"5f", x"60", x"60", 
        x"5f", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"60", x"60", x"61", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"61", x"61", x"60", x"5f", x"5f", x"5f", 
        x"63", x"63", x"65", x"65", x"64", x"62", x"63", x"62", x"62", x"63", x"63", x"63", x"63", x"62", x"62", 
        x"63", x"63", x"62", x"63", x"64", x"64", x"63", x"61", x"61", x"62", x"63", x"63", x"61", x"61", x"63", 
        x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", 
        x"62", x"63", x"63", x"63", x"62", x"64", x"64", x"62", x"63", x"63", x"63", x"63", x"63", x"62", x"62", 
        x"62", x"64", x"64", x"63", x"62", x"61", x"61", x"61", x"62", x"62", x"63", x"64", x"65", x"65", x"64", 
        x"63", x"64", x"63", x"63", x"62", x"62", x"63", x"63", x"63", x"63", x"64", x"64", x"63", x"63", x"64", 
        x"64", x"63", x"64", x"65", x"64", x"64", x"64", x"65", x"65", x"65", x"65", x"65", x"64", x"65", x"65", 
        x"65", x"66", x"66", x"65", x"66", x"64", x"64", x"63", x"64", x"65", x"65", x"64", x"66", x"66", x"66", 
        x"65", x"62", x"67", x"69", x"68", x"66", x"64", x"63", x"64", x"66", x"67", x"69", x"66", x"65", x"65", 
        x"66", x"65", x"66", x"65", x"65", x"66", x"64", x"65", x"66", x"66", x"65", x"66", x"65", x"67", x"68", 
        x"67", x"66", x"66", x"66", x"62", x"65", x"69", x"66", x"67", x"68", x"64", x"66", x"69", x"69", x"66", 
        x"67", x"67", x"67", x"66", x"68", x"6a", x"68", x"68", x"67", x"66", x"66", x"67", x"67", x"69", x"6a", 
        x"68", x"69", x"6a", x"66", x"68", x"67", x"67", x"67", x"5c", x"75", x"b2", x"d0", x"a1", x"87", x"ac", 
        x"d2", x"cf", x"ca", x"c8", x"c7", x"cb", x"cf", x"c8", x"cf", x"cf", x"ce", x"ce", x"ce", x"ca", x"a5", 
        x"67", x"5d", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5e", x"5f", 
        x"5e", x"5e", x"5c", x"5b", x"5a", x"5c", x"5f", x"5d", x"5e", x"62", x"73", x"8a", x"b4", x"d9", x"ef", 
        x"e8", x"c3", x"9b", x"71", x"5c", x"5f", x"67", x"6c", x"6c", x"69", x"6a", x"6b", x"6d", x"6b", x"6b", 
        x"6c", x"6b", x"6b", x"6a", x"68", x"69", x"6c", x"6d", x"6b", x"6a", x"68", x"6d", x"6c", x"6c", x"6c", 
        x"6d", x"6b", x"6c", x"69", x"6c", x"6d", x"6b", x"6d", x"6e", x"6d", x"6e", x"6c", x"6b", x"6c", x"6b", 
        x"6a", x"6d", x"6d", x"6b", x"6b", x"6c", x"6d", x"6d", x"6d", x"6e", x"6d", x"6d", x"6f", x"6d", x"69", 
        x"69", x"6c", x"6d", x"6e", x"6c", x"6c", x"6d", x"6b", x"6d", x"6e", x"6d", x"6e", x"6b", x"6b", x"6e", 
        x"6d", x"6d", x"6d", x"6e", x"6e", x"6b", x"6a", x"6d", x"6d", x"6a", x"6a", x"6c", x"6c", x"6b", x"6b", 
        x"6b", x"6b", x"6b", x"6d", x"6d", x"6c", x"6d", x"6d", x"6b", x"6b", x"6c", x"6b", x"6a", x"6a", x"6c", 
        x"6e", x"6c", x"6d", x"6c", x"6c", x"6e", x"6c", x"6b", x"6c", x"6c", x"6d", x"6c", x"6a", x"6a", x"6b", 
        x"69", x"6a", x"6a", x"6b", x"6d", x"6d", x"6f", x"6f", x"6c", x"6a", x"6d", x"6e", x"6c", x"6c", x"69", 
        x"69", x"6d", x"6e", x"6c", x"6b", x"6c", x"6c", x"6a", x"6d", x"6d", x"6b", x"6b", x"6a", x"69", x"6a", 
        x"6a", x"6a", x"6b", x"6c", x"6c", x"6d", x"6d", x"6d", x"6b", x"6c", x"6c", x"6c", x"6a", x"6a", x"6c", 
        x"6d", x"6d", x"6d", x"6c", x"6c", x"6a", x"6c", x"6e", x"6f", x"70", x"6f", x"6f", x"6e", x"6f", x"70", 
        x"6f", x"6f", x"70", x"70", x"6e", x"6e", x"6e", x"6f", x"6e", x"6c", x"6b", x"6c", x"69", x"6e", x"6e", 
        x"6b", x"6b", x"6a", x"6e", x"6d", x"6b", x"69", x"6a", x"6a", x"69", x"6a", x"69", x"67", x"6d", x"6f", 
        x"6c", x"6b", x"6b", x"6b", x"6e", x"6f", x"6d", x"6c", x"69", x"69", x"6b", x"6c", x"6b", x"6a", x"6b", 
        x"6a", x"69", x"69", x"68", x"69", x"68", x"6b", x"67", x"6a", x"6a", x"6b", x"6b", x"6b", x"6a", x"69", 
        x"69", x"6b", x"6d", x"70", x"6e", x"6d", x"6b", x"6a", x"6b", x"66", x"66", x"67", x"68", x"65", x"66", 
        x"68", x"68", x"69", x"69", x"67", x"66", x"66", x"67", x"67", x"68", x"69", x"69", x"67", x"67", x"6b", 
        x"6a", x"6a", x"6b", x"6b", x"6b", x"6b", x"6b", x"69", x"6b", x"6b", x"68", x"68", x"68", x"69", x"6a", 
        x"69", x"6b", x"6a", x"6a", x"68", x"67", x"6b", x"69", x"68", x"67", x"67", x"68", x"6a", x"6b", x"69", 
        x"69", x"6a", x"67", x"65", x"68", x"69", x"68", x"67", x"67", x"68", x"6a", x"6a", x"6a", x"6c", x"6c", 
        x"6c", x"69", x"6a", x"6a", x"68", x"68", x"6a", x"6a", x"6a", x"68", x"67", x"68", x"68", x"67", x"69", 
        x"69", x"67", x"67", x"67", x"66", x"68", x"6c", x"67", x"67", x"67", x"67", x"66", x"65", x"67", x"65", 
        x"65", x"66", x"66", x"67", x"65", x"65", x"64", x"64", x"68", x"69", x"66", x"64", x"64", x"64", x"65", 
        x"66", x"65", x"64", x"64", x"66", x"65", x"64", x"62", x"64", x"65", x"62", x"64", x"64", x"63", x"64", 
        x"65", x"65", x"64", x"63", x"65", x"65", x"65", x"62", x"62", x"62", x"65", x"65", x"65", x"66", x"64", 
        x"63", x"64", x"64", x"65", x"66", x"64", x"64", x"64", x"63", x"64", x"64", x"64", x"62", x"64", x"64", 
        x"63", x"63", x"63", x"64", x"64", x"64", x"65", x"64", x"64", x"64", x"64", x"64", x"63", x"63", x"63", 
        x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"61", x"61", x"62", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", 
        x"61", x"60", x"60", x"60", x"60", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", 
        x"5f", x"5f", x"5f", x"60", x"61", x"61", x"60", x"60", x"60", x"61", x"61", x"60", x"60", x"5f", x"5e", 
        x"64", x"64", x"65", x"66", x"64", x"62", x"63", x"63", x"63", x"63", x"63", x"62", x"63", x"62", x"62", 
        x"62", x"62", x"62", x"62", x"63", x"64", x"62", x"61", x"62", x"62", x"64", x"64", x"62", x"62", x"65", 
        x"64", x"62", x"62", x"62", x"63", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"63", x"62", x"62", 
        x"62", x"63", x"62", x"61", x"61", x"65", x"64", x"63", x"63", x"63", x"62", x"63", x"64", x"64", x"64", 
        x"63", x"63", x"64", x"61", x"60", x"62", x"62", x"61", x"62", x"63", x"64", x"64", x"65", x"65", x"64", 
        x"64", x"64", x"65", x"65", x"64", x"64", x"64", x"63", x"63", x"62", x"63", x"65", x"64", x"64", x"66", 
        x"64", x"62", x"63", x"66", x"65", x"64", x"66", x"67", x"66", x"64", x"64", x"63", x"62", x"64", x"66", 
        x"65", x"67", x"68", x"66", x"66", x"65", x"63", x"63", x"63", x"64", x"63", x"63", x"64", x"66", x"67", 
        x"65", x"62", x"62", x"65", x"67", x"65", x"65", x"66", x"65", x"67", x"69", x"68", x"65", x"65", x"67", 
        x"66", x"64", x"65", x"65", x"64", x"65", x"67", x"67", x"65", x"66", x"66", x"67", x"66", x"68", x"69", 
        x"68", x"67", x"67", x"69", x"66", x"66", x"69", x"66", x"67", x"69", x"66", x"69", x"6a", x"67", x"67", 
        x"67", x"67", x"68", x"69", x"6b", x"6b", x"6a", x"69", x"65", x"66", x"67", x"68", x"68", x"68", x"6b", 
        x"6b", x"68", x"69", x"66", x"66", x"6a", x"65", x"68", x"87", x"bf", x"c0", x"97", x"94", x"b7", x"ce", 
        x"cf", x"cc", x"ce", x"cc", x"ca", x"c8", x"cb", x"c8", x"cc", x"ce", x"cd", x"ce", x"ce", x"c9", x"a4", 
        x"67", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"60", x"6d", x"8a", x"ab", 
        x"cb", x"e5", x"e4", x"cc", x"a1", x"7f", x"68", x"64", x"67", x"67", x"6a", x"6a", x"6a", x"6b", x"6e", 
        x"6b", x"6c", x"6d", x"6c", x"6b", x"6a", x"6c", x"6b", x"6c", x"6f", x"6d", x"6e", x"6d", x"6d", x"6e", 
        x"6c", x"69", x"6b", x"68", x"6d", x"6e", x"6b", x"6c", x"6e", x"6b", x"6e", x"6d", x"6c", x"6d", x"6c", 
        x"6b", x"6c", x"6b", x"6b", x"6b", x"6c", x"6d", x"6e", x"6f", x"6f", x"6e", x"6e", x"70", x"6f", x"6b", 
        x"6a", x"6d", x"70", x"6f", x"6d", x"6c", x"6d", x"6b", x"6e", x"6f", x"6e", x"6f", x"6c", x"6a", x"6e", 
        x"6f", x"6f", x"6e", x"6e", x"6e", x"6b", x"6a", x"6d", x"6e", x"6c", x"6c", x"6d", x"6e", x"6d", x"6c", 
        x"6c", x"6d", x"6e", x"6d", x"6c", x"6d", x"70", x"6f", x"6b", x"6b", x"6c", x"6d", x"6d", x"6d", x"6e", 
        x"6e", x"6d", x"6c", x"6a", x"6b", x"6d", x"67", x"69", x"6d", x"6c", x"6e", x"70", x"6c", x"6c", x"70", 
        x"6f", x"70", x"6e", x"6b", x"6c", x"6b", x"6d", x"6f", x"6d", x"69", x"6a", x"6d", x"6d", x"6b", x"6a", 
        x"6b", x"6e", x"6e", x"6a", x"6a", x"6d", x"6e", x"6c", x"6d", x"6d", x"69", x"68", x"6a", x"6a", x"6d", 
        x"6d", x"6b", x"6c", x"6d", x"6c", x"6c", x"6c", x"6e", x"6a", x"6a", x"6a", x"6e", x"6d", x"6c", x"6c", 
        x"6c", x"6c", x"6b", x"69", x"6b", x"6b", x"6b", x"6a", x"6a", x"6c", x"6b", x"6d", x"6e", x"6e", x"6e", 
        x"6e", x"6f", x"6f", x"70", x"72", x"72", x"71", x"70", x"6f", x"6f", x"6f", x"6e", x"6c", x"6d", x"6e", 
        x"6e", x"6d", x"6b", x"6e", x"6c", x"6a", x"6a", x"6b", x"6d", x"6c", x"6a", x"69", x"69", x"6d", x"6d", 
        x"6a", x"68", x"6a", x"6c", x"6c", x"6b", x"6b", x"6b", x"6b", x"6b", x"6b", x"6b", x"6b", x"6c", x"6d", 
        x"6c", x"6a", x"6a", x"68", x"68", x"67", x"6c", x"67", x"6b", x"6d", x"6d", x"6d", x"6c", x"6b", x"6b", 
        x"6d", x"6b", x"6d", x"6e", x"6c", x"6b", x"69", x"6a", x"6c", x"69", x"67", x"6a", x"6a", x"67", x"68", 
        x"6a", x"6b", x"6e", x"6b", x"68", x"68", x"69", x"68", x"69", x"68", x"69", x"69", x"66", x"67", x"6b", 
        x"69", x"68", x"68", x"6c", x"6b", x"6a", x"6b", x"69", x"6b", x"6b", x"6a", x"6a", x"69", x"6b", x"6c", 
        x"6a", x"6b", x"69", x"6a", x"68", x"68", x"6c", x"68", x"69", x"69", x"69", x"68", x"67", x"68", x"6a", 
        x"6a", x"69", x"66", x"64", x"65", x"66", x"69", x"68", x"68", x"69", x"6a", x"68", x"67", x"69", x"6b", 
        x"6c", x"69", x"6b", x"6a", x"66", x"68", x"6a", x"6a", x"6a", x"68", x"68", x"68", x"68", x"68", x"6a", 
        x"6a", x"68", x"68", x"69", x"67", x"66", x"68", x"64", x"67", x"66", x"66", x"67", x"68", x"67", x"67", 
        x"66", x"65", x"66", x"67", x"65", x"66", x"65", x"64", x"68", x"6a", x"66", x"64", x"65", x"65", x"66", 
        x"66", x"65", x"64", x"63", x"64", x"64", x"65", x"62", x"65", x"68", x"63", x"64", x"63", x"63", x"63", 
        x"64", x"63", x"63", x"63", x"65", x"64", x"64", x"61", x"63", x"62", x"65", x"67", x"65", x"66", x"65", 
        x"62", x"65", x"63", x"65", x"65", x"64", x"64", x"64", x"62", x"64", x"63", x"65", x"62", x"63", x"65", 
        x"64", x"64", x"63", x"63", x"63", x"64", x"65", x"66", x"65", x"63", x"65", x"65", x"63", x"64", x"62", 
        x"62", x"63", x"64", x"64", x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"62", x"63", x"63", x"62", x"61", x"61", x"62", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", 
        x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"61", x"5f", 
        x"5f", x"5f", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5f", 
        x"65", x"67", x"67", x"66", x"64", x"63", x"63", x"63", x"63", x"63", x"62", x"62", x"62", x"63", x"63", 
        x"61", x"62", x"62", x"62", x"62", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"62", x"62", x"65", 
        x"64", x"62", x"61", x"62", x"64", x"65", x"65", x"65", x"65", x"65", x"65", x"65", x"65", x"63", x"63", 
        x"63", x"63", x"62", x"61", x"61", x"64", x"63", x"63", x"64", x"63", x"62", x"64", x"64", x"63", x"63", 
        x"63", x"64", x"65", x"63", x"61", x"62", x"61", x"61", x"63", x"64", x"65", x"65", x"65", x"65", x"64", 
        x"64", x"64", x"65", x"65", x"64", x"64", x"63", x"63", x"62", x"62", x"62", x"65", x"64", x"65", x"66", 
        x"65", x"62", x"61", x"65", x"66", x"65", x"66", x"67", x"66", x"65", x"64", x"63", x"62", x"64", x"65", 
        x"65", x"67", x"67", x"65", x"65", x"66", x"66", x"66", x"66", x"65", x"64", x"63", x"64", x"64", x"65", 
        x"65", x"64", x"64", x"66", x"65", x"63", x"64", x"66", x"66", x"67", x"68", x"67", x"64", x"65", x"66", 
        x"66", x"64", x"63", x"65", x"65", x"66", x"68", x"66", x"65", x"66", x"67", x"67", x"68", x"68", x"67", 
        x"68", x"69", x"68", x"6a", x"69", x"67", x"67", x"66", x"66", x"68", x"66", x"68", x"69", x"67", x"66", 
        x"68", x"69", x"6a", x"6a", x"6b", x"6b", x"6b", x"6a", x"68", x"69", x"6b", x"6b", x"68", x"68", x"6c", 
        x"6d", x"69", x"66", x"69", x"69", x"60", x"62", x"9a", x"d1", x"b6", x"8a", x"9f", x"c3", x"d2", x"ca", 
        x"cb", x"cc", x"cf", x"cd", x"cb", x"c8", x"cb", x"c7", x"cb", x"cc", x"cc", x"ce", x"cf", x"c9", x"a4", 
        x"67", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", x"64", 
        x"7a", x"a1", x"c8", x"eb", x"ea", x"d7", x"b5", x"84", x"63", x"5a", x"67", x"6d", x"6d", x"6a", x"6a", 
        x"68", x"6a", x"69", x"6d", x"71", x"6d", x"6d", x"6a", x"69", x"6e", x"6d", x"6f", x"6e", x"6e", x"6c", 
        x"6b", x"6b", x"69", x"68", x"6b", x"6c", x"6c", x"6b", x"6a", x"6a", x"6c", x"6c", x"6b", x"69", x"69", 
        x"6a", x"6b", x"6b", x"6b", x"6b", x"6c", x"6c", x"6d", x"6d", x"6f", x"6e", x"6d", x"6f", x"6f", x"6d", 
        x"6c", x"6e", x"6e", x"6d", x"6c", x"6a", x"6c", x"6b", x"6d", x"70", x"6f", x"6f", x"6c", x"6a", x"6d", 
        x"6d", x"6c", x"6c", x"6d", x"6d", x"6c", x"6b", x"6c", x"6d", x"6e", x"6f", x"6d", x"6f", x"70", x"6d", 
        x"6b", x"6d", x"6e", x"6e", x"6d", x"6d", x"6e", x"6d", x"6b", x"6a", x"6b", x"6d", x"6f", x"6e", x"6e", 
        x"6c", x"6b", x"6c", x"6b", x"6c", x"6d", x"68", x"69", x"6c", x"6c", x"6e", x"6f", x"6d", x"6d", x"6f", 
        x"6c", x"6d", x"6d", x"6a", x"69", x"69", x"6c", x"6f", x"6d", x"6a", x"69", x"6b", x"6d", x"6d", x"6c", 
        x"6d", x"6e", x"6e", x"6b", x"6b", x"6d", x"6e", x"6e", x"6d", x"6b", x"6b", x"6a", x"6a", x"6d", x"6d", 
        x"6b", x"69", x"6a", x"6c", x"6b", x"6c", x"6c", x"6d", x"6a", x"6b", x"6a", x"6b", x"6b", x"6b", x"6b", 
        x"6c", x"6c", x"6c", x"6a", x"6b", x"6c", x"6c", x"6a", x"6a", x"6d", x"6d", x"6e", x"6d", x"6e", x"6f", 
        x"70", x"70", x"70", x"72", x"74", x"73", x"71", x"70", x"70", x"72", x"73", x"70", x"6d", x"6c", x"6d", 
        x"6f", x"6c", x"6b", x"6c", x"6a", x"69", x"6a", x"6d", x"6c", x"6b", x"6b", x"6b", x"6c", x"6d", x"6d", 
        x"6a", x"6a", x"6d", x"6d", x"6b", x"68", x"68", x"6b", x"6e", x"6e", x"6b", x"68", x"6a", x"6d", x"6c", 
        x"69", x"6a", x"6c", x"6b", x"69", x"66", x"6b", x"6a", x"6d", x"6a", x"6a", x"6c", x"6c", x"6c", x"6c", 
        x"6d", x"6b", x"6a", x"6a", x"69", x"68", x"69", x"6a", x"6b", x"6a", x"69", x"6a", x"6b", x"6a", x"6b", 
        x"6c", x"6c", x"6d", x"6b", x"6a", x"6b", x"6b", x"6a", x"6d", x"6b", x"6a", x"69", x"65", x"67", x"6a", 
        x"6b", x"68", x"67", x"6a", x"69", x"68", x"68", x"68", x"6a", x"68", x"67", x"69", x"68", x"69", x"6a", 
        x"69", x"6a", x"69", x"6a", x"68", x"69", x"6c", x"69", x"6a", x"6a", x"6a", x"68", x"67", x"67", x"6a", 
        x"6a", x"6a", x"67", x"65", x"64", x"65", x"67", x"6a", x"6a", x"69", x"6b", x"6a", x"67", x"69", x"6a", 
        x"6a", x"6b", x"6c", x"6b", x"69", x"68", x"68", x"68", x"68", x"68", x"69", x"69", x"67", x"67", x"69", 
        x"69", x"69", x"68", x"67", x"66", x"63", x"65", x"63", x"67", x"67", x"67", x"68", x"69", x"67", x"68", 
        x"68", x"65", x"64", x"68", x"67", x"67", x"67", x"68", x"67", x"65", x"64", x"65", x"66", x"66", x"66", 
        x"66", x"66", x"66", x"64", x"65", x"65", x"65", x"64", x"65", x"67", x"65", x"66", x"64", x"63", x"63", 
        x"64", x"63", x"63", x"65", x"65", x"64", x"64", x"63", x"65", x"65", x"65", x"68", x"65", x"64", x"64", 
        x"63", x"65", x"62", x"61", x"63", x"65", x"64", x"63", x"62", x"64", x"64", x"66", x"64", x"65", x"65", 
        x"64", x"66", x"66", x"65", x"64", x"64", x"67", x"68", x"68", x"63", x"64", x"64", x"63", x"64", x"62", 
        x"62", x"63", x"64", x"64", x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"62", x"63", x"63", x"62", x"61", x"61", x"62", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"61", x"61", x"61", x"60", x"60", x"60", x"5f", 
        x"5f", x"5f", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5f", 
        x"64", x"67", x"67", x"64", x"63", x"64", x"63", x"63", x"64", x"63", x"63", x"63", x"63", x"63", x"64", 
        x"64", x"63", x"62", x"61", x"61", x"61", x"62", x"64", x"64", x"64", x"64", x"63", x"61", x"61", x"64", 
        x"63", x"62", x"62", x"63", x"64", x"66", x"66", x"66", x"66", x"66", x"66", x"66", x"65", x"64", x"64", 
        x"64", x"64", x"63", x"63", x"63", x"64", x"63", x"63", x"64", x"63", x"63", x"66", x"64", x"62", x"63", 
        x"63", x"65", x"66", x"65", x"63", x"63", x"63", x"63", x"63", x"64", x"64", x"65", x"65", x"65", x"65", 
        x"65", x"65", x"65", x"64", x"62", x"62", x"62", x"63", x"64", x"64", x"63", x"65", x"65", x"65", x"66", 
        x"66", x"63", x"61", x"64", x"65", x"65", x"65", x"65", x"64", x"64", x"65", x"66", x"65", x"65", x"65", 
        x"64", x"65", x"65", x"65", x"64", x"65", x"67", x"69", x"69", x"68", x"66", x"65", x"65", x"64", x"64", 
        x"66", x"68", x"65", x"66", x"66", x"64", x"66", x"67", x"66", x"68", x"69", x"68", x"66", x"67", x"68", 
        x"68", x"69", x"67", x"68", x"66", x"66", x"68", x"66", x"67", x"67", x"68", x"66", x"68", x"68", x"66", 
        x"69", x"6a", x"66", x"68", x"69", x"66", x"65", x"68", x"66", x"67", x"66", x"68", x"68", x"67", x"66", 
        x"68", x"68", x"68", x"67", x"67", x"68", x"6a", x"6b", x"6a", x"6a", x"6c", x"6c", x"68", x"68", x"6a", 
        x"6b", x"70", x"6d", x"66", x"63", x"72", x"b1", x"c9", x"a4", x"8a", x"b4", x"cc", x"ce", x"cb", x"cc", 
        x"cd", x"ca", x"ca", x"c9", x"cb", x"ca", x"cf", x"ca", x"ce", x"ce", x"cd", x"cf", x"d0", x"cb", x"a5", 
        x"68", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5f", x"5f", x"5e", x"5d", x"5d", x"5d", x"5e", 
        x"5d", x"61", x"74", x"91", x"bc", x"d8", x"e6", x"dd", x"be", x"95", x"69", x"63", x"6d", x"6c", x"6d", 
        x"6c", x"6a", x"6c", x"6e", x"67", x"6a", x"6e", x"6f", x"6e", x"72", x"6e", x"6b", x"6b", x"6c", x"69", 
        x"6a", x"6d", x"69", x"6c", x"6c", x"6f", x"71", x"70", x"6e", x"70", x"6e", x"6e", x"6f", x"6d", x"6c", 
        x"6d", x"6d", x"6e", x"6e", x"6d", x"6d", x"6c", x"6b", x"6a", x"6d", x"6d", x"6c", x"6f", x"70", x"6e", 
        x"6e", x"6f", x"6c", x"6d", x"6e", x"6d", x"6d", x"6a", x"6b", x"6c", x"6c", x"6c", x"6c", x"6d", x"70", 
        x"71", x"6d", x"6d", x"6e", x"6e", x"6d", x"6c", x"6c", x"6d", x"6e", x"6d", x"6b", x"6d", x"6e", x"6d", 
        x"6c", x"6c", x"6d", x"6d", x"6e", x"6d", x"6b", x"6c", x"6e", x"6b", x"6b", x"6d", x"6f", x"6e", x"6d", 
        x"6e", x"6e", x"6e", x"6e", x"6d", x"6d", x"6a", x"69", x"6a", x"6c", x"6d", x"6e", x"6d", x"6c", x"6d", 
        x"6a", x"6c", x"6e", x"6b", x"6b", x"6b", x"6c", x"6e", x"6e", x"6c", x"6a", x"6b", x"6c", x"6c", x"6c", 
        x"6e", x"6f", x"6e", x"6c", x"6b", x"6c", x"6d", x"6d", x"6c", x"6c", x"6d", x"6d", x"6c", x"6b", x"6a", 
        x"69", x"69", x"6b", x"6c", x"6c", x"6c", x"6b", x"6d", x"6d", x"6f", x"6f", x"6f", x"6c", x"6b", x"6b", 
        x"6d", x"6f", x"70", x"6f", x"6e", x"6c", x"6e", x"6d", x"6e", x"70", x"6e", x"6f", x"6d", x"6c", x"6c", 
        x"6d", x"6f", x"70", x"72", x"70", x"6f", x"6e", x"6d", x"6e", x"70", x"72", x"6e", x"6f", x"6c", x"6d", 
        x"6f", x"6c", x"6d", x"6d", x"6e", x"6a", x"6a", x"6d", x"6a", x"6a", x"6b", x"6c", x"6d", x"6d", x"6c", 
        x"6c", x"6d", x"6e", x"6c", x"6b", x"6a", x"6a", x"6b", x"6d", x"6e", x"6d", x"69", x"69", x"6b", x"6b", 
        x"6b", x"6c", x"6d", x"6e", x"6c", x"68", x"6b", x"6d", x"6e", x"68", x"68", x"6b", x"6d", x"6c", x"6a", 
        x"68", x"6a", x"69", x"6a", x"6c", x"6b", x"6c", x"6b", x"69", x"6b", x"6a", x"6a", x"6a", x"6b", x"6c", 
        x"6c", x"6c", x"6d", x"6b", x"6a", x"6a", x"6a", x"68", x"6a", x"69", x"6a", x"6a", x"67", x"67", x"6b", 
        x"6c", x"69", x"67", x"6a", x"6a", x"68", x"68", x"6b", x"6c", x"69", x"69", x"6b", x"69", x"68", x"6a", 
        x"6a", x"6a", x"6a", x"6a", x"6a", x"6a", x"6b", x"69", x"68", x"68", x"69", x"69", x"6a", x"69", x"69", 
        x"6b", x"6b", x"6a", x"69", x"68", x"66", x"65", x"68", x"68", x"67", x"6a", x"6b", x"67", x"68", x"68", 
        x"68", x"6a", x"6a", x"69", x"67", x"68", x"68", x"67", x"67", x"68", x"69", x"68", x"65", x"65", x"67", 
        x"66", x"68", x"66", x"65", x"65", x"63", x"65", x"66", x"6a", x"6a", x"69", x"6a", x"68", x"69", x"68", 
        x"65", x"66", x"66", x"66", x"65", x"65", x"66", x"68", x"68", x"67", x"68", x"67", x"67", x"67", x"67", 
        x"67", x"67", x"67", x"66", x"66", x"65", x"66", x"64", x"64", x"65", x"65", x"66", x"63", x"63", x"64", 
        x"65", x"65", x"64", x"64", x"63", x"63", x"62", x"62", x"64", x"64", x"65", x"69", x"66", x"64", x"65", 
        x"65", x"66", x"64", x"63", x"64", x"66", x"66", x"64", x"66", x"65", x"65", x"65", x"65", x"65", x"65", 
        x"65", x"66", x"66", x"65", x"63", x"63", x"65", x"66", x"66", x"64", x"64", x"64", x"63", x"64", x"62", 
        x"63", x"63", x"64", x"64", x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"62", x"63", x"62", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"60", x"60", x"60", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"61", x"62", x"61", x"60", x"60", x"60", x"61", 
        x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5f", 
        x"63", x"65", x"65", x"62", x"63", x"64", x"64", x"64", x"64", x"64", x"64", x"63", x"63", x"63", x"64", 
        x"64", x"63", x"62", x"62", x"61", x"61", x"61", x"61", x"62", x"64", x"64", x"65", x"64", x"64", x"63", 
        x"63", x"64", x"64", x"65", x"65", x"65", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"63", x"62", 
        x"62", x"63", x"64", x"65", x"66", x"66", x"64", x"63", x"63", x"63", x"63", x"67", x"65", x"63", x"64", 
        x"63", x"64", x"65", x"65", x"65", x"66", x"65", x"64", x"63", x"62", x"62", x"63", x"64", x"65", x"65", 
        x"65", x"65", x"65", x"64", x"63", x"62", x"61", x"63", x"65", x"64", x"64", x"66", x"66", x"65", x"64", 
        x"65", x"65", x"63", x"64", x"65", x"64", x"64", x"63", x"63", x"63", x"64", x"64", x"65", x"64", x"65", 
        x"65", x"66", x"66", x"68", x"66", x"65", x"67", x"68", x"69", x"69", x"66", x"68", x"68", x"66", x"65", 
        x"67", x"6a", x"66", x"67", x"67", x"66", x"67", x"68", x"66", x"66", x"66", x"65", x"66", x"66", x"66", 
        x"67", x"69", x"68", x"69", x"67", x"65", x"66", x"65", x"67", x"67", x"68", x"66", x"68", x"68", x"67", 
        x"6a", x"69", x"65", x"66", x"69", x"67", x"65", x"6a", x"67", x"67", x"67", x"68", x"67", x"67", x"66", 
        x"66", x"67", x"69", x"69", x"69", x"68", x"68", x"68", x"67", x"67", x"69", x"6a", x"6a", x"6b", x"6c", 
        x"6c", x"6e", x"67", x"63", x"89", x"c2", x"c5", x"90", x"8e", x"c5", x"cf", x"ca", x"c8", x"c9", x"ca", 
        x"cd", x"cb", x"cb", x"ca", x"cd", x"cc", x"d0", x"cc", x"ce", x"ce", x"cc", x"cf", x"d0", x"cb", x"a5", 
        x"68", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", 
        x"5d", x"5d", x"5f", x"63", x"6c", x"88", x"af", x"d4", x"e6", x"e5", x"ce", x"a4", x"79", x"61", x"66", 
        x"69", x"6a", x"6d", x"6d", x"68", x"6b", x"6f", x"6d", x"6c", x"6f", x"6d", x"6e", x"6e", x"6f", x"6d", 
        x"6d", x"70", x"6c", x"6c", x"6a", x"6c", x"6f", x"6f", x"6d", x"6f", x"6b", x"6c", x"6d", x"6b", x"6a", 
        x"6b", x"6b", x"6d", x"6e", x"6d", x"6d", x"6c", x"6b", x"6b", x"6c", x"6c", x"6c", x"70", x"72", x"6f", 
        x"6e", x"6e", x"6d", x"6e", x"6f", x"6e", x"6f", x"6c", x"6e", x"71", x"70", x"6d", x"6c", x"6c", x"6b", 
        x"6c", x"6e", x"6f", x"6f", x"6f", x"6e", x"6e", x"6d", x"6f", x"6d", x"6b", x"6b", x"6c", x"6d", x"6e", 
        x"71", x"70", x"6c", x"6a", x"6b", x"6d", x"6e", x"6f", x"6f", x"6c", x"6c", x"6d", x"6f", x"6e", x"6d", 
        x"6e", x"6e", x"6e", x"6e", x"6d", x"6c", x"6e", x"6c", x"6d", x"6f", x"70", x"6f", x"6e", x"6d", x"6e", 
        x"6b", x"6d", x"70", x"6e", x"6f", x"70", x"6e", x"6d", x"6e", x"6e", x"6d", x"6b", x"6a", x"69", x"69", 
        x"6c", x"6e", x"6d", x"6c", x"6b", x"6c", x"6d", x"6c", x"6d", x"6e", x"6d", x"6d", x"6d", x"6b", x"6b", 
        x"6c", x"6d", x"6e", x"6f", x"70", x"6f", x"6d", x"6e", x"6e", x"70", x"6e", x"6c", x"6d", x"6e", x"6d", 
        x"6e", x"6e", x"6e", x"6c", x"6b", x"6a", x"6c", x"6c", x"6c", x"6d", x"6c", x"6d", x"6c", x"6b", x"6b", 
        x"6c", x"6e", x"70", x"71", x"70", x"6f", x"6f", x"6f", x"6f", x"71", x"71", x"6e", x"71", x"6f", x"6e", 
        x"6d", x"6a", x"6e", x"70", x"70", x"6b", x"6a", x"6c", x"6b", x"6c", x"6d", x"6f", x"6f", x"6d", x"6b", 
        x"6c", x"6c", x"6d", x"6d", x"6d", x"6c", x"6b", x"6c", x"6c", x"6d", x"6e", x"6d", x"6b", x"6b", x"6e", 
        x"6e", x"6d", x"6c", x"6e", x"6e", x"6b", x"6c", x"6e", x"6d", x"6c", x"6c", x"6b", x"6c", x"6b", x"6b", 
        x"6b", x"6b", x"6a", x"6b", x"6e", x"6d", x"6e", x"6b", x"6a", x"6c", x"6c", x"6b", x"6b", x"6b", x"6b", 
        x"6c", x"6d", x"6e", x"6b", x"69", x"69", x"69", x"67", x"68", x"68", x"6a", x"6c", x"6a", x"68", x"6b", 
        x"6c", x"68", x"66", x"6b", x"6b", x"6a", x"6a", x"6c", x"6d", x"6a", x"6a", x"6d", x"6c", x"6b", x"6a", 
        x"6a", x"69", x"69", x"6a", x"6b", x"6b", x"69", x"68", x"69", x"69", x"6a", x"6a", x"69", x"68", x"67", 
        x"68", x"6a", x"6b", x"6a", x"69", x"67", x"69", x"6a", x"68", x"66", x"67", x"69", x"68", x"68", x"69", 
        x"67", x"6a", x"69", x"67", x"66", x"67", x"68", x"67", x"67", x"68", x"67", x"66", x"65", x"67", x"68", 
        x"66", x"69", x"67", x"65", x"67", x"67", x"68", x"68", x"69", x"69", x"66", x"66", x"65", x"67", x"67", 
        x"65", x"65", x"66", x"65", x"65", x"67", x"66", x"65", x"67", x"68", x"68", x"66", x"66", x"67", x"68", 
        x"68", x"67", x"66", x"66", x"66", x"65", x"65", x"66", x"64", x"65", x"65", x"64", x"63", x"63", x"64", 
        x"66", x"67", x"66", x"65", x"65", x"66", x"66", x"67", x"66", x"65", x"63", x"68", x"67", x"65", x"66", 
        x"65", x"66", x"65", x"64", x"64", x"65", x"65", x"65", x"67", x"65", x"64", x"64", x"64", x"64", x"64", 
        x"64", x"64", x"65", x"64", x"64", x"63", x"63", x"63", x"64", x"65", x"65", x"64", x"63", x"64", x"64", 
        x"65", x"64", x"64", x"64", x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"63", x"63", x"62", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"60", x"60", x"60", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"61", x"62", x"61", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5f", 
        x"64", x"64", x"63", x"63", x"64", x"65", x"65", x"64", x"64", x"64", x"64", x"64", x"63", x"63", x"63", 
        x"62", x"62", x"62", x"62", x"63", x"63", x"62", x"62", x"63", x"64", x"64", x"64", x"63", x"63", x"62", 
        x"63", x"64", x"65", x"65", x"65", x"65", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"62", x"62", 
        x"62", x"62", x"64", x"65", x"67", x"68", x"65", x"62", x"63", x"64", x"65", x"66", x"65", x"65", x"65", 
        x"63", x"62", x"63", x"64", x"64", x"64", x"64", x"64", x"63", x"63", x"64", x"65", x"64", x"65", x"65", 
        x"65", x"65", x"65", x"64", x"66", x"64", x"62", x"63", x"65", x"64", x"62", x"64", x"66", x"65", x"64", 
        x"64", x"66", x"65", x"64", x"65", x"64", x"64", x"63", x"63", x"64", x"64", x"64", x"66", x"65", x"65", 
        x"66", x"66", x"66", x"67", x"65", x"65", x"65", x"68", x"6a", x"69", x"66", x"67", x"68", x"68", x"66", 
        x"67", x"69", x"68", x"68", x"67", x"65", x"68", x"69", x"68", x"66", x"65", x"65", x"67", x"67", x"66", 
        x"67", x"68", x"66", x"67", x"68", x"67", x"65", x"64", x"66", x"68", x"67", x"66", x"67", x"68", x"69", 
        x"6a", x"67", x"65", x"66", x"6b", x"68", x"64", x"69", x"67", x"67", x"69", x"69", x"66", x"69", x"67", 
        x"68", x"6a", x"6b", x"6a", x"68", x"69", x"6b", x"69", x"68", x"68", x"68", x"69", x"6b", x"6c", x"6a", 
        x"67", x"62", x"69", x"99", x"c6", x"bb", x"8e", x"a0", x"cb", x"d4", x"ce", x"cc", x"cd", x"ce", x"cc", 
        x"cc", x"ca", x"cb", x"cb", x"cd", x"cc", x"cd", x"c8", x"cb", x"cc", x"cc", x"cf", x"d0", x"cb", x"a6", 
        x"69", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5d", x"5d", x"5c", x"5e", x"5f", 
        x"5f", x"5e", x"5f", x"60", x"5d", x"5d", x"66", x"7e", x"a2", x"c7", x"e1", x"e6", x"d6", x"aa", x"82", 
        x"6c", x"69", x"69", x"6c", x"6f", x"6f", x"70", x"6c", x"6c", x"71", x"71", x"71", x"70", x"70", x"6e", 
        x"6e", x"6e", x"6c", x"6d", x"6a", x"6a", x"6d", x"6d", x"6b", x"6c", x"6e", x"6f", x"70", x"6e", x"6e", 
        x"6e", x"6e", x"6d", x"6c", x"6c", x"6d", x"6d", x"6e", x"6e", x"6e", x"6b", x"6c", x"70", x"71", x"6e", 
        x"6d", x"6f", x"6f", x"6e", x"6e", x"6d", x"6f", x"6e", x"70", x"6e", x"6e", x"6b", x"6d", x"6f", x"6d", 
        x"6e", x"6f", x"70", x"6f", x"6e", x"6f", x"6f", x"6d", x"70", x"6d", x"6c", x"6d", x"6e", x"6d", x"6e", 
        x"71", x"71", x"6f", x"6d", x"6e", x"6f", x"6f", x"70", x"71", x"6e", x"6c", x"6c", x"6d", x"6c", x"6c", 
        x"6c", x"6c", x"6b", x"6c", x"6c", x"6b", x"70", x"6d", x"6c", x"6f", x"70", x"6e", x"6e", x"6c", x"6c", 
        x"6a", x"6b", x"6c", x"6c", x"6e", x"70", x"6e", x"6d", x"6e", x"6e", x"6e", x"6b", x"6a", x"69", x"69", 
        x"6d", x"6d", x"6c", x"6d", x"6c", x"6c", x"6e", x"6f", x"6f", x"6e", x"6c", x"6c", x"6d", x"6c", x"6c", 
        x"6d", x"6d", x"6b", x"6b", x"6e", x"6e", x"6d", x"6d", x"6d", x"6d", x"6b", x"6a", x"6c", x"6d", x"6c", 
        x"6c", x"6c", x"6b", x"69", x"6b", x"6d", x"6d", x"6b", x"6b", x"6e", x"6e", x"6e", x"6c", x"6c", x"6d", 
        x"6e", x"6e", x"6f", x"6f", x"6f", x"6f", x"70", x"70", x"70", x"71", x"71", x"6f", x"72", x"72", x"6f", 
        x"6b", x"69", x"6c", x"6f", x"6e", x"6c", x"6b", x"6c", x"6d", x"6f", x"6d", x"6e", x"6f", x"6d", x"6d", 
        x"6e", x"6d", x"6e", x"6e", x"6e", x"6c", x"6c", x"6c", x"6c", x"6c", x"6a", x"6b", x"6a", x"6a", x"6d", 
        x"6c", x"69", x"6b", x"6c", x"6e", x"6d", x"6c", x"6d", x"6c", x"6c", x"6c", x"6b", x"6c", x"6b", x"6a", 
        x"68", x"6b", x"6b", x"6b", x"6c", x"6c", x"6c", x"6a", x"6c", x"6d", x"6c", x"6c", x"6c", x"6b", x"6b", 
        x"6c", x"6d", x"6e", x"6c", x"6a", x"6b", x"6a", x"6a", x"6c", x"6b", x"6d", x"6d", x"6c", x"69", x"6b", 
        x"6d", x"6a", x"67", x"6b", x"6c", x"6c", x"6d", x"6e", x"6e", x"6b", x"6a", x"6d", x"6a", x"69", x"6a", 
        x"6a", x"69", x"69", x"69", x"6b", x"6b", x"6a", x"6b", x"6a", x"69", x"69", x"68", x"69", x"68", x"66", 
        x"66", x"67", x"69", x"68", x"67", x"67", x"6a", x"6a", x"69", x"69", x"68", x"6a", x"6b", x"69", x"6b", 
        x"68", x"6a", x"69", x"6a", x"67", x"66", x"68", x"68", x"68", x"68", x"67", x"66", x"67", x"69", x"6a", 
        x"69", x"68", x"67", x"67", x"67", x"67", x"67", x"66", x"66", x"66", x"64", x"66", x"64", x"64", x"66", 
        x"67", x"65", x"64", x"67", x"6a", x"6a", x"67", x"66", x"66", x"66", x"65", x"65", x"66", x"67", x"68", 
        x"68", x"67", x"65", x"65", x"67", x"64", x"66", x"67", x"64", x"65", x"65", x"63", x"64", x"64", x"64", 
        x"65", x"68", x"67", x"64", x"64", x"65", x"65", x"66", x"63", x"63", x"64", x"68", x"67", x"67", x"66", 
        x"64", x"66", x"65", x"64", x"64", x"64", x"64", x"64", x"64", x"65", x"65", x"64", x"64", x"64", x"64", 
        x"65", x"64", x"65", x"65", x"65", x"65", x"64", x"63", x"65", x"66", x"66", x"65", x"64", x"65", x"64", 
        x"64", x"64", x"64", x"64", x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"63", x"63", x"61", x"61", x"62", x"62", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"61", 
        x"61", x"62", x"62", x"62", x"62", x"62", x"61", x"60", x"61", x"61", x"61", x"60", x"60", x"60", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5f", 
        x"69", x"65", x"63", x"65", x"66", x"65", x"65", x"65", x"65", x"64", x"63", x"63", x"63", x"63", x"64", 
        x"64", x"63", x"62", x"61", x"61", x"61", x"61", x"62", x"64", x"65", x"63", x"61", x"61", x"61", x"63", 
        x"63", x"64", x"65", x"66", x"66", x"66", x"65", x"65", x"65", x"65", x"65", x"65", x"64", x"63", x"62", 
        x"62", x"62", x"63", x"64", x"66", x"6a", x"66", x"61", x"62", x"65", x"65", x"65", x"66", x"68", x"67", 
        x"64", x"61", x"62", x"62", x"63", x"65", x"64", x"63", x"63", x"64", x"65", x"65", x"64", x"65", x"65", 
        x"66", x"65", x"65", x"64", x"66", x"64", x"63", x"64", x"66", x"65", x"62", x"62", x"65", x"67", x"65", 
        x"65", x"66", x"65", x"66", x"66", x"66", x"66", x"64", x"63", x"65", x"65", x"65", x"67", x"65", x"65", 
        x"66", x"65", x"62", x"63", x"64", x"65", x"65", x"66", x"68", x"69", x"64", x"65", x"68", x"68", x"67", 
        x"66", x"66", x"66", x"68", x"68", x"68", x"6a", x"6b", x"68", x"67", x"66", x"67", x"6b", x"6a", x"68", 
        x"68", x"68", x"68", x"68", x"6b", x"6a", x"66", x"69", x"6a", x"69", x"67", x"67", x"65", x"67", x"6a", 
        x"6a", x"69", x"68", x"67", x"6b", x"69", x"64", x"69", x"69", x"69", x"6b", x"6b", x"67", x"6a", x"69", 
        x"69", x"6b", x"6b", x"69", x"67", x"68", x"6b", x"6a", x"6b", x"6c", x"69", x"69", x"6b", x"6a", x"66", 
        x"62", x"76", x"af", x"c8", x"a0", x"8d", x"b4", x"d0", x"cd", x"ca", x"cb", x"cc", x"cc", x"cb", x"cc", 
        x"cb", x"ca", x"cd", x"cc", x"ca", x"ca", x"cd", x"c9", x"cc", x"cd", x"cd", x"d0", x"d1", x"cc", x"a7", 
        x"69", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5a", x"5d", x"5f", 
        x"5d", x"5c", x"5e", x"61", x"5e", x"5c", x"5b", x"5b", x"5b", x"6e", x"97", x"bd", x"da", x"e9", x"e3", 
        x"c0", x"8f", x"6b", x"66", x"69", x"6e", x"73", x"71", x"6f", x"72", x"6f", x"6e", x"6d", x"6c", x"6e", 
        x"6c", x"69", x"6c", x"6f", x"6d", x"6d", x"6f", x"70", x"6f", x"6f", x"6e", x"6c", x"6e", x"6f", x"6f", 
        x"6d", x"6c", x"6d", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6d", x"6d", x"6d", x"6f", x"70", x"6c", 
        x"6c", x"6f", x"70", x"6e", x"6c", x"6b", x"6f", x"6f", x"71", x"6f", x"6f", x"6d", x"6e", x"6f", x"6b", 
        x"6b", x"6e", x"6f", x"6e", x"6d", x"6e", x"70", x"6e", x"6d", x"6c", x"6d", x"6d", x"6e", x"6e", x"6c", 
        x"6d", x"6d", x"6e", x"6f", x"6f", x"6e", x"6d", x"6e", x"70", x"6e", x"6c", x"6c", x"6b", x"6c", x"6d", 
        x"6f", x"6e", x"6b", x"6c", x"6a", x"6a", x"70", x"6c", x"6a", x"6f", x"70", x"6d", x"6e", x"6c", x"6f", 
        x"6e", x"6e", x"6c", x"6b", x"6f", x"70", x"70", x"6e", x"6d", x"6e", x"6e", x"6c", x"6c", x"6d", x"6d", 
        x"6f", x"6c", x"6a", x"6c", x"6e", x"6c", x"6d", x"72", x"70", x"6c", x"6d", x"6f", x"6f", x"6e", x"6e", 
        x"6d", x"6b", x"67", x"68", x"6e", x"6e", x"6c", x"6d", x"6c", x"6e", x"6c", x"6c", x"6b", x"6a", x"6a", 
        x"6b", x"6c", x"6c", x"6b", x"6e", x"6f", x"70", x"6e", x"6d", x"6e", x"6d", x"6f", x"6f", x"6e", x"6f", 
        x"6f", x"6f", x"6f", x"6f", x"6e", x"6f", x"6f", x"6f", x"6f", x"70", x"6f", x"6e", x"6d", x"70", x"6f", 
        x"6e", x"6e", x"6d", x"6e", x"6d", x"6d", x"6c", x"6b", x"6d", x"6e", x"6b", x"6c", x"6d", x"6c", x"6d", 
        x"6f", x"6e", x"6c", x"6d", x"6d", x"6c", x"6c", x"6d", x"6e", x"6d", x"6a", x"69", x"69", x"6b", x"6b", 
        x"6a", x"69", x"6b", x"69", x"6d", x"6e", x"6c", x"6c", x"6a", x"6c", x"6b", x"6b", x"6c", x"6b", x"6a", 
        x"67", x"6a", x"6d", x"6b", x"6a", x"6c", x"6a", x"69", x"6c", x"6c", x"69", x"6c", x"6c", x"6a", x"6b", 
        x"6d", x"6d", x"70", x"6e", x"6c", x"6d", x"6e", x"6f", x"6f", x"6c", x"6c", x"6b", x"6a", x"68", x"6b", 
        x"6d", x"6b", x"6a", x"6d", x"6c", x"6d", x"6f", x"6f", x"6f", x"6c", x"6c", x"6c", x"69", x"69", x"6a", 
        x"6b", x"69", x"6a", x"68", x"6a", x"6b", x"68", x"6b", x"6b", x"68", x"68", x"68", x"69", x"6a", x"69", 
        x"69", x"69", x"6a", x"69", x"67", x"67", x"69", x"67", x"68", x"6a", x"68", x"67", x"6b", x"66", x"6a", 
        x"66", x"68", x"69", x"6b", x"67", x"63", x"66", x"68", x"6a", x"6a", x"68", x"68", x"69", x"6a", x"69", 
        x"68", x"65", x"65", x"67", x"66", x"67", x"67", x"65", x"66", x"67", x"65", x"68", x"67", x"67", x"69", 
        x"68", x"66", x"66", x"67", x"69", x"66", x"66", x"68", x"68", x"67", x"66", x"66", x"66", x"67", x"67", 
        x"67", x"66", x"66", x"65", x"66", x"63", x"65", x"68", x"64", x"65", x"65", x"63", x"65", x"65", x"64", 
        x"64", x"66", x"68", x"68", x"66", x"66", x"65", x"67", x"64", x"64", x"67", x"69", x"67", x"67", x"65", 
        x"62", x"66", x"64", x"65", x"66", x"66", x"66", x"65", x"63", x"64", x"67", x"64", x"65", x"64", x"64", 
        x"67", x"64", x"64", x"63", x"63", x"63", x"64", x"64", x"64", x"64", x"65", x"66", x"65", x"66", x"63", 
        x"63", x"63", x"64", x"64", x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"64", x"63", x"61", x"61", x"62", x"62", x"61", x"60", x"61", x"61", x"61", x"61", x"60", x"60", x"60", 
        x"61", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"60", x"60", x"60", x"61", x"61", x"5f", 
        x"5f", x"5f", x"60", x"61", x"61", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5f", 
        x"67", x"65", x"62", x"65", x"64", x"64", x"64", x"64", x"65", x"63", x"62", x"63", x"63", x"63", x"63", 
        x"63", x"64", x"64", x"63", x"63", x"63", x"63", x"63", x"64", x"64", x"63", x"63", x"63", x"63", x"63", 
        x"63", x"62", x"63", x"65", x"67", x"66", x"64", x"63", x"63", x"64", x"64", x"63", x"64", x"64", x"63", 
        x"61", x"62", x"63", x"64", x"64", x"67", x"65", x"62", x"62", x"64", x"65", x"65", x"65", x"65", x"65", 
        x"63", x"62", x"63", x"64", x"65", x"65", x"65", x"65", x"65", x"65", x"64", x"64", x"65", x"66", x"65", 
        x"64", x"64", x"65", x"66", x"65", x"64", x"62", x"64", x"66", x"67", x"67", x"63", x"65", x"67", x"65", 
        x"66", x"67", x"65", x"65", x"65", x"66", x"67", x"66", x"65", x"67", x"67", x"66", x"66", x"65", x"64", 
        x"64", x"64", x"64", x"65", x"66", x"65", x"65", x"65", x"64", x"65", x"64", x"64", x"65", x"66", x"66", 
        x"66", x"67", x"67", x"68", x"69", x"69", x"69", x"68", x"63", x"64", x"65", x"64", x"66", x"66", x"65", 
        x"65", x"68", x"6a", x"68", x"6a", x"6a", x"67", x"6b", x"6c", x"69", x"68", x"69", x"67", x"67", x"6a", 
        x"6a", x"6b", x"6b", x"69", x"6a", x"69", x"67", x"6a", x"68", x"6a", x"6b", x"6a", x"69", x"6c", x"6a", 
        x"69", x"6a", x"6b", x"69", x"68", x"67", x"68", x"69", x"6a", x"6d", x"6a", x"67", x"6d", x"67", x"63", 
        x"8f", x"c0", x"c0", x"94", x"97", x"c5", x"d1", x"cd", x"ce", x"cc", x"cd", x"c9", x"cc", x"cb", x"cc", 
        x"cb", x"cb", x"cf", x"ce", x"cb", x"ca", x"cf", x"cc", x"ce", x"ce", x"ce", x"ce", x"d0", x"cd", x"a9", 
        x"6a", x"5e", x"5f", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5d", x"5c", 
        x"5e", x"61", x"60", x"5c", x"5e", x"5e", x"5f", x"5e", x"5d", x"5f", x"61", x"6f", x"8a", x"ad", x"ce", 
        x"e5", x"ea", x"c9", x"a0", x"7f", x"6a", x"64", x"67", x"71", x"75", x"71", x"6d", x"6f", x"71", x"6e", 
        x"6d", x"6f", x"6f", x"6d", x"6b", x"6c", x"6f", x"70", x"70", x"6f", x"71", x"70", x"6f", x"72", x"73", 
        x"72", x"71", x"70", x"70", x"6f", x"6e", x"6e", x"6e", x"6f", x"6f", x"6f", x"6d", x"6f", x"70", x"6e", 
        x"6e", x"6f", x"6e", x"6d", x"6e", x"6e", x"6f", x"6e", x"6f", x"70", x"70", x"6e", x"70", x"70", x"6d", 
        x"6e", x"6f", x"6e", x"6f", x"6e", x"6e", x"71", x"70", x"6d", x"6d", x"6d", x"6d", x"6c", x"6c", x"6a", 
        x"6b", x"6d", x"6d", x"6c", x"6c", x"6d", x"6e", x"6d", x"6c", x"6e", x"6d", x"6d", x"6e", x"6f", x"70", 
        x"6d", x"6e", x"6c", x"6c", x"6c", x"6e", x"73", x"6e", x"6d", x"6f", x"6f", x"6e", x"70", x"6e", x"6d", 
        x"6e", x"6f", x"6e", x"6e", x"71", x"71", x"71", x"70", x"6d", x"6d", x"6d", x"6c", x"6d", x"6d", x"6e", 
        x"6f", x"6e", x"6d", x"6e", x"6e", x"6c", x"6a", x"6e", x"6e", x"6c", x"6e", x"6f", x"6e", x"70", x"6f", 
        x"6e", x"6d", x"6b", x"6b", x"70", x"70", x"6e", x"6f", x"6d", x"6b", x"6a", x"6a", x"69", x"6b", x"6c", 
        x"6c", x"6e", x"70", x"6d", x"6b", x"6a", x"6b", x"6c", x"6d", x"6e", x"6e", x"70", x"70", x"6f", x"6e", 
        x"6d", x"6e", x"6f", x"71", x"70", x"6f", x"6d", x"6f", x"70", x"6f", x"70", x"70", x"6e", x"6f", x"6e", 
        x"6d", x"6e", x"6b", x"6c", x"6d", x"6f", x"6d", x"6b", x"6c", x"6b", x"6a", x"6d", x"6e", x"6d", x"6e", 
        x"6f", x"6d", x"6b", x"6c", x"6c", x"6d", x"6e", x"6d", x"6c", x"6c", x"6e", x"6d", x"6e", x"6f", x"6e", 
        x"6e", x"6e", x"6c", x"68", x"69", x"6b", x"69", x"6d", x"6c", x"6e", x"6d", x"6c", x"6c", x"6c", x"6c", 
        x"6b", x"6d", x"6e", x"6d", x"6b", x"6d", x"6c", x"6c", x"6d", x"6d", x"6a", x"6b", x"6e", x"6b", x"6b", 
        x"6c", x"6a", x"6d", x"6c", x"6b", x"6c", x"6c", x"6b", x"6c", x"6c", x"6b", x"69", x"68", x"69", x"6c", 
        x"6b", x"6b", x"6c", x"6d", x"6c", x"6c", x"6e", x"6c", x"6d", x"6d", x"6c", x"6b", x"69", x"69", x"6b", 
        x"6c", x"6b", x"6b", x"6a", x"6b", x"6a", x"68", x"69", x"6a", x"6a", x"6b", x"6b", x"6a", x"69", x"6a", 
        x"6b", x"6b", x"6a", x"6a", x"69", x"6a", x"6d", x"6c", x"6c", x"6c", x"69", x"66", x"6a", x"68", x"6a", 
        x"67", x"69", x"6a", x"6c", x"68", x"65", x"66", x"6a", x"6a", x"69", x"69", x"68", x"69", x"68", x"69", 
        x"68", x"64", x"65", x"66", x"67", x"6b", x"69", x"67", x"67", x"69", x"68", x"69", x"69", x"69", x"6a", 
        x"68", x"68", x"69", x"68", x"68", x"66", x"67", x"69", x"68", x"66", x"67", x"66", x"65", x"67", x"66", 
        x"65", x"67", x"66", x"66", x"67", x"65", x"65", x"67", x"64", x"65", x"66", x"65", x"66", x"66", x"64", 
        x"63", x"65", x"66", x"66", x"65", x"65", x"64", x"66", x"64", x"65", x"67", x"68", x"66", x"64", x"63", 
        x"63", x"65", x"64", x"64", x"66", x"67", x"66", x"66", x"63", x"64", x"68", x"64", x"66", x"66", x"64", 
        x"67", x"64", x"63", x"64", x"65", x"65", x"65", x"67", x"66", x"63", x"65", x"65", x"65", x"65", x"63", 
        x"63", x"63", x"62", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"63", x"62", x"62", x"61", x"62", x"62", x"61", x"60", x"60", x"61", x"61", x"61", x"61", x"60", x"60", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"5f", x"60", x"61", x"61", x"60", x"5f", 
        x"60", x"60", x"61", x"61", x"60", x"61", x"61", x"60", x"60", x"60", x"60", x"60", x"60", x"5f", x"5f", 
        x"62", x"63", x"62", x"63", x"62", x"63", x"63", x"64", x"66", x"63", x"62", x"64", x"62", x"63", x"64", 
        x"64", x"65", x"66", x"65", x"64", x"65", x"64", x"64", x"64", x"65", x"64", x"64", x"64", x"65", x"65", 
        x"65", x"62", x"61", x"65", x"66", x"64", x"64", x"63", x"64", x"65", x"64", x"63", x"64", x"64", x"63", 
        x"62", x"63", x"64", x"64", x"64", x"64", x"63", x"63", x"63", x"63", x"65", x"66", x"66", x"65", x"64", 
        x"64", x"64", x"65", x"65", x"63", x"62", x"62", x"63", x"66", x"66", x"65", x"64", x"66", x"64", x"63", 
        x"63", x"64", x"67", x"68", x"64", x"65", x"62", x"64", x"64", x"66", x"68", x"65", x"66", x"66", x"66", 
        x"66", x"67", x"66", x"65", x"67", x"66", x"67", x"67", x"66", x"67", x"66", x"67", x"65", x"66", x"66", 
        x"65", x"65", x"68", x"69", x"69", x"67", x"68", x"69", x"66", x"67", x"66", x"65", x"64", x"65", x"66", 
        x"67", x"68", x"67", x"67", x"67", x"68", x"69", x"69", x"67", x"6a", x"69", x"65", x"66", x"66", x"66", 
        x"67", x"69", x"69", x"68", x"68", x"68", x"69", x"6a", x"6a", x"68", x"68", x"6a", x"6a", x"67", x"66", 
        x"67", x"67", x"6b", x"6a", x"6a", x"6b", x"6a", x"6a", x"67", x"6b", x"69", x"69", x"69", x"6c", x"6a", 
        x"6d", x"6c", x"6a", x"6a", x"6b", x"68", x"6a", x"6c", x"69", x"6d", x"6c", x"69", x"67", x"72", x"9c", 
        x"c4", x"b3", x"8e", x"a8", x"cc", x"d2", x"ca", x"cc", x"cc", x"cc", x"cd", x"cd", x"cd", x"ce", x"ce", 
        x"cd", x"cd", x"ce", x"cf", x"cd", x"cc", x"cf", x"cc", x"ce", x"ce", x"ce", x"cd", x"cf", x"ce", x"ab", 
        x"69", x"5d", x"5f", x"5c", x"5d", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5d", x"5e", x"5d", x"60", x"61", x"5e", x"5f", x"60", x"5d", x"60", x"6b", x"82", 
        x"a3", x"c6", x"df", x"e4", x"d4", x"ad", x"89", x"70", x"6a", x"6d", x"71", x"70", x"6e", x"72", x"71", 
        x"6d", x"6e", x"71", x"71", x"6d", x"6e", x"6f", x"6f", x"73", x"71", x"71", x"70", x"70", x"71", x"72", 
        x"72", x"71", x"6f", x"6f", x"6e", x"6e", x"6f", x"70", x"71", x"70", x"6f", x"6f", x"6e", x"6f", x"6f", 
        x"6f", x"6e", x"6d", x"6d", x"6f", x"71", x"6f", x"6d", x"6d", x"6f", x"6d", x"6e", x"70", x"6f", x"6f", 
        x"71", x"71", x"6e", x"70", x"70", x"6f", x"71", x"70", x"70", x"6d", x"6e", x"6f", x"6d", x"6d", x"6e", 
        x"6c", x"6d", x"6e", x"6c", x"6b", x"6d", x"6f", x"6d", x"6d", x"72", x"71", x"6e", x"70", x"6e", x"6e", 
        x"6a", x"6d", x"6f", x"6e", x"6d", x"6f", x"70", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6f", 
        x"70", x"70", x"6e", x"6d", x"6f", x"71", x"6f", x"6e", x"6e", x"6e", x"6d", x"6d", x"6c", x"6c", x"6d", 
        x"6e", x"6f", x"6f", x"70", x"6f", x"6d", x"6b", x"6c", x"6c", x"6e", x"6e", x"6d", x"6b", x"6c", x"6f", 
        x"6d", x"6d", x"6d", x"6c", x"6f", x"6d", x"6c", x"6f", x"6e", x"6a", x"6c", x"6b", x"69", x"6d", x"6d", 
        x"6c", x"6e", x"70", x"6c", x"6c", x"6d", x"6b", x"6d", x"6e", x"6d", x"6e", x"6e", x"6c", x"6e", x"6e", 
        x"6c", x"6d", x"6c", x"6e", x"6f", x"6e", x"6a", x"6d", x"6f", x"6d", x"6e", x"6e", x"6f", x"6f", x"6d", 
        x"6d", x"6e", x"6c", x"6a", x"6c", x"6f", x"6b", x"6d", x"6d", x"6c", x"6c", x"6e", x"6e", x"6c", x"6c", 
        x"6e", x"6d", x"6c", x"6b", x"6b", x"6c", x"6d", x"6c", x"69", x"69", x"6e", x"6f", x"70", x"70", x"70", 
        x"70", x"6f", x"6c", x"6d", x"6b", x"6c", x"6b", x"6d", x"6d", x"6c", x"6d", x"6d", x"6e", x"6d", x"6c", 
        x"6c", x"6b", x"6b", x"6b", x"6b", x"6c", x"6d", x"6e", x"6c", x"6e", x"6d", x"6b", x"6f", x"6c", x"69", 
        x"6d", x"6d", x"6c", x"6d", x"6d", x"6d", x"6a", x"69", x"6b", x"6e", x"6d", x"6c", x"6b", x"6d", x"6c", 
        x"6a", x"6b", x"6d", x"6d", x"6c", x"6c", x"6d", x"6c", x"6c", x"70", x"6e", x"6c", x"6b", x"6b", x"6c", 
        x"6a", x"6c", x"6a", x"6a", x"6a", x"68", x"6a", x"6a", x"69", x"69", x"6a", x"6b", x"6b", x"6b", x"69", 
        x"69", x"6a", x"68", x"68", x"6b", x"6c", x"6b", x"6d", x"6b", x"6c", x"6a", x"68", x"69", x"69", x"68", 
        x"68", x"68", x"6a", x"68", x"66", x"68", x"68", x"6a", x"68", x"67", x"68", x"67", x"67", x"68", x"6a", 
        x"68", x"67", x"68", x"68", x"6a", x"6d", x"6a", x"68", x"69", x"6a", x"69", x"68", x"69", x"68", x"69", 
        x"67", x"67", x"69", x"67", x"68", x"68", x"67", x"67", x"67", x"67", x"67", x"65", x"64", x"68", x"65", 
        x"64", x"67", x"66", x"67", x"68", x"68", x"67", x"66", x"66", x"66", x"68", x"67", x"67", x"68", x"64", 
        x"65", x"66", x"64", x"65", x"65", x"65", x"67", x"68", x"67", x"66", x"66", x"67", x"66", x"63", x"63", 
        x"65", x"65", x"66", x"65", x"66", x"67", x"65", x"65", x"63", x"63", x"69", x"64", x"66", x"66", x"64", 
        x"67", x"64", x"63", x"65", x"66", x"65", x"65", x"65", x"65", x"65", x"65", x"64", x"64", x"64", x"65", 
        x"65", x"65", x"63", x"63", x"64", x"63", x"61", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"61", x"61", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"61", x"62", x"62", x"62", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"60", x"5f", x"5f", x"61", x"62", x"61", x"61", x"60", 
        x"61", x"61", x"61", x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"60", 
        x"63", x"64", x"63", x"65", x"63", x"64", x"64", x"64", x"66", x"64", x"63", x"64", x"63", x"64", x"64", 
        x"65", x"65", x"65", x"64", x"64", x"65", x"64", x"64", x"64", x"64", x"63", x"63", x"64", x"64", x"65", 
        x"65", x"63", x"61", x"64", x"65", x"63", x"64", x"64", x"65", x"65", x"63", x"62", x"65", x"64", x"64", 
        x"65", x"64", x"63", x"64", x"66", x"65", x"64", x"64", x"63", x"64", x"64", x"64", x"66", x"66", x"65", 
        x"65", x"65", x"65", x"64", x"63", x"63", x"61", x"61", x"63", x"65", x"65", x"65", x"64", x"62", x"61", 
        x"63", x"65", x"65", x"65", x"65", x"66", x"64", x"64", x"63", x"64", x"65", x"66", x"66", x"65", x"68", 
        x"67", x"67", x"68", x"68", x"69", x"66", x"66", x"66", x"65", x"67", x"68", x"68", x"67", x"69", x"69", 
        x"68", x"67", x"68", x"69", x"6a", x"68", x"69", x"68", x"67", x"68", x"65", x"66", x"67", x"68", x"68", 
        x"66", x"65", x"69", x"68", x"66", x"68", x"6a", x"6b", x"6a", x"6c", x"6a", x"68", x"69", x"69", x"69", 
        x"6a", x"69", x"67", x"67", x"67", x"67", x"68", x"69", x"69", x"68", x"67", x"69", x"6a", x"68", x"67", 
        x"66", x"65", x"69", x"68", x"69", x"6b", x"6a", x"6b", x"69", x"6a", x"69", x"6a", x"69", x"69", x"6a", 
        x"6b", x"6e", x"6e", x"6e", x"6e", x"6b", x"68", x"69", x"69", x"6d", x"6a", x"61", x"7d", x"b6", x"ce", 
        x"9d", x"93", x"bb", x"d1", x"d1", x"ce", x"cb", x"cc", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"ce", 
        x"cd", x"cd", x"cd", x"ce", x"cd", x"cb", x"cf", x"cd", x"ce", x"cf", x"cf", x"ce", x"cf", x"ce", x"ac", 
        x"6a", x"5d", x"5f", x"5c", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5b", x"5f", x"60", x"5b", x"5b", x"5f", x"5e", x"5c", x"5a", x"5c", 
        x"63", x"77", x"97", x"bb", x"dd", x"e9", x"df", x"c0", x"92", x"73", x"62", x"64", x"6d", x"71", x"71", 
        x"71", x"71", x"72", x"74", x"70", x"6f", x"6f", x"70", x"74", x"74", x"6e", x"6d", x"6c", x"6d", x"6f", 
        x"6f", x"6f", x"6f", x"70", x"70", x"70", x"70", x"71", x"72", x"6f", x"6d", x"6f", x"6e", x"6c", x"6d", 
        x"6f", x"70", x"6e", x"6d", x"6f", x"70", x"6e", x"6d", x"6e", x"6e", x"6d", x"6e", x"70", x"6e", x"6e", 
        x"6f", x"6e", x"6b", x"6d", x"6e", x"6e", x"6f", x"6c", x"6d", x"6c", x"6f", x"71", x"70", x"71", x"70", 
        x"6f", x"6f", x"6f", x"6c", x"6c", x"6e", x"6f", x"6e", x"6f", x"72", x"71", x"6e", x"70", x"6d", x"6d", 
        x"6c", x"6d", x"70", x"72", x"70", x"6f", x"70", x"6e", x"6e", x"6f", x"6e", x"6d", x"6d", x"6f", x"6e", 
        x"6e", x"6e", x"6d", x"6d", x"6f", x"71", x"6e", x"6d", x"6f", x"70", x"6f", x"6d", x"6b", x"6c", x"6f", 
        x"6e", x"6e", x"6e", x"6f", x"70", x"6f", x"6c", x"6c", x"6d", x"6e", x"6f", x"6e", x"6d", x"6a", x"70", 
        x"70", x"6f", x"6d", x"6b", x"6e", x"6d", x"6c", x"6f", x"6e", x"6b", x"6c", x"6c", x"6c", x"6f", x"6d", 
        x"6d", x"6c", x"6d", x"6d", x"6e", x"6f", x"6c", x"6d", x"6e", x"6d", x"6d", x"6e", x"6c", x"6e", x"6f", 
        x"6f", x"70", x"6d", x"6d", x"6f", x"6f", x"6d", x"6f", x"70", x"6d", x"6e", x"6c", x"6e", x"70", x"6e", 
        x"6e", x"6e", x"6d", x"6b", x"6d", x"6f", x"6c", x"6d", x"6f", x"70", x"70", x"70", x"6d", x"6a", x"6a", 
        x"6d", x"6e", x"6e", x"6e", x"6d", x"6d", x"6e", x"6e", x"6d", x"6c", x"6c", x"6e", x"6e", x"6e", x"6f", 
        x"70", x"70", x"6d", x"6f", x"6d", x"6f", x"6c", x"6c", x"6a", x"6a", x"6c", x"6c", x"6e", x"6d", x"6d", 
        x"6c", x"6a", x"6a", x"6b", x"6b", x"6b", x"6b", x"6b", x"68", x"6a", x"6b", x"6b", x"70", x"6d", x"69", 
        x"6d", x"6d", x"6c", x"6c", x"6d", x"6e", x"6d", x"6c", x"6d", x"6d", x"6b", x"6c", x"6e", x"6e", x"6a", 
        x"6d", x"6e", x"6e", x"6d", x"6d", x"6e", x"70", x"6c", x"6a", x"6e", x"6c", x"6c", x"6b", x"6b", x"6c", 
        x"6a", x"6a", x"69", x"68", x"69", x"69", x"6a", x"6a", x"69", x"69", x"68", x"69", x"6a", x"6c", x"6c", 
        x"6a", x"69", x"69", x"6a", x"6c", x"6b", x"68", x"6b", x"6b", x"6d", x"6d", x"6a", x"6a", x"66", x"68", 
        x"6a", x"69", x"67", x"66", x"68", x"69", x"68", x"6a", x"69", x"67", x"67", x"66", x"67", x"69", x"68", 
        x"65", x"65", x"67", x"69", x"6a", x"6a", x"69", x"69", x"69", x"69", x"68", x"66", x"68", x"6a", x"67", 
        x"66", x"67", x"67", x"65", x"69", x"67", x"65", x"67", x"69", x"69", x"68", x"66", x"66", x"66", x"63", 
        x"64", x"67", x"68", x"68", x"67", x"68", x"69", x"68", x"68", x"67", x"68", x"67", x"67", x"68", x"66", 
        x"66", x"67", x"66", x"66", x"64", x"65", x"68", x"6a", x"68", x"66", x"67", x"67", x"68", x"67", x"67", 
        x"66", x"65", x"67", x"66", x"67", x"67", x"64", x"65", x"65", x"66", x"69", x"64", x"65", x"64", x"64", 
        x"67", x"66", x"66", x"65", x"65", x"68", x"69", x"65", x"64", x"67", x"66", x"66", x"65", x"65", x"64", 
        x"64", x"64", x"63", x"63", x"65", x"63", x"63", x"64", x"63", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"60", x"60", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"60", x"60", x"62", x"62", x"61", x"61", 
        x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"60", x"5f", x"5f", x"5f", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", 
        x"65", x"65", x"64", x"66", x"65", x"65", x"65", x"65", x"65", x"64", x"64", x"64", x"64", x"65", x"65", 
        x"65", x"66", x"66", x"66", x"66", x"65", x"64", x"64", x"63", x"63", x"63", x"63", x"64", x"63", x"63", 
        x"65", x"63", x"61", x"63", x"65", x"65", x"63", x"64", x"66", x"66", x"63", x"62", x"65", x"63", x"64", 
        x"65", x"64", x"63", x"64", x"66", x"66", x"65", x"65", x"64", x"64", x"64", x"64", x"64", x"64", x"64", 
        x"65", x"66", x"66", x"64", x"64", x"65", x"63", x"62", x"63", x"65", x"67", x"66", x"64", x"63", x"63", 
        x"63", x"63", x"63", x"63", x"65", x"66", x"65", x"64", x"63", x"64", x"64", x"67", x"67", x"66", x"67", 
        x"67", x"67", x"69", x"65", x"65", x"63", x"64", x"65", x"67", x"6a", x"6a", x"6a", x"6a", x"6a", x"69", 
        x"66", x"63", x"63", x"67", x"68", x"67", x"67", x"66", x"66", x"67", x"64", x"66", x"68", x"69", x"69", 
        x"67", x"66", x"67", x"66", x"65", x"67", x"69", x"69", x"69", x"6b", x"69", x"68", x"69", x"69", x"69", 
        x"69", x"69", x"69", x"69", x"69", x"68", x"69", x"69", x"69", x"6a", x"69", x"6b", x"6c", x"6c", x"6b", 
        x"69", x"68", x"6b", x"69", x"68", x"68", x"67", x"68", x"69", x"69", x"69", x"69", x"69", x"6a", x"6a", 
        x"68", x"6c", x"6e", x"6b", x"6a", x"6d", x"6d", x"6d", x"6e", x"66", x"62", x"8f", x"c8", x"b9", x"93", 
        x"a6", x"c8", x"d1", x"ca", x"ca", x"cd", x"ca", x"cc", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"cd", 
        x"cd", x"cd", x"cd", x"ce", x"cc", x"cb", x"cf", x"cd", x"d0", x"d0", x"d0", x"cf", x"cf", x"cf", x"af", 
        x"6c", x"5d", x"5f", x"5c", x"5c", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5c", x"5c", x"5e", x"5d", x"5b", x"5c", x"61", 
        x"5f", x"5c", x"62", x"70", x"89", x"b7", x"db", x"f0", x"e6", x"cf", x"ac", x"7f", x"69", x"69", x"6c", 
        x"6c", x"73", x"78", x"78", x"72", x"72", x"72", x"70", x"71", x"6f", x"6e", x"6c", x"6d", x"6e", x"71", 
        x"72", x"71", x"71", x"71", x"71", x"71", x"71", x"71", x"71", x"70", x"70", x"71", x"6f", x"6c", x"6b", 
        x"6d", x"6e", x"6e", x"6e", x"6f", x"6f", x"6d", x"6e", x"6f", x"6e", x"6e", x"6f", x"70", x"6f", x"6e", 
        x"6e", x"6e", x"6e", x"6f", x"6f", x"6e", x"6f", x"6e", x"70", x"6f", x"70", x"71", x"6f", x"6f", x"6f", 
        x"6d", x"6f", x"6d", x"6b", x"6c", x"6e", x"6c", x"6d", x"71", x"71", x"6f", x"6e", x"70", x"6f", x"6e", 
        x"6e", x"6b", x"6c", x"6e", x"6e", x"6e", x"6f", x"70", x"71", x"70", x"6f", x"6c", x"6c", x"6d", x"6c", 
        x"6d", x"70", x"70", x"6f", x"6e", x"6e", x"6f", x"6f", x"6e", x"6e", x"6e", x"6e", x"6e", x"6d", x"6e", 
        x"6f", x"70", x"70", x"6f", x"6f", x"6d", x"6b", x"6d", x"6e", x"6e", x"6e", x"6f", x"70", x"6d", x"6e", 
        x"6e", x"70", x"6f", x"6d", x"6d", x"6d", x"6e", x"6f", x"6f", x"6d", x"6d", x"6d", x"6e", x"6f", x"6d", 
        x"6e", x"6c", x"6b", x"6e", x"6f", x"6f", x"6d", x"6d", x"6f", x"6e", x"6d", x"6c", x"6b", x"6c", x"6e", 
        x"6e", x"6e", x"6b", x"6b", x"6d", x"6f", x"6f", x"70", x"6f", x"6e", x"6e", x"6d", x"70", x"70", x"6d", 
        x"6c", x"6e", x"6e", x"6c", x"6c", x"6c", x"6b", x"6c", x"6e", x"6f", x"6e", x"6d", x"6b", x"6a", x"6d", 
        x"6f", x"6e", x"6c", x"6d", x"6c", x"6c", x"6c", x"6d", x"6d", x"6c", x"6c", x"6e", x"6d", x"6c", x"6c", 
        x"6e", x"71", x"6d", x"6d", x"6d", x"6e", x"6d", x"6e", x"6d", x"6c", x"6c", x"6b", x"6e", x"6d", x"6c", 
        x"6b", x"6e", x"6f", x"6e", x"6d", x"6c", x"6c", x"6b", x"6c", x"6f", x"6e", x"6d", x"6f", x"6e", x"6c", 
        x"6e", x"6e", x"6c", x"6c", x"6d", x"6f", x"6e", x"6c", x"6b", x"6d", x"6c", x"6c", x"6c", x"6d", x"6a", 
        x"6f", x"6f", x"6e", x"6d", x"6e", x"6f", x"71", x"6d", x"6b", x"6d", x"6d", x"6d", x"6d", x"6b", x"6d", 
        x"6b", x"6d", x"6c", x"6a", x"6c", x"6c", x"6c", x"6b", x"6b", x"6a", x"68", x"68", x"69", x"6b", x"6c", 
        x"6b", x"6a", x"6a", x"6b", x"6b", x"6a", x"6a", x"6d", x"6c", x"6c", x"6b", x"68", x"68", x"66", x"69", 
        x"6d", x"6d", x"6a", x"6a", x"6c", x"6b", x"6b", x"6d", x"6c", x"6a", x"69", x"68", x"68", x"68", x"68", 
        x"67", x"67", x"67", x"68", x"68", x"68", x"67", x"68", x"69", x"6a", x"6a", x"68", x"68", x"6c", x"68", 
        x"67", x"6b", x"6a", x"67", x"66", x"67", x"68", x"68", x"68", x"68", x"69", x"68", x"68", x"67", x"63", 
        x"66", x"66", x"68", x"67", x"65", x"66", x"66", x"66", x"66", x"65", x"66", x"67", x"67", x"68", x"67", 
        x"66", x"67", x"67", x"67", x"66", x"66", x"69", x"69", x"68", x"66", x"67", x"66", x"67", x"6a", x"69", 
        x"66", x"65", x"65", x"65", x"69", x"6a", x"66", x"66", x"64", x"65", x"67", x"65", x"67", x"64", x"64", 
        x"65", x"65", x"67", x"64", x"65", x"68", x"6a", x"66", x"65", x"66", x"66", x"66", x"66", x"65", x"64", 
        x"63", x"64", x"63", x"64", x"65", x"64", x"64", x"65", x"63", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"61", x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"62", x"61", x"61", x"60", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", x"61", x"62", x"61", x"61", x"61", x"61", x"60", 
        x"60", x"60", x"60", x"60", x"60", x"5f", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", 
        x"65", x"65", x"65", x"65", x"65", x"65", x"65", x"65", x"65", x"65", x"64", x"64", x"65", x"65", x"63", 
        x"62", x"63", x"65", x"65", x"64", x"62", x"62", x"64", x"64", x"65", x"64", x"64", x"65", x"64", x"63", 
        x"65", x"64", x"61", x"63", x"65", x"64", x"63", x"64", x"67", x"67", x"63", x"62", x"65", x"64", x"63", 
        x"62", x"63", x"63", x"64", x"65", x"64", x"65", x"65", x"65", x"65", x"64", x"65", x"64", x"63", x"64", 
        x"64", x"66", x"66", x"65", x"64", x"64", x"62", x"61", x"62", x"64", x"64", x"64", x"63", x"64", x"64", 
        x"63", x"62", x"65", x"67", x"65", x"64", x"65", x"64", x"64", x"64", x"64", x"67", x"68", x"66", x"66", 
        x"66", x"68", x"69", x"65", x"66", x"65", x"66", x"67", x"67", x"68", x"67", x"67", x"68", x"69", x"69", 
        x"68", x"66", x"66", x"69", x"6a", x"6a", x"69", x"67", x"68", x"69", x"6a", x"6a", x"69", x"68", x"67", 
        x"67", x"66", x"68", x"67", x"67", x"69", x"6a", x"6a", x"69", x"6a", x"68", x"66", x"68", x"67", x"67", 
        x"66", x"67", x"68", x"69", x"69", x"6a", x"6a", x"6b", x"6a", x"68", x"67", x"67", x"69", x"6a", x"69", 
        x"68", x"68", x"6b", x"69", x"69", x"69", x"68", x"68", x"68", x"6a", x"6a", x"68", x"6a", x"6d", x"6c", 
        x"6d", x"6d", x"6b", x"69", x"66", x"6a", x"6f", x"6f", x"67", x"72", x"9c", x"c8", x"ab", x"8f", x"ac", 
        x"cc", x"cf", x"c5", x"ce", x"d1", x"ca", x"cb", x"cc", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"cd", 
        x"cd", x"cd", x"cd", x"ce", x"cc", x"ca", x"ce", x"ce", x"d0", x"d1", x"d0", x"cf", x"cf", x"cf", x"af", 
        x"6d", x"5d", x"5f", x"5d", x"5c", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5c", x"5e", x"5f", x"5e", x"5e", x"5f", x"60", x"60", x"5d", x"5c", x"60", 
        x"61", x"67", x"78", x"8c", x"a5", x"c6", x"df", x"f0", x"f6", x"f6", x"ec", x"d7", x"b3", x"87", x"6a", 
        x"65", x"6b", x"72", x"71", x"6e", x"70", x"71", x"6c", x"6d", x"70", x"71", x"70", x"6f", x"70", x"70", 
        x"70", x"6e", x"70", x"72", x"72", x"72", x"72", x"71", x"71", x"71", x"72", x"71", x"70", x"6f", x"6f", 
        x"6d", x"6d", x"6e", x"6e", x"6f", x"6e", x"6c", x"6e", x"70", x"6f", x"6f", x"70", x"70", x"70", x"6e", 
        x"6e", x"6e", x"71", x"71", x"6f", x"6d", x"6e", x"72", x"71", x"6d", x"6f", x"6f", x"6e", x"70", x"70", 
        x"6f", x"71", x"71", x"70", x"71", x"72", x"6f", x"6f", x"74", x"71", x"6d", x"6c", x"6e", x"6e", x"6d", 
        x"6d", x"6d", x"6d", x"6e", x"6f", x"6d", x"6b", x"6e", x"70", x"70", x"6f", x"6e", x"6e", x"6e", x"70", 
        x"71", x"72", x"71", x"6e", x"6c", x"6b", x"6e", x"6f", x"6e", x"6c", x"6c", x"6e", x"70", x"70", x"6f", 
        x"6f", x"6f", x"6f", x"6f", x"6f", x"6d", x"6a", x"6c", x"6d", x"6d", x"6e", x"70", x"71", x"6f", x"6d", 
        x"6d", x"6f", x"70", x"6f", x"6d", x"6f", x"70", x"71", x"70", x"6f", x"6e", x"6f", x"6e", x"6d", x"6c", 
        x"70", x"6e", x"6c", x"6f", x"6f", x"6e", x"6d", x"6d", x"6f", x"70", x"6f", x"6e", x"6e", x"6e", x"6f", 
        x"70", x"70", x"6f", x"6d", x"6d", x"6d", x"6f", x"6f", x"6e", x"6e", x"6d", x"70", x"72", x"70", x"6c", 
        x"6c", x"6d", x"6d", x"6f", x"70", x"6f", x"6f", x"6f", x"6f", x"6f", x"6d", x"6c", x"6b", x"6b", x"6e", 
        x"70", x"6d", x"6c", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6f", x"6e", x"6b", x"69", 
        x"6c", x"6e", x"6a", x"6c", x"6f", x"70", x"6f", x"6d", x"6b", x"6d", x"6d", x"6c", x"6e", x"6d", x"6c", 
        x"6a", x"6d", x"6f", x"6f", x"6e", x"6e", x"6d", x"6d", x"6f", x"71", x"70", x"6e", x"6e", x"6d", x"6c", 
        x"6d", x"6d", x"6c", x"6c", x"6d", x"6e", x"6c", x"6b", x"6b", x"6e", x"6d", x"6d", x"6c", x"6d", x"6b", 
        x"6e", x"6e", x"6d", x"6d", x"6e", x"6f", x"70", x"6f", x"6e", x"6d", x"6e", x"6f", x"6d", x"6b", x"6d", 
        x"6b", x"6e", x"6f", x"6c", x"6d", x"6c", x"6a", x"69", x"6a", x"6b", x"6a", x"6b", x"6d", x"6c", x"68", 
        x"6a", x"6c", x"6b", x"6a", x"6b", x"6b", x"6a", x"6c", x"6a", x"6b", x"6a", x"69", x"6b", x"68", x"69", 
        x"6b", x"6d", x"6d", x"6d", x"6d", x"6c", x"6d", x"6e", x"6e", x"6c", x"6a", x"69", x"6a", x"6a", x"6b", 
        x"6b", x"6b", x"69", x"67", x"68", x"6a", x"6a", x"68", x"68", x"69", x"6a", x"68", x"67", x"6b", x"66", 
        x"66", x"6c", x"6a", x"67", x"68", x"6a", x"6c", x"6a", x"68", x"66", x"66", x"67", x"69", x"68", x"66", 
        x"68", x"66", x"67", x"68", x"66", x"66", x"65", x"65", x"65", x"65", x"66", x"67", x"67", x"67", x"67", 
        x"67", x"67", x"67", x"66", x"68", x"69", x"68", x"67", x"67", x"67", x"67", x"65", x"65", x"68", x"67", 
        x"66", x"66", x"65", x"65", x"69", x"6a", x"67", x"67", x"64", x"66", x"67", x"66", x"68", x"64", x"64", 
        x"64", x"65", x"68", x"67", x"66", x"66", x"65", x"65", x"64", x"64", x"65", x"65", x"65", x"65", x"64", 
        x"64", x"68", x"66", x"66", x"66", x"63", x"62", x"63", x"63", x"62", x"62", x"62", x"62", x"62", x"63", 
        x"62", x"62", x"61", x"61", x"61", x"60", x"60", x"61", x"62", x"61", x"61", x"62", x"61", x"60", x"60", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"61", x"62", x"62", x"61", x"61", x"61", x"62", x"60", 
        x"60", x"60", x"61", x"61", x"60", x"5f", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", 
        x"64", x"64", x"65", x"64", x"65", x"64", x"64", x"65", x"64", x"65", x"65", x"64", x"65", x"66", x"64", 
        x"64", x"66", x"68", x"69", x"67", x"64", x"62", x"65", x"65", x"65", x"65", x"65", x"65", x"64", x"63", 
        x"65", x"64", x"62", x"64", x"66", x"65", x"64", x"64", x"67", x"67", x"64", x"63", x"65", x"65", x"63", 
        x"61", x"62", x"65", x"65", x"64", x"64", x"65", x"66", x"66", x"65", x"66", x"66", x"66", x"65", x"65", 
        x"65", x"66", x"65", x"64", x"64", x"65", x"63", x"62", x"63", x"64", x"64", x"63", x"63", x"66", x"66", 
        x"63", x"62", x"65", x"69", x"64", x"63", x"65", x"65", x"65", x"64", x"65", x"66", x"68", x"67", x"65", 
        x"66", x"68", x"68", x"67", x"6a", x"69", x"6a", x"69", x"67", x"68", x"65", x"66", x"68", x"68", x"6a", 
        x"6b", x"6b", x"6b", x"6a", x"69", x"6a", x"68", x"67", x"69", x"69", x"6c", x"6a", x"68", x"66", x"66", 
        x"67", x"69", x"68", x"68", x"68", x"69", x"6a", x"69", x"67", x"6b", x"6a", x"67", x"68", x"67", x"67", 
        x"67", x"68", x"69", x"6a", x"6a", x"6b", x"6b", x"6b", x"6a", x"68", x"69", x"68", x"68", x"6a", x"6b", 
        x"69", x"67", x"6b", x"69", x"69", x"6a", x"69", x"6a", x"69", x"6b", x"6b", x"66", x"6a", x"6e", x"6b", 
        x"6a", x"6c", x"6c", x"6e", x"6f", x"6c", x"66", x"5e", x"7b", x"b7", x"ce", x"9e", x"92", x"bd", x"d4", 
        x"ce", x"cc", x"cd", x"cc", x"ca", x"c9", x"cb", x"cc", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"cd", 
        x"cd", x"cd", x"cd", x"ce", x"cc", x"cb", x"cf", x"ce", x"d0", x"d0", x"cf", x"ce", x"d0", x"cf", x"b0", 
        x"6e", x"5d", x"5f", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"5e", x"5f", x"61", x"5f", x"5c", x"5e", x"62", x"6c", x"83", 
        x"a3", x"c3", x"d9", x"e4", x"ec", x"ef", x"f1", x"f1", x"ee", x"eb", x"ea", x"ef", x"eb", x"e0", x"bd", 
        x"88", x"64", x"60", x"6e", x"6e", x"73", x"73", x"6f", x"71", x"75", x"75", x"74", x"72", x"72", x"72", 
        x"71", x"70", x"70", x"72", x"72", x"72", x"71", x"71", x"71", x"71", x"70", x"70", x"70", x"73", x"73", 
        x"70", x"6e", x"6e", x"6e", x"6f", x"6f", x"6d", x"6e", x"6f", x"70", x"71", x"70", x"70", x"70", x"6f", 
        x"6e", x"6e", x"72", x"71", x"6d", x"6a", x"6c", x"72", x"70", x"6c", x"6d", x"6e", x"6d", x"71", x"72", 
        x"6e", x"6e", x"70", x"6f", x"70", x"70", x"6d", x"6e", x"74", x"70", x"6c", x"6c", x"6e", x"71", x"6f", 
        x"6f", x"71", x"70", x"6f", x"71", x"6f", x"6c", x"6f", x"70", x"6f", x"6f", x"6f", x"6f", x"6e", x"70", 
        x"71", x"72", x"71", x"70", x"6f", x"6f", x"6e", x"6f", x"6f", x"6f", x"6f", x"6f", x"70", x"70", x"6f", 
        x"70", x"71", x"70", x"70", x"6e", x"6d", x"6c", x"6c", x"6d", x"6d", x"6e", x"6f", x"70", x"70", x"6e", 
        x"6f", x"6d", x"6d", x"6f", x"6f", x"6d", x"6f", x"6f", x"6e", x"6e", x"6c", x"6d", x"6d", x"6c", x"6c", 
        x"70", x"6f", x"6d", x"70", x"6f", x"6e", x"6e", x"6e", x"6f", x"71", x"6f", x"6d", x"6e", x"6d", x"6d", 
        x"6e", x"6d", x"6e", x"6d", x"6e", x"6e", x"6f", x"6f", x"6e", x"6f", x"6e", x"6e", x"70", x"6f", x"6e", 
        x"6f", x"6f", x"6d", x"6f", x"6f", x"6c", x"6e", x"6d", x"6c", x"6c", x"6e", x"70", x"6f", x"6d", x"6e", 
        x"70", x"6e", x"6b", x"6b", x"6c", x"6c", x"6b", x"6b", x"6b", x"6c", x"6e", x"70", x"6e", x"6b", x"6a", 
        x"6b", x"6b", x"69", x"69", x"6c", x"6c", x"6e", x"6c", x"6c", x"6d", x"6e", x"6d", x"6e", x"6d", x"6c", 
        x"6a", x"6b", x"6c", x"6e", x"6f", x"6e", x"6c", x"6a", x"69", x"6a", x"6b", x"6d", x"6e", x"6e", x"6e", 
        x"6d", x"6d", x"6c", x"6c", x"6d", x"6d", x"6c", x"6a", x"6b", x"6c", x"6a", x"6c", x"6d", x"6d", x"69", 
        x"6c", x"6c", x"6c", x"6d", x"6e", x"6e", x"6e", x"6f", x"70", x"6e", x"70", x"6f", x"6d", x"6b", x"6b", 
        x"68", x"6d", x"6e", x"6a", x"6c", x"6a", x"69", x"6b", x"6b", x"6b", x"6b", x"6c", x"6d", x"6c", x"67", 
        x"6b", x"6d", x"6a", x"69", x"6b", x"6c", x"6a", x"6b", x"69", x"69", x"6a", x"6a", x"6d", x"6a", x"68", 
        x"68", x"6a", x"6c", x"6d", x"6b", x"6a", x"6c", x"6c", x"6c", x"6a", x"69", x"69", x"6b", x"6c", x"6b", 
        x"6b", x"6b", x"69", x"68", x"6a", x"6c", x"6b", x"6a", x"68", x"69", x"6b", x"6b", x"6a", x"6b", x"66", 
        x"66", x"6a", x"6a", x"67", x"68", x"67", x"68", x"6a", x"6b", x"6a", x"67", x"69", x"69", x"6b", x"69", 
        x"69", x"67", x"68", x"6a", x"69", x"68", x"66", x"65", x"65", x"66", x"66", x"67", x"67", x"66", x"67", 
        x"66", x"65", x"66", x"66", x"69", x"69", x"67", x"65", x"66", x"67", x"66", x"64", x"64", x"66", x"66", 
        x"66", x"66", x"64", x"61", x"63", x"65", x"65", x"68", x"68", x"68", x"68", x"67", x"66", x"64", x"65", 
        x"66", x"65", x"66", x"67", x"66", x"64", x"63", x"65", x"66", x"64", x"64", x"65", x"65", x"65", x"64", 
        x"65", x"66", x"64", x"65", x"66", x"65", x"64", x"65", x"63", x"62", x"62", x"62", x"62", x"62", x"63", 
        x"63", x"63", x"63", x"61", x"61", x"60", x"60", x"62", x"63", x"62", x"61", x"62", x"61", x"60", x"60", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"62", x"61", x"61", x"62", x"61", x"61", 
        x"61", x"60", x"60", x"60", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"60", x"60", 
        x"65", x"64", x"65", x"64", x"65", x"65", x"65", x"66", x"63", x"65", x"65", x"64", x"66", x"67", x"64", 
        x"63", x"63", x"65", x"66", x"65", x"62", x"62", x"64", x"64", x"64", x"64", x"64", x"64", x"65", x"67", 
        x"67", x"65", x"63", x"65", x"65", x"63", x"63", x"64", x"66", x"68", x"66", x"64", x"64", x"65", x"65", 
        x"64", x"64", x"65", x"66", x"66", x"67", x"67", x"67", x"67", x"67", x"66", x"65", x"65", x"64", x"64", 
        x"64", x"66", x"68", x"68", x"68", x"67", x"66", x"65", x"65", x"66", x"67", x"66", x"65", x"65", x"65", 
        x"65", x"65", x"64", x"64", x"63", x"62", x"65", x"65", x"66", x"64", x"65", x"66", x"66", x"66", x"67", 
        x"66", x"67", x"67", x"67", x"6a", x"68", x"69", x"68", x"67", x"68", x"66", x"68", x"69", x"66", x"67", 
        x"6a", x"6b", x"6a", x"69", x"67", x"69", x"67", x"67", x"69", x"67", x"6a", x"68", x"67", x"66", x"68", 
        x"69", x"6b", x"6a", x"69", x"67", x"67", x"68", x"67", x"65", x"6a", x"6a", x"67", x"67", x"67", x"67", 
        x"69", x"69", x"67", x"68", x"69", x"69", x"68", x"67", x"67", x"6b", x"6d", x"6b", x"6a", x"6d", x"6f", 
        x"6e", x"6a", x"6d", x"6c", x"6b", x"6b", x"69", x"6a", x"6c", x"6c", x"6b", x"67", x"6a", x"6a", x"69", 
        x"6b", x"72", x"71", x"6e", x"6c", x"61", x"69", x"8f", x"c6", x"b9", x"8f", x"a2", x"ce", x"d2", x"ca", 
        x"cc", x"cd", x"cb", x"c7", x"ca", x"ce", x"ca", x"cc", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"ce", 
        x"ce", x"ce", x"ce", x"cf", x"cd", x"cc", x"cf", x"cd", x"cf", x"cf", x"cf", x"cf", x"d0", x"cf", x"b0", 
        x"6e", x"5d", x"5f", x"5f", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5d", x"5c", x"67", x"7e", x"a1", x"cd", x"e7", 
        x"f0", x"f5", x"f2", x"e7", x"d9", x"c7", x"b8", x"a6", x"92", x"89", x"8a", x"95", x"af", x"d3", x"e8", 
        x"e6", x"d3", x"a5", x"77", x"68", x"68", x"72", x"74", x"72", x"6d", x"72", x"73", x"72", x"73", x"73", 
        x"74", x"73", x"73", x"73", x"71", x"70", x"70", x"70", x"71", x"70", x"70", x"70", x"71", x"71", x"72", 
        x"72", x"70", x"6d", x"6d", x"6f", x"71", x"6f", x"6d", x"6e", x"70", x"71", x"6f", x"6d", x"6e", x"70", 
        x"6e", x"6e", x"72", x"6f", x"6c", x"6d", x"6d", x"70", x"71", x"6f", x"70", x"70", x"6e", x"70", x"6f", 
        x"6c", x"6f", x"71", x"70", x"70", x"71", x"70", x"6f", x"6f", x"6e", x"6d", x"6e", x"6f", x"73", x"70", 
        x"72", x"71", x"6f", x"6e", x"6f", x"6e", x"6f", x"71", x"70", x"6e", x"6f", x"70", x"70", x"6d", x"6e", 
        x"6e", x"6d", x"6c", x"6d", x"70", x"74", x"70", x"6d", x"6f", x"71", x"72", x"71", x"6f", x"6f", x"6f", 
        x"70", x"72", x"72", x"70", x"6e", x"6d", x"6f", x"6e", x"6d", x"6e", x"6f", x"70", x"70", x"71", x"6e", 
        x"6f", x"6d", x"6d", x"70", x"6f", x"6e", x"71", x"71", x"70", x"70", x"6e", x"6f", x"70", x"6e", x"6c", 
        x"6e", x"6e", x"6e", x"6f", x"6e", x"6f", x"6f", x"6e", x"70", x"72", x"6f", x"6d", x"71", x"71", x"71", 
        x"71", x"6f", x"71", x"71", x"71", x"6e", x"6f", x"6f", x"70", x"72", x"6f", x"6e", x"6e", x"6d", x"6e", 
        x"71", x"71", x"6e", x"72", x"70", x"6c", x"6f", x"6e", x"6e", x"6e", x"70", x"70", x"6e", x"6c", x"6c", 
        x"6e", x"6e", x"6e", x"70", x"70", x"6e", x"6c", x"6c", x"6d", x"6e", x"6e", x"6e", x"6e", x"6e", x"6d", 
        x"6c", x"6c", x"6e", x"6c", x"6c", x"6a", x"6e", x"6f", x"72", x"6d", x"6e", x"6e", x"70", x"6e", x"6e", 
        x"6e", x"6e", x"6e", x"6e", x"6d", x"6c", x"6b", x"6b", x"6b", x"6b", x"6c", x"6d", x"6d", x"6c", x"6b", 
        x"6b", x"6e", x"6b", x"6b", x"6d", x"6f", x"6e", x"6d", x"6d", x"6e", x"6c", x"6d", x"6d", x"6e", x"6b", 
        x"6c", x"6b", x"6b", x"6c", x"6e", x"6e", x"6d", x"6d", x"6f", x"6d", x"6f", x"6e", x"6d", x"6c", x"6c", 
        x"67", x"6c", x"6d", x"68", x"6b", x"6b", x"6b", x"6e", x"6d", x"6b", x"6b", x"6a", x"69", x"6a", x"6b", 
        x"6b", x"6b", x"6a", x"6a", x"6c", x"6e", x"6c", x"6d", x"6a", x"6a", x"6a", x"68", x"6b", x"6a", x"69", 
        x"68", x"69", x"6a", x"6b", x"6b", x"6a", x"6d", x"6b", x"6c", x"6a", x"69", x"6a", x"6b", x"6a", x"68", 
        x"69", x"6b", x"6a", x"6a", x"6b", x"6b", x"6b", x"6b", x"6a", x"6a", x"6b", x"6d", x"6d", x"69", x"67", 
        x"67", x"69", x"6b", x"69", x"68", x"66", x"66", x"68", x"6b", x"6c", x"6b", x"6c", x"68", x"6b", x"6b", 
        x"68", x"68", x"69", x"69", x"68", x"68", x"68", x"68", x"68", x"67", x"67", x"68", x"68", x"65", x"67", 
        x"66", x"63", x"66", x"66", x"68", x"68", x"67", x"65", x"65", x"65", x"65", x"66", x"65", x"65", x"66", 
        x"67", x"68", x"6b", x"66", x"65", x"66", x"67", x"69", x"67", x"67", x"68", x"67", x"65", x"66", x"66", 
        x"67", x"67", x"66", x"66", x"66", x"65", x"65", x"68", x"69", x"67", x"66", x"66", x"66", x"66", x"66", 
        x"65", x"64", x"63", x"65", x"67", x"66", x"66", x"67", x"63", x"62", x"62", x"62", x"62", x"62", x"63", 
        x"64", x"64", x"63", x"62", x"61", x"61", x"61", x"63", x"64", x"63", x"63", x"63", x"62", x"61", x"60", 
        x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"61", x"61", x"61", x"62", x"62", x"61", x"61", 
        x"62", x"61", x"60", x"60", x"61", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"66", x"65", x"67", x"65", x"66", x"66", x"66", x"66", x"63", x"64", x"64", x"63", x"65", x"66", x"64", 
        x"64", x"64", x"65", x"66", x"66", x"64", x"63", x"63", x"64", x"64", x"64", x"63", x"65", x"66", x"64", 
        x"64", x"63", x"64", x"67", x"68", x"66", x"65", x"65", x"65", x"67", x"65", x"64", x"64", x"65", x"66", 
        x"67", x"66", x"65", x"66", x"67", x"68", x"68", x"68", x"67", x"66", x"64", x"64", x"66", x"66", x"65", 
        x"65", x"66", x"67", x"67", x"66", x"67", x"66", x"64", x"65", x"66", x"65", x"65", x"63", x"62", x"63", 
        x"65", x"67", x"65", x"63", x"65", x"65", x"67", x"66", x"67", x"64", x"65", x"66", x"65", x"65", x"68", 
        x"67", x"65", x"67", x"67", x"69", x"68", x"65", x"65", x"64", x"65", x"66", x"68", x"67", x"65", x"64", 
        x"67", x"69", x"69", x"69", x"68", x"69", x"67", x"68", x"6a", x"67", x"68", x"69", x"69", x"68", x"67", 
        x"68", x"69", x"6c", x"6c", x"6a", x"69", x"6a", x"6a", x"69", x"6a", x"69", x"65", x"65", x"66", x"67", 
        x"69", x"69", x"67", x"68", x"69", x"6a", x"6a", x"6a", x"69", x"6a", x"6b", x"6a", x"69", x"6b", x"6c", 
        x"6c", x"6c", x"6e", x"6b", x"6b", x"6c", x"6c", x"6b", x"6f", x"6e", x"6e", x"6a", x"6a", x"68", x"69", 
        x"6b", x"6e", x"6d", x"6c", x"64", x"74", x"a7", x"c8", x"ae", x"94", x"b2", x"d3", x"ce", x"cb", x"c8", 
        x"cc", x"cc", x"cb", x"cc", x"ca", x"cb", x"ce", x"cd", x"cd", x"cc", x"cc", x"cd", x"cd", x"cd", x"cd", 
        x"cd", x"cd", x"cd", x"ce", x"cd", x"cc", x"cf", x"ce", x"cf", x"ce", x"ce", x"ce", x"d1", x"d0", x"af", 
        x"6d", x"5d", x"5f", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5c", x"5e", x"5f", x"5b", x"62", x"7e", x"ab", x"d4", x"ed", x"f7", x"f5", 
        x"ec", x"d8", x"b9", x"9c", x"82", x"6c", x"65", x"63", x"5e", x"5c", x"5c", x"5e", x"69", x"81", x"a7", 
        x"ca", x"e1", x"e8", x"d9", x"af", x"86", x"6f", x"68", x"6e", x"75", x"73", x"70", x"70", x"70", x"72", 
        x"70", x"6f", x"71", x"70", x"70", x"71", x"71", x"72", x"71", x"70", x"72", x"73", x"72", x"70", x"70", 
        x"71", x"72", x"6e", x"6d", x"6f", x"72", x"71", x"6e", x"6e", x"6f", x"70", x"6f", x"6d", x"6e", x"70", 
        x"6f", x"70", x"72", x"6f", x"70", x"73", x"71", x"71", x"71", x"70", x"72", x"71", x"6e", x"70", x"70", 
        x"6c", x"6e", x"70", x"6e", x"6d", x"6f", x"70", x"6f", x"70", x"70", x"6f", x"6f", x"70", x"73", x"70", 
        x"70", x"6f", x"6f", x"70", x"6e", x"6b", x"6d", x"6f", x"6e", x"6e", x"6f", x"70", x"71", x"6f", x"6d", 
        x"6d", x"6e", x"6f", x"6f", x"6f", x"6f", x"70", x"6f", x"6f", x"71", x"72", x"71", x"71", x"71", x"71", 
        x"6f", x"6e", x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"70", x"70", x"70", x"71", x"73", x"6e", 
        x"6e", x"6f", x"6f", x"70", x"6c", x"6d", x"70", x"71", x"6e", x"6e", x"6d", x"6f", x"71", x"70", x"6c", 
        x"6d", x"6e", x"6e", x"6f", x"6f", x"70", x"71", x"6f", x"70", x"71", x"6f", x"6c", x"6f", x"71", x"71", 
        x"71", x"6e", x"6f", x"70", x"73", x"70", x"70", x"70", x"70", x"71", x"70", x"73", x"71", x"6e", x"6e", 
        x"70", x"70", x"6d", x"6f", x"6c", x"6a", x"6d", x"6b", x"6d", x"6e", x"6f", x"70", x"6f", x"6f", x"6e", 
        x"6f", x"6f", x"6f", x"6f", x"70", x"6e", x"6c", x"6c", x"6f", x"6f", x"6d", x"6e", x"6f", x"70", x"6f", 
        x"6d", x"6e", x"6e", x"6e", x"6f", x"6d", x"6d", x"6c", x"6d", x"6b", x"6d", x"6d", x"6f", x"6e", x"6f", 
        x"70", x"71", x"70", x"6d", x"6d", x"6d", x"6d", x"6f", x"6f", x"6d", x"6e", x"6e", x"6e", x"6d", x"6d", 
        x"6e", x"6f", x"6c", x"6c", x"6e", x"6e", x"6e", x"6d", x"6b", x"6f", x"6e", x"6b", x"69", x"6c", x"6d", 
        x"6d", x"6c", x"6b", x"6c", x"6d", x"6e", x"6e", x"6c", x"6e", x"6d", x"6e", x"6d", x"6d", x"6c", x"6d", 
        x"6c", x"6e", x"6d", x"69", x"6d", x"6c", x"6d", x"6e", x"6c", x"6b", x"6b", x"6c", x"6a", x"6a", x"6e", 
        x"6c", x"6a", x"6a", x"6b", x"6d", x"6d", x"6d", x"6d", x"6c", x"6b", x"6a", x"69", x"6a", x"6a", x"6b", 
        x"6a", x"6a", x"6a", x"6a", x"6c", x"6d", x"6d", x"6b", x"6c", x"6c", x"6b", x"6c", x"6a", x"69", x"67", 
        x"67", x"6b", x"69", x"69", x"6b", x"6c", x"6c", x"6b", x"6a", x"67", x"68", x"69", x"69", x"64", x"64", 
        x"65", x"67", x"69", x"6a", x"6b", x"6b", x"68", x"67", x"67", x"68", x"6a", x"6b", x"68", x"6a", x"6b", 
        x"69", x"69", x"69", x"68", x"67", x"68", x"69", x"67", x"67", x"67", x"67", x"69", x"68", x"65", x"68", 
        x"66", x"64", x"66", x"66", x"66", x"66", x"66", x"66", x"65", x"64", x"64", x"68", x"68", x"66", x"67", 
        x"68", x"68", x"69", x"66", x"65", x"67", x"68", x"69", x"67", x"66", x"68", x"67", x"66", x"67", x"67", 
        x"66", x"68", x"67", x"66", x"66", x"66", x"66", x"67", x"68", x"68", x"67", x"67", x"65", x"65", x"65", 
        x"67", x"69", x"68", x"68", x"67", x"64", x"63", x"65", x"64", x"63", x"63", x"62", x"61", x"62", x"63", 
        x"64", x"63", x"63", x"62", x"61", x"62", x"62", x"63", x"64", x"63", x"63", x"63", x"62", x"61", x"61", 
        x"62", x"62", x"61", x"61", x"61", x"62", x"62", x"62", x"61", x"61", x"62", x"63", x"62", x"61", x"61", 
        x"62", x"63", x"62", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"62", x"61", 
        x"65", x"64", x"66", x"66", x"65", x"66", x"65", x"64", x"64", x"63", x"64", x"64", x"64", x"63", x"64", 
        x"64", x"64", x"64", x"64", x"65", x"66", x"64", x"64", x"65", x"63", x"64", x"64", x"66", x"69", x"65", 
        x"65", x"64", x"65", x"66", x"66", x"66", x"65", x"67", x"64", x"64", x"64", x"62", x"66", x"66", x"65", 
        x"64", x"65", x"65", x"65", x"64", x"65", x"65", x"67", x"67", x"65", x"63", x"65", x"67", x"66", x"67", 
        x"68", x"68", x"67", x"66", x"64", x"66", x"66", x"65", x"66", x"69", x"65", x"64", x"64", x"64", x"64", 
        x"64", x"64", x"65", x"67", x"67", x"68", x"67", x"66", x"67", x"66", x"69", x"69", x"66", x"65", x"66", 
        x"65", x"65", x"67", x"65", x"6a", x"6d", x"67", x"66", x"67", x"67", x"69", x"68", x"68", x"67", x"68", 
        x"69", x"6a", x"69", x"67", x"68", x"67", x"67", x"67", x"67", x"65", x"65", x"6a", x"6b", x"68", x"67", 
        x"68", x"6a", x"68", x"68", x"69", x"69", x"69", x"6a", x"6b", x"6b", x"69", x"67", x"67", x"69", x"6a", 
        x"69", x"69", x"69", x"6a", x"6b", x"6a", x"6a", x"6b", x"69", x"68", x"69", x"6a", x"69", x"68", x"67", 
        x"67", x"6c", x"6c", x"68", x"69", x"6b", x"70", x"6e", x"6c", x"6d", x"70", x"6f", x"6c", x"6a", x"6a", 
        x"6d", x"6f", x"6b", x"6b", x"7f", x"b7", x"c4", x"a0", x"95", x"be", x"d2", x"ce", x"ce", x"ca", x"cc", 
        x"cd", x"cd", x"cd", x"cd", x"cd", x"cc", x"cd", x"cd", x"cd", x"cc", x"cc", x"cc", x"cc", x"cb", x"cb", 
        x"cc", x"cb", x"cb", x"cd", x"cd", x"cb", x"cc", x"ce", x"d0", x"cf", x"cd", x"ce", x"d1", x"d3", x"ab", 
        x"6a", x"5e", x"5e", x"5f", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5e", 
        x"5e", x"5f", x"5d", x"5d", x"5f", x"5c", x"60", x"74", x"9c", x"ce", x"f0", x"f6", x"f5", x"e6", x"cb", 
        x"a8", x"83", x"69", x"5f", x"5d", x"5d", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5f", x"60", x"66", 
        x"7d", x"9f", x"bf", x"dd", x"e5", x"dd", x"b9", x"92", x"75", x"6b", x"6c", x"6d", x"73", x"74", x"75", 
        x"71", x"70", x"70", x"6e", x"71", x"74", x"72", x"73", x"72", x"6f", x"72", x"71", x"71", x"71", x"72", 
        x"73", x"73", x"70", x"6f", x"70", x"73", x"74", x"72", x"6f", x"71", x"72", x"72", x"71", x"71", x"71", 
        x"72", x"70", x"71", x"73", x"74", x"74", x"73", x"72", x"71", x"71", x"71", x"70", x"6e", x"70", x"71", 
        x"70", x"70", x"72", x"72", x"6f", x"6f", x"70", x"72", x"72", x"72", x"6f", x"70", x"73", x"73", x"70", 
        x"70", x"70", x"6d", x"6e", x"6f", x"6d", x"70", x"6f", x"6e", x"70", x"6e", x"6c", x"6f", x"71", x"6f", 
        x"6d", x"6c", x"6d", x"6f", x"71", x"71", x"74", x"71", x"6f", x"70", x"71", x"70", x"72", x"73", x"71", 
        x"6d", x"6f", x"72", x"72", x"6e", x"6d", x"6c", x"70", x"71", x"71", x"6f", x"6f", x"70", x"72", x"70", 
        x"70", x"72", x"71", x"6d", x"6c", x"6f", x"70", x"74", x"6e", x"6e", x"73", x"73", x"70", x"70", x"6e", 
        x"6e", x"70", x"6e", x"6f", x"71", x"71", x"71", x"70", x"6e", x"6d", x"6f", x"6f", x"6f", x"71", x"70", 
        x"71", x"6f", x"6d", x"6f", x"6f", x"71", x"6f", x"70", x"6f", x"6c", x"6f", x"70", x"6e", x"6e", x"70", 
        x"72", x"71", x"6f", x"6f", x"6b", x"6f", x"6f", x"69", x"6e", x"6e", x"6e", x"6e", x"6d", x"6e", x"6e", 
        x"6c", x"6c", x"6d", x"6e", x"70", x"71", x"6f", x"70", x"72", x"73", x"70", x"70", x"70", x"72", x"71", 
        x"6d", x"6d", x"6b", x"6e", x"71", x"70", x"6d", x"6b", x"6c", x"6d", x"6e", x"6e", x"6e", x"6f", x"6f", 
        x"70", x"6f", x"6f", x"6d", x"71", x"6f", x"6c", x"6d", x"6d", x"6c", x"6e", x"70", x"71", x"6c", x"6c", 
        x"6e", x"71", x"6f", x"6f", x"6f", x"6b", x"69", x"6b", x"6e", x"6f", x"6e", x"6c", x"6c", x"6d", x"6d", 
        x"6d", x"6b", x"6c", x"6d", x"6b", x"6b", x"6e", x"6c", x"6e", x"6f", x"6d", x"6c", x"6c", x"6a", x"6c", 
        x"70", x"6e", x"6a", x"6b", x"6b", x"6a", x"6c", x"6c", x"6a", x"6d", x"6a", x"6c", x"6c", x"6b", x"6e", 
        x"6c", x"6b", x"6c", x"6d", x"6c", x"6c", x"70", x"6d", x"6d", x"6c", x"6c", x"6d", x"6a", x"6a", x"6c", 
        x"69", x"6a", x"6c", x"6a", x"6c", x"6e", x"6b", x"68", x"6a", x"6c", x"6b", x"6a", x"6a", x"6b", x"6b", 
        x"66", x"6c", x"69", x"68", x"6a", x"69", x"69", x"69", x"6a", x"66", x"69", x"68", x"6b", x"6a", x"68", 
        x"6a", x"6a", x"69", x"6c", x"6a", x"68", x"66", x"65", x"69", x"6b", x"67", x"67", x"67", x"68", x"6b", 
        x"6c", x"6b", x"68", x"69", x"69", x"6b", x"6c", x"67", x"67", x"68", x"68", x"6a", x"68", x"67", x"6a", 
        x"6a", x"68", x"67", x"67", x"66", x"65", x"66", x"68", x"68", x"65", x"65", x"6b", x"6e", x"6b", x"69", 
        x"6a", x"6a", x"6c", x"69", x"68", x"6b", x"69", x"67", x"68", x"68", x"6b", x"6a", x"69", x"66", x"68", 
        x"67", x"66", x"66", x"65", x"65", x"66", x"66", x"66", x"65", x"68", x"67", x"68", x"66", x"66", x"66", 
        x"69", x"69", x"6a", x"6a", x"67", x"64", x"65", x"67", x"65", x"64", x"66", x"63", x"5f", x"62", x"64", 
        x"65", x"62", x"63", x"63", x"62", x"65", x"63", x"61", x"61", x"62", x"63", x"63", x"62", x"61", x"61", 
        x"61", x"62", x"62", x"62", x"62", x"62", x"62", x"61", x"61", x"62", x"63", x"63", x"63", x"63", x"62", 
        x"63", x"62", x"60", x"61", x"62", x"61", x"60", x"61", x"62", x"62", x"61", x"61", x"61", x"61", x"62", 
        x"66", x"66", x"66", x"65", x"65", x"65", x"64", x"66", x"66", x"64", x"65", x"66", x"65", x"64", x"65", 
        x"65", x"65", x"64", x"63", x"64", x"66", x"66", x"65", x"65", x"63", x"63", x"63", x"63", x"65", x"65", 
        x"65", x"65", x"66", x"66", x"65", x"64", x"64", x"65", x"63", x"63", x"65", x"64", x"67", x"67", x"66", 
        x"65", x"64", x"64", x"63", x"64", x"65", x"63", x"62", x"65", x"68", x"68", x"66", x"67", x"67", x"68", 
        x"68", x"66", x"66", x"68", x"66", x"64", x"64", x"62", x"64", x"69", x"67", x"67", x"64", x"65", x"66", 
        x"65", x"65", x"65", x"67", x"66", x"66", x"65", x"64", x"64", x"67", x"69", x"65", x"64", x"67", x"67", 
        x"65", x"64", x"67", x"67", x"6a", x"6b", x"66", x"68", x"6a", x"69", x"67", x"67", x"67", x"68", x"6a", 
        x"6b", x"6c", x"6a", x"67", x"68", x"69", x"6a", x"6a", x"6a", x"68", x"68", x"6b", x"6a", x"67", x"66", 
        x"68", x"6a", x"67", x"6a", x"6b", x"6a", x"68", x"68", x"6c", x"6b", x"6a", x"6a", x"6a", x"6b", x"6b", 
        x"69", x"6b", x"6b", x"6c", x"6d", x"6b", x"6d", x"6d", x"6b", x"68", x"6a", x"6b", x"6c", x"6c", x"6b", 
        x"6a", x"69", x"6c", x"6a", x"6a", x"6b", x"6f", x"6f", x"69", x"6d", x"6f", x"6f", x"6e", x"6d", x"6c", 
        x"6d", x"6c", x"6c", x"90", x"c7", x"ba", x"92", x"a0", x"c9", x"d0", x"c7", x"ce", x"cc", x"c9", x"d0", 
        x"cd", x"cd", x"ce", x"ce", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"cc", x"cc", x"cc", 
        x"cd", x"cc", x"cb", x"cb", x"cc", x"cb", x"cc", x"cf", x"cf", x"ce", x"cc", x"ce", x"d2", x"d2", x"aa", 
        x"69", x"5d", x"5d", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"61", x"5c", 
        x"60", x"5e", x"5e", x"5e", x"61", x"64", x"88", x"ce", x"ee", x"f5", x"f6", x"e5", x"c4", x"92", x"6e", 
        x"5f", x"5b", x"5d", x"5d", x"5d", x"5f", x"60", x"60", x"5e", x"5e", x"5d", x"5d", x"5f", x"5e", x"5c", 
        x"5c", x"61", x"6c", x"8a", x"ae", x"d1", x"e8", x"e7", x"cb", x"9d", x"7c", x"69", x"6a", x"6d", x"71", 
        x"77", x"75", x"75", x"73", x"73", x"73", x"6e", x"70", x"72", x"6e", x"6a", x"6d", x"6f", x"71", x"72", 
        x"71", x"72", x"75", x"74", x"73", x"74", x"75", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", 
        x"73", x"72", x"72", x"72", x"72", x"71", x"71", x"71", x"72", x"72", x"72", x"71", x"6f", x"6f", x"70", 
        x"70", x"71", x"71", x"6f", x"6e", x"6e", x"71", x"72", x"72", x"72", x"70", x"70", x"73", x"71", x"6f", 
        x"71", x"6f", x"6c", x"6f", x"72", x"70", x"70", x"6f", x"6d", x"6f", x"6c", x"6a", x"6e", x"71", x"71", 
        x"70", x"6f", x"6f", x"70", x"71", x"72", x"72", x"71", x"70", x"70", x"70", x"70", x"71", x"74", x"74", 
        x"72", x"73", x"75", x"73", x"71", x"71", x"6f", x"6f", x"70", x"70", x"70", x"6f", x"6d", x"6e", x"6d", 
        x"6e", x"71", x"72", x"70", x"6f", x"70", x"6f", x"72", x"6d", x"6e", x"71", x"71", x"6f", x"70", x"6f", 
        x"6e", x"70", x"6f", x"6f", x"6f", x"6e", x"6f", x"6f", x"6e", x"6e", x"70", x"70", x"70", x"71", x"70", 
        x"71", x"70", x"6e", x"70", x"6e", x"6f", x"6e", x"71", x"72", x"70", x"71", x"71", x"6f", x"6e", x"71", 
        x"72", x"71", x"70", x"6f", x"6f", x"72", x"6d", x"69", x"70", x"6e", x"6e", x"6f", x"6d", x"6e", x"6d", 
        x"6c", x"6e", x"70", x"70", x"72", x"72", x"71", x"71", x"72", x"71", x"6f", x"70", x"70", x"70", x"70", 
        x"6e", x"6c", x"6c", x"6f", x"70", x"6f", x"6d", x"6d", x"6c", x"6e", x"6f", x"6e", x"6e", x"6e", x"6f", 
        x"6f", x"6e", x"6f", x"6d", x"6f", x"6e", x"6e", x"70", x"6f", x"6d", x"6d", x"6e", x"6f", x"6b", x"6b", 
        x"6c", x"6d", x"6c", x"6f", x"70", x"6e", x"6d", x"6f", x"71", x"6f", x"6c", x"6c", x"6e", x"6d", x"6a", 
        x"6e", x"6e", x"6e", x"6e", x"6b", x"6a", x"69", x"6e", x"70", x"6e", x"6c", x"6d", x"6d", x"68", x"69", 
        x"6f", x"6d", x"6a", x"6c", x"6b", x"6a", x"6b", x"69", x"68", x"6a", x"66", x"69", x"6d", x"6e", x"6d", 
        x"6c", x"6b", x"6d", x"6e", x"6e", x"6d", x"6e", x"6b", x"6d", x"6c", x"6c", x"6d", x"6b", x"69", x"6c", 
        x"6a", x"6b", x"6c", x"69", x"69", x"6d", x"6c", x"6a", x"6c", x"6e", x"6d", x"6e", x"6e", x"6c", x"6f", 
        x"6d", x"6f", x"6d", x"6c", x"6a", x"6a", x"69", x"69", x"6b", x"69", x"6c", x"6b", x"6c", x"6c", x"6c", 
        x"69", x"6b", x"6e", x"6b", x"67", x"68", x"68", x"66", x"68", x"69", x"67", x"64", x"67", x"6a", x"6c", 
        x"6a", x"6a", x"6b", x"6a", x"68", x"69", x"6a", x"66", x"65", x"66", x"67", x"6a", x"68", x"68", x"69", 
        x"6b", x"6c", x"6b", x"6a", x"69", x"68", x"68", x"6a", x"6a", x"68", x"64", x"68", x"6b", x"6a", x"69", 
        x"6a", x"6b", x"6c", x"68", x"66", x"6a", x"6c", x"6a", x"67", x"66", x"68", x"68", x"68", x"66", x"69", 
        x"68", x"69", x"69", x"66", x"65", x"65", x"65", x"65", x"67", x"6a", x"69", x"6b", x"64", x"66", x"69", 
        x"69", x"66", x"68", x"6a", x"69", x"67", x"65", x"64", x"63", x"62", x"65", x"64", x"62", x"64", x"64", 
        x"66", x"64", x"64", x"64", x"62", x"64", x"63", x"62", x"62", x"62", x"62", x"62", x"62", x"62", x"62", 
        x"63", x"63", x"63", x"62", x"62", x"62", x"62", x"61", x"61", x"61", x"61", x"63", x"64", x"64", x"63", 
        x"64", x"63", x"62", x"63", x"64", x"62", x"60", x"61", x"62", x"62", x"61", x"61", x"61", x"62", x"62", 
        x"67", x"67", x"65", x"65", x"65", x"64", x"66", x"67", x"65", x"65", x"66", x"67", x"66", x"65", x"66", 
        x"66", x"65", x"64", x"63", x"64", x"66", x"67", x"66", x"65", x"64", x"65", x"65", x"64", x"65", x"64", 
        x"63", x"64", x"66", x"67", x"66", x"64", x"66", x"65", x"63", x"64", x"65", x"64", x"65", x"67", x"67", 
        x"66", x"65", x"64", x"64", x"65", x"64", x"63", x"64", x"66", x"68", x"67", x"66", x"66", x"67", x"69", 
        x"69", x"67", x"66", x"67", x"68", x"67", x"66", x"62", x"63", x"66", x"64", x"65", x"65", x"66", x"67", 
        x"67", x"67", x"66", x"67", x"6a", x"68", x"68", x"67", x"64", x"68", x"69", x"65", x"65", x"67", x"68", 
        x"66", x"65", x"68", x"68", x"6b", x"6c", x"68", x"67", x"68", x"68", x"66", x"67", x"68", x"69", x"6a", 
        x"6a", x"6a", x"69", x"67", x"67", x"6a", x"6c", x"6c", x"6c", x"6d", x"6a", x"6a", x"69", x"67", x"68", 
        x"69", x"69", x"6a", x"6a", x"6a", x"6a", x"6a", x"6a", x"6a", x"6a", x"6a", x"68", x"67", x"67", x"69", 
        x"6a", x"6b", x"6a", x"6a", x"6c", x"6a", x"6b", x"6c", x"69", x"67", x"68", x"69", x"6b", x"6b", x"6b", 
        x"6a", x"69", x"6c", x"6c", x"6b", x"6b", x"6e", x"6e", x"6d", x"6e", x"6f", x"6c", x"6c", x"6f", x"6e", 
        x"68", x"7b", x"ad", x"c4", x"a8", x"9a", x"b9", x"cf", x"ce", x"c8", x"cb", x"cd", x"c8", x"c9", x"cb", 
        x"cc", x"cd", x"ce", x"ce", x"cd", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"cd", x"cc", x"cb", x"cc", 
        x"cd", x"cc", x"cb", x"cb", x"cb", x"ca", x"ce", x"cf", x"ce", x"cd", x"cc", x"cf", x"d3", x"d1", x"ab", 
        x"69", x"5c", x"5d", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"5f", 
        x"5d", x"5f", x"60", x"5d", x"75", x"ab", x"dc", x"f3", x"f7", x"ed", x"c7", x"9a", x"75", x"5f", x"5b", 
        x"5f", x"5e", x"5f", x"5f", x"5e", x"5f", x"60", x"60", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5f", 
        x"5f", x"5e", x"5d", x"60", x"6e", x"81", x"9f", x"bf", x"d9", x"e5", x"d3", x"b5", x"8d", x"6f", x"68", 
        x"6d", x"73", x"78", x"73", x"6f", x"70", x"72", x"74", x"73", x"71", x"71", x"72", x"73", x"74", x"74", 
        x"74", x"74", x"74", x"74", x"73", x"72", x"72", x"72", x"73", x"74", x"73", x"73", x"74", x"74", x"74", 
        x"73", x"72", x"72", x"72", x"72", x"72", x"73", x"73", x"72", x"72", x"72", x"71", x"6f", x"6f", x"6e", 
        x"6e", x"6f", x"71", x"71", x"70", x"6f", x"6f", x"70", x"70", x"71", x"71", x"72", x"74", x"73", x"70", 
        x"6f", x"70", x"70", x"71", x"71", x"70", x"71", x"6e", x"6e", x"70", x"6e", x"6c", x"6e", x"70", x"71", 
        x"71", x"71", x"70", x"6f", x"71", x"72", x"71", x"70", x"71", x"71", x"70", x"6f", x"70", x"72", x"73", 
        x"74", x"73", x"72", x"70", x"70", x"70", x"70", x"71", x"71", x"6f", x"6d", x"6f", x"6f", x"6d", x"6e", 
        x"6f", x"6f", x"71", x"71", x"6f", x"72", x"71", x"72", x"6f", x"70", x"71", x"70", x"6f", x"70", x"6f", 
        x"6f", x"70", x"6f", x"6f", x"6e", x"6e", x"70", x"71", x"6f", x"6f", x"6f", x"6e", x"6d", x"6f", x"6e", 
        x"6e", x"6d", x"6d", x"6f", x"72", x"73", x"72", x"71", x"70", x"6d", x"6e", x"75", x"73", x"70", x"70", 
        x"70", x"6f", x"6e", x"6e", x"70", x"72", x"6e", x"6a", x"71", x"70", x"6f", x"70", x"6e", x"6e", x"6e", 
        x"6e", x"70", x"70", x"70", x"71", x"70", x"71", x"72", x"72", x"71", x"6e", x"6e", x"6f", x"6e", x"6f", 
        x"6f", x"6b", x"6e", x"6f", x"6f", x"6f", x"6f", x"6e", x"6d", x"70", x"70", x"6f", x"6e", x"6e", x"6e", 
        x"6e", x"6c", x"6d", x"6d", x"6d", x"6e", x"70", x"71", x"6f", x"6c", x"6d", x"6c", x"6e", x"6c", x"6d", 
        x"6d", x"6d", x"6d", x"6f", x"70", x"6e", x"6e", x"71", x"73", x"6f", x"6c", x"6c", x"6f", x"6e", x"6a", 
        x"6d", x"6f", x"6f", x"6e", x"6f", x"6e", x"6a", x"6c", x"6e", x"6e", x"6d", x"6d", x"6d", x"6b", x"6a", 
        x"6b", x"6b", x"6b", x"6d", x"6c", x"6c", x"6c", x"6c", x"6c", x"6c", x"6a", x"6c", x"6e", x"70", x"6e", 
        x"6d", x"6c", x"6c", x"6c", x"6c", x"6b", x"6c", x"6b", x"6d", x"6d", x"6d", x"6e", x"6c", x"6a", x"6c", 
        x"6b", x"6c", x"6c", x"69", x"69", x"6b", x"6b", x"6b", x"6e", x"6e", x"6e", x"71", x"70", x"6d", x"6f", 
        x"6f", x"6f", x"6e", x"6d", x"6b", x"6b", x"6a", x"68", x"6b", x"6b", x"6d", x"6c", x"6a", x"6a", x"6b", 
        x"67", x"69", x"6d", x"68", x"68", x"6b", x"6b", x"69", x"6b", x"6c", x"69", x"65", x"68", x"6c", x"6c", 
        x"69", x"6a", x"6c", x"6b", x"69", x"6a", x"6a", x"67", x"67", x"66", x"68", x"6b", x"6a", x"68", x"68", 
        x"69", x"6b", x"6a", x"67", x"68", x"68", x"6a", x"6a", x"68", x"66", x"62", x"66", x"69", x"6a", x"6a", 
        x"6b", x"69", x"68", x"68", x"69", x"6b", x"6b", x"6a", x"69", x"66", x"66", x"67", x"67", x"66", x"68", 
        x"68", x"68", x"68", x"65", x"65", x"66", x"68", x"69", x"69", x"68", x"69", x"69", x"61", x"65", x"69", 
        x"68", x"67", x"68", x"69", x"6a", x"69", x"68", x"67", x"65", x"64", x"66", x"66", x"64", x"64", x"63", 
        x"65", x"65", x"65", x"64", x"64", x"64", x"63", x"62", x"62", x"63", x"63", x"63", x"63", x"62", x"62", 
        x"63", x"64", x"63", x"62", x"63", x"63", x"62", x"62", x"61", x"62", x"62", x"62", x"64", x"64", x"64", 
        x"64", x"64", x"63", x"65", x"65", x"63", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", 
        x"66", x"67", x"65", x"65", x"66", x"65", x"68", x"67", x"65", x"64", x"65", x"66", x"66", x"65", x"67", 
        x"67", x"65", x"64", x"63", x"65", x"66", x"67", x"66", x"64", x"64", x"64", x"64", x"63", x"63", x"67", 
        x"64", x"63", x"65", x"66", x"64", x"63", x"67", x"66", x"64", x"65", x"65", x"65", x"63", x"65", x"66", 
        x"66", x"65", x"64", x"65", x"67", x"64", x"64", x"66", x"67", x"67", x"67", x"67", x"66", x"66", x"69", 
        x"6a", x"67", x"66", x"67", x"68", x"68", x"68", x"63", x"65", x"67", x"65", x"65", x"66", x"67", x"68", 
        x"69", x"68", x"67", x"67", x"6a", x"67", x"69", x"67", x"64", x"66", x"65", x"65", x"64", x"64", x"66", 
        x"67", x"67", x"68", x"66", x"67", x"6b", x"68", x"65", x"66", x"68", x"67", x"67", x"69", x"6a", x"6b", 
        x"6b", x"6a", x"6a", x"6c", x"6a", x"6c", x"6e", x"6d", x"6d", x"6e", x"69", x"69", x"69", x"6a", x"6a", 
        x"6a", x"6a", x"6b", x"6a", x"69", x"6a", x"6b", x"6b", x"69", x"6a", x"6a", x"6b", x"6a", x"6a", x"6a", 
        x"6b", x"6c", x"6a", x"6b", x"6c", x"6a", x"6c", x"6d", x"6a", x"6a", x"6a", x"6b", x"6b", x"6c", x"6b", 
        x"6a", x"69", x"6a", x"6c", x"6d", x"6e", x"6e", x"6e", x"6e", x"6c", x"6f", x"6f", x"6b", x"68", x"65", 
        x"81", x"b8", x"c2", x"9c", x"9d", x"c3", x"d3", x"ce", x"ca", x"c8", x"c8", x"cc", x"cb", x"ca", x"cb", 
        x"cd", x"ce", x"ce", x"ce", x"ce", x"cd", x"cd", x"ce", x"ce", x"cf", x"ce", x"cd", x"cc", x"cb", x"cb", 
        x"cb", x"cc", x"cc", x"cb", x"cc", x"cc", x"cf", x"cf", x"ce", x"cd", x"cd", x"cf", x"d3", x"d0", x"ac", 
        x"6a", x"5b", x"5d", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"5f", x"60", 
        x"5e", x"5c", x"5b", x"77", x"bc", x"ea", x"f9", x"f6", x"e3", x"b7", x"7c", x"62", x"5b", x"5e", x"5d", 
        x"5c", x"5f", x"60", x"5e", x"5d", x"5d", x"5e", x"5f", x"5f", x"5e", x"5e", x"60", x"5f", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5f", x"5b", x"5c", x"67", x"78", x"94", x"bb", x"d8", x"e8", x"dc", x"b8", x"92", 
        x"71", x"65", x"6d", x"72", x"71", x"74", x"75", x"73", x"73", x"75", x"76", x"73", x"71", x"71", x"72", 
        x"73", x"73", x"72", x"74", x"75", x"73", x"72", x"73", x"74", x"76", x"74", x"73", x"74", x"75", x"74", 
        x"72", x"71", x"72", x"72", x"73", x"74", x"75", x"75", x"73", x"72", x"71", x"71", x"71", x"71", x"71", 
        x"6e", x"6d", x"72", x"74", x"73", x"70", x"6d", x"6f", x"71", x"72", x"73", x"74", x"74", x"72", x"70", 
        x"70", x"73", x"74", x"71", x"6e", x"6e", x"70", x"6e", x"6f", x"71", x"71", x"70", x"6f", x"6f", x"71", 
        x"71", x"71", x"70", x"6f", x"70", x"72", x"70", x"70", x"72", x"72", x"70", x"70", x"6f", x"71", x"72", 
        x"74", x"72", x"70", x"6e", x"6e", x"6f", x"6f", x"71", x"71", x"6e", x"6d", x"6f", x"72", x"6e", x"70", 
        x"6f", x"6e", x"70", x"70", x"6f", x"73", x"73", x"72", x"71", x"71", x"71", x"71", x"70", x"71", x"70", 
        x"70", x"70", x"6f", x"6f", x"6f", x"6f", x"71", x"73", x"71", x"70", x"70", x"70", x"70", x"71", x"71", 
        x"70", x"70", x"71", x"70", x"6e", x"71", x"72", x"70", x"6e", x"6f", x"72", x"74", x"72", x"70", x"70", 
        x"70", x"71", x"71", x"72", x"70", x"72", x"71", x"6d", x"6e", x"6f", x"70", x"71", x"70", x"6f", x"6f", 
        x"6f", x"6f", x"6e", x"6e", x"6e", x"6f", x"70", x"72", x"72", x"71", x"6d", x"6c", x"6f", x"6e", x"6d", 
        x"6f", x"6d", x"71", x"6f", x"6e", x"6f", x"70", x"6f", x"6f", x"71", x"70", x"6f", x"6e", x"6e", x"6e", 
        x"6e", x"6c", x"6e", x"6f", x"6e", x"6e", x"70", x"6f", x"6f", x"70", x"70", x"70", x"6e", x"6e", x"6c", 
        x"6c", x"6c", x"6b", x"6e", x"70", x"6f", x"70", x"71", x"6f", x"6e", x"6c", x"6c", x"6d", x"6e", x"6c", 
        x"6b", x"6e", x"6d", x"6d", x"70", x"72", x"6e", x"6b", x"6d", x"6e", x"6e", x"6c", x"6d", x"6f", x"6d", 
        x"6a", x"6c", x"6c", x"6d", x"6c", x"6b", x"6d", x"6d", x"6b", x"6b", x"6d", x"6e", x"6d", x"6e", x"70", 
        x"6f", x"6e", x"6d", x"6c", x"6c", x"6c", x"6b", x"6b", x"6e", x"6e", x"6d", x"6e", x"6d", x"6b", x"6b", 
        x"6b", x"6b", x"6b", x"6b", x"6b", x"6d", x"6c", x"6d", x"6e", x"6d", x"6c", x"6e", x"6c", x"6c", x"6c", 
        x"6c", x"70", x"6f", x"6d", x"6f", x"6c", x"6a", x"68", x"69", x"6a", x"6a", x"6a", x"6a", x"6a", x"6b", 
        x"6c", x"6b", x"6a", x"6a", x"6a", x"6a", x"68", x"67", x"6a", x"6b", x"68", x"67", x"69", x"6b", x"6c", 
        x"6a", x"6a", x"6a", x"6b", x"6b", x"6a", x"6a", x"69", x"68", x"67", x"68", x"6b", x"6a", x"69", x"68", 
        x"68", x"68", x"68", x"67", x"66", x"66", x"69", x"69", x"68", x"6a", x"65", x"68", x"6a", x"6a", x"6b", 
        x"6b", x"68", x"68", x"67", x"67", x"6a", x"6d", x"6d", x"68", x"67", x"69", x"6a", x"6a", x"68", x"67", 
        x"67", x"68", x"6a", x"69", x"68", x"67", x"68", x"67", x"67", x"68", x"69", x"6a", x"62", x"65", x"68", 
        x"67", x"66", x"66", x"67", x"67", x"68", x"68", x"68", x"66", x"65", x"65", x"65", x"65", x"66", x"66", 
        x"66", x"66", x"65", x"65", x"64", x"63", x"63", x"62", x"62", x"63", x"64", x"64", x"63", x"62", x"62", 
        x"63", x"63", x"63", x"64", x"64", x"65", x"64", x"64", x"64", x"64", x"64", x"63", x"64", x"64", x"64", 
        x"64", x"63", x"62", x"64", x"66", x"65", x"62", x"61", x"62", x"62", x"62", x"61", x"61", x"61", x"61", 
        x"64", x"66", x"64", x"65", x"67", x"66", x"68", x"67", x"65", x"64", x"64", x"65", x"64", x"64", x"66", 
        x"67", x"65", x"64", x"65", x"66", x"65", x"65", x"63", x"63", x"64", x"65", x"66", x"66", x"66", x"69", 
        x"66", x"64", x"64", x"64", x"63", x"63", x"65", x"64", x"65", x"66", x"66", x"66", x"64", x"64", x"65", 
        x"65", x"64", x"65", x"66", x"68", x"69", x"68", x"68", x"67", x"67", x"67", x"64", x"64", x"69", x"69", 
        x"68", x"66", x"66", x"68", x"68", x"67", x"68", x"65", x"68", x"69", x"67", x"66", x"67", x"68", x"68", 
        x"68", x"69", x"67", x"66", x"67", x"65", x"68", x"69", x"66", x"67", x"65", x"68", x"66", x"65", x"68", 
        x"6b", x"6a", x"6a", x"6a", x"69", x"68", x"67", x"65", x"66", x"66", x"67", x"6a", x"6a", x"69", x"69", 
        x"67", x"66", x"68", x"6c", x"6b", x"6b", x"6b", x"69", x"6a", x"6b", x"69", x"68", x"6a", x"6d", x"6c", 
        x"6b", x"6b", x"6a", x"6a", x"6a", x"6a", x"6a", x"6a", x"6a", x"6b", x"6c", x"6c", x"6c", x"6c", x"6c", 
        x"6b", x"6c", x"6b", x"6b", x"6b", x"6b", x"6c", x"6c", x"6c", x"6c", x"6c", x"6c", x"6c", x"6b", x"6b", 
        x"6c", x"6b", x"6a", x"6c", x"6e", x"70", x"6e", x"6e", x"6f", x"6d", x"6c", x"6f", x"66", x"68", x"9b", 
        x"ca", x"b0", x"8d", x"aa", x"ca", x"d4", x"cd", x"cc", x"c8", x"ca", x"cd", x"ca", x"ca", x"cc", x"cf", 
        x"ce", x"ce", x"cf", x"cf", x"ce", x"ce", x"cd", x"cd", x"cd", x"ce", x"ce", x"cd", x"cc", x"cb", x"ca", 
        x"ca", x"cc", x"cc", x"cb", x"cc", x"ce", x"cf", x"cf", x"cd", x"cd", x"ce", x"cf", x"d2", x"d0", x"ae", 
        x"6c", x"5b", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"61", 
        x"5d", x"5e", x"84", x"ca", x"f1", x"f8", x"f7", x"da", x"95", x"67", x"5e", x"5f", x"5c", x"5a", x"5d", 
        x"60", x"5e", x"5d", x"5c", x"5b", x"5b", x"5c", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"5e", 
        x"5d", x"5d", x"5e", x"5f", x"5b", x"5b", x"5f", x"60", x"62", x"70", x"86", x"aa", x"d2", x"e7", x"e4", 
        x"cd", x"a7", x"7a", x"66", x"65", x"6e", x"76", x"74", x"71", x"72", x"74", x"72", x"70", x"70", x"71", 
        x"72", x"72", x"70", x"73", x"76", x"75", x"73", x"73", x"74", x"73", x"72", x"72", x"74", x"75", x"75", 
        x"74", x"72", x"72", x"73", x"73", x"73", x"73", x"72", x"71", x"70", x"6f", x"6f", x"70", x"71", x"70", 
        x"6f", x"6f", x"71", x"73", x"73", x"71", x"6f", x"71", x"74", x"73", x"74", x"75", x"74", x"72", x"72", 
        x"71", x"70", x"72", x"71", x"70", x"71", x"6f", x"71", x"73", x"72", x"72", x"72", x"71", x"72", x"72", 
        x"71", x"70", x"6f", x"6f", x"71", x"73", x"71", x"71", x"73", x"72", x"71", x"72", x"71", x"71", x"73", 
        x"74", x"72", x"71", x"71", x"70", x"70", x"70", x"70", x"6f", x"6f", x"70", x"72", x"72", x"6f", x"70", 
        x"70", x"6f", x"70", x"71", x"70", x"71", x"71", x"6f", x"71", x"71", x"6f", x"70", x"72", x"71", x"71", 
        x"71", x"6f", x"6f", x"6f", x"6e", x"6f", x"72", x"74", x"73", x"72", x"72", x"72", x"70", x"71", x"72", 
        x"70", x"70", x"72", x"70", x"6c", x"70", x"74", x"70", x"6d", x"6f", x"72", x"72", x"70", x"6f", x"71", 
        x"71", x"72", x"73", x"71", x"6d", x"6f", x"73", x"71", x"6e", x"71", x"71", x"71", x"71", x"70", x"70", 
        x"70", x"6f", x"6e", x"6f", x"6f", x"6f", x"6e", x"6e", x"6f", x"6f", x"6d", x"6b", x"6e", x"6e", x"6d", 
        x"6e", x"6f", x"71", x"6f", x"6e", x"6e", x"6f", x"6f", x"6e", x"70", x"70", x"6f", x"6f", x"6f", x"6f", 
        x"6e", x"6d", x"6d", x"6f", x"6f", x"6f", x"70", x"6d", x"6c", x"6e", x"6f", x"70", x"70", x"72", x"70", 
        x"6f", x"6f", x"6d", x"6e", x"70", x"6f", x"70", x"71", x"6d", x"6f", x"6e", x"6c", x"6e", x"70", x"70", 
        x"6c", x"6c", x"6b", x"6a", x"6e", x"6f", x"6d", x"6e", x"6c", x"6b", x"6d", x"6d", x"6d", x"6e", x"6f", 
        x"6e", x"6e", x"6e", x"6b", x"6a", x"69", x"6b", x"6e", x"69", x"67", x"6d", x"6f", x"6f", x"6d", x"6c", 
        x"6c", x"6c", x"6b", x"6c", x"6d", x"6e", x"6c", x"6d", x"71", x"70", x"6f", x"70", x"6e", x"6c", x"6b", 
        x"6b", x"6b", x"6b", x"6e", x"6e", x"6e", x"6d", x"6d", x"6d", x"6b", x"69", x"6c", x"6a", x"6d", x"6a", 
        x"68", x"6c", x"6b", x"68", x"6e", x"6e", x"6b", x"6a", x"68", x"6a", x"68", x"69", x"6a", x"6b", x"6a", 
        x"6f", x"6d", x"67", x"6c", x"6c", x"6a", x"67", x"66", x"6b", x"6d", x"69", x"69", x"6b", x"6b", x"6b", 
        x"6a", x"69", x"68", x"6a", x"6b", x"69", x"67", x"68", x"67", x"66", x"67", x"68", x"68", x"68", x"68", 
        x"68", x"68", x"68", x"69", x"67", x"66", x"6a", x"6a", x"69", x"6f", x"6b", x"6b", x"69", x"67", x"69", 
        x"6a", x"69", x"68", x"67", x"66", x"68", x"6d", x"6d", x"68", x"66", x"66", x"68", x"69", x"6a", x"69", 
        x"6b", x"6b", x"6a", x"6b", x"6b", x"69", x"67", x"66", x"65", x"66", x"67", x"68", x"64", x"66", x"65", 
        x"66", x"64", x"65", x"66", x"66", x"66", x"66", x"66", x"66", x"66", x"65", x"65", x"66", x"66", x"67", 
        x"67", x"67", x"66", x"64", x"64", x"63", x"63", x"65", x"64", x"63", x"63", x"63", x"63", x"64", x"64", 
        x"63", x"63", x"64", x"65", x"65", x"66", x"66", x"65", x"65", x"66", x"66", x"64", x"63", x"62", x"64", 
        x"64", x"61", x"60", x"63", x"67", x"67", x"63", x"62", x"62", x"63", x"63", x"62", x"61", x"61", x"61", 
        x"66", x"65", x"66", x"66", x"66", x"67", x"66", x"68", x"68", x"66", x"65", x"65", x"64", x"63", x"66", 
        x"66", x"65", x"66", x"66", x"65", x"64", x"66", x"67", x"67", x"68", x"67", x"67", x"66", x"64", x"65", 
        x"64", x"64", x"66", x"67", x"67", x"66", x"64", x"64", x"67", x"66", x"65", x"67", x"65", x"65", x"65", 
        x"65", x"66", x"66", x"67", x"67", x"68", x"69", x"68", x"67", x"68", x"6a", x"67", x"67", x"69", x"68", 
        x"67", x"66", x"67", x"69", x"69", x"68", x"69", x"64", x"68", x"68", x"66", x"65", x"68", x"67", x"67", 
        x"67", x"68", x"67", x"66", x"68", x"68", x"67", x"69", x"6a", x"68", x"67", x"68", x"67", x"66", x"69", 
        x"6a", x"69", x"68", x"68", x"65", x"65", x"68", x"68", x"6b", x"6b", x"68", x"69", x"69", x"69", x"69", 
        x"69", x"6a", x"6a", x"6c", x"6c", x"6c", x"6a", x"6a", x"6a", x"69", x"6a", x"69", x"6b", x"6c", x"6b", 
        x"6a", x"6b", x"69", x"69", x"69", x"69", x"6a", x"6a", x"6b", x"6d", x"6c", x"69", x"69", x"6a", x"6c", 
        x"6c", x"6a", x"6c", x"6a", x"69", x"6c", x"6b", x"69", x"6c", x"6b", x"6a", x"6b", x"6b", x"6b", x"6c", 
        x"6d", x"6d", x"6b", x"6e", x"6e", x"70", x"6e", x"71", x"6e", x"6b", x"68", x"66", x"7b", x"ab", x"c1", 
        x"a2", x"97", x"bc", x"cf", x"ce", x"cf", x"cf", x"cc", x"ca", x"cc", x"cd", x"cc", x"cb", x"cb", x"cf", 
        x"ce", x"ce", x"cf", x"cf", x"ce", x"ce", x"cd", x"cd", x"cd", x"cd", x"cd", x"cc", x"cc", x"cb", x"cb", 
        x"ca", x"cc", x"cc", x"ca", x"ca", x"ce", x"cf", x"ce", x"cd", x"ce", x"cf", x"d0", x"d1", x"d0", x"b1", 
        x"6f", x"5b", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"5f", x"63", 
        x"5e", x"80", x"c6", x"f3", x"f8", x"f5", x"d6", x"8a", x"65", x"5c", x"5c", x"5e", x"60", x"5f", x"5b", 
        x"5c", x"60", x"5f", x"5d", x"5d", x"5c", x"5c", x"5e", x"5f", x"5e", x"5d", x"5d", x"5f", x"5f", x"5e", 
        x"5d", x"5d", x"5e", x"5e", x"5d", x"5c", x"5e", x"60", x"5e", x"5d", x"60", x"6a", x"7f", x"a1", x"bf", 
        x"dd", x"e2", x"d3", x"b3", x"85", x"6d", x"6b", x"6e", x"75", x"78", x"74", x"74", x"73", x"73", x"74", 
        x"75", x"74", x"71", x"73", x"74", x"73", x"72", x"72", x"73", x"73", x"73", x"73", x"73", x"72", x"72", 
        x"72", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"72", x"71", x"72", x"73", x"72", x"71", 
        x"71", x"71", x"71", x"71", x"71", x"71", x"71", x"73", x"73", x"71", x"72", x"74", x"74", x"73", x"74", 
        x"71", x"6d", x"6f", x"70", x"72", x"74", x"71", x"71", x"73", x"71", x"72", x"73", x"71", x"72", x"73", 
        x"71", x"70", x"70", x"71", x"73", x"74", x"73", x"73", x"74", x"72", x"73", x"75", x"72", x"72", x"74", 
        x"74", x"72", x"73", x"75", x"73", x"70", x"71", x"70", x"70", x"70", x"71", x"71", x"71", x"6f", x"70", 
        x"70", x"70", x"71", x"71", x"72", x"6f", x"71", x"6e", x"71", x"71", x"6e", x"71", x"72", x"70", x"71", 
        x"71", x"6f", x"70", x"6f", x"6e", x"70", x"72", x"73", x"73", x"71", x"72", x"72", x"70", x"70", x"72", 
        x"6e", x"6f", x"72", x"6f", x"6c", x"6d", x"72", x"70", x"70", x"72", x"72", x"72", x"72", x"71", x"72", 
        x"71", x"71", x"71", x"73", x"71", x"70", x"71", x"6f", x"6c", x"70", x"71", x"72", x"71", x"6f", x"6f", 
        x"70", x"70", x"6f", x"70", x"71", x"70", x"6e", x"6d", x"6e", x"6e", x"6d", x"6d", x"6d", x"6e", x"6e", 
        x"6e", x"6f", x"6f", x"6f", x"6e", x"6e", x"6f", x"6e", x"6e", x"6e", x"6f", x"70", x"71", x"71", x"70", 
        x"6f", x"6f", x"6e", x"70", x"6f", x"6f", x"6e", x"6c", x"6f", x"72", x"71", x"70", x"6d", x"70", x"6e", 
        x"6f", x"71", x"6f", x"6f", x"6f", x"6d", x"6e", x"6f", x"6d", x"6d", x"6c", x"6b", x"6d", x"6f", x"6e", 
        x"6c", x"6c", x"6d", x"6e", x"6d", x"6d", x"6d", x"6f", x"6b", x"6a", x"6c", x"6e", x"6d", x"6e", x"70", 
        x"6d", x"6d", x"6f", x"6b", x"6b", x"6c", x"6d", x"6f", x"6b", x"68", x"6f", x"70", x"6f", x"6e", x"6c", 
        x"6d", x"6d", x"6d", x"6d", x"6f", x"70", x"6b", x"6b", x"6f", x"6e", x"6c", x"6e", x"6c", x"6d", x"6c", 
        x"6e", x"6d", x"6c", x"6e", x"6e", x"6d", x"6b", x"6b", x"6d", x"6d", x"6c", x"6f", x"6d", x"6f", x"6d", 
        x"6d", x"6f", x"6f", x"6c", x"70", x"6e", x"6d", x"6d", x"6a", x"6c", x"69", x"6b", x"6a", x"6a", x"68", 
        x"6a", x"69", x"68", x"6b", x"6a", x"6a", x"68", x"67", x"6b", x"6c", x"69", x"68", x"6a", x"6b", x"6a", 
        x"68", x"68", x"69", x"6b", x"6c", x"69", x"67", x"69", x"68", x"66", x"68", x"67", x"66", x"67", x"69", 
        x"6a", x"69", x"68", x"69", x"69", x"68", x"6c", x"69", x"67", x"6d", x"6b", x"6b", x"6a", x"67", x"68", 
        x"69", x"68", x"65", x"68", x"69", x"68", x"68", x"6a", x"69", x"69", x"68", x"6a", x"69", x"69", x"66", 
        x"6a", x"68", x"67", x"6a", x"6a", x"6a", x"68", x"68", x"66", x"67", x"65", x"63", x"64", x"65", x"62", 
        x"66", x"68", x"69", x"6a", x"68", x"68", x"69", x"6a", x"67", x"69", x"68", x"66", x"65", x"63", x"66", 
        x"67", x"69", x"68", x"66", x"67", x"64", x"65", x"67", x"65", x"63", x"62", x"62", x"63", x"64", x"64", 
        x"63", x"63", x"64", x"65", x"66", x"66", x"66", x"66", x"66", x"66", x"66", x"65", x"64", x"63", x"64", 
        x"65", x"62", x"62", x"64", x"68", x"68", x"64", x"62", x"62", x"63", x"64", x"63", x"61", x"63", x"63", 
        x"69", x"66", x"68", x"68", x"66", x"67", x"65", x"69", x"6a", x"68", x"66", x"66", x"65", x"63", x"65", 
        x"67", x"66", x"67", x"67", x"66", x"65", x"66", x"66", x"66", x"68", x"66", x"66", x"66", x"64", x"64", 
        x"65", x"66", x"67", x"67", x"67", x"66", x"65", x"65", x"69", x"66", x"64", x"66", x"65", x"67", x"66", 
        x"65", x"67", x"67", x"67", x"66", x"66", x"6a", x"6b", x"68", x"66", x"67", x"68", x"68", x"69", x"68", 
        x"67", x"67", x"68", x"68", x"67", x"68", x"68", x"63", x"67", x"66", x"65", x"65", x"68", x"67", x"66", 
        x"66", x"67", x"66", x"66", x"69", x"6a", x"66", x"67", x"68", x"66", x"65", x"68", x"69", x"69", x"6c", 
        x"6b", x"68", x"68", x"68", x"66", x"68", x"6a", x"69", x"6a", x"6c", x"6a", x"69", x"69", x"68", x"68", 
        x"68", x"69", x"69", x"69", x"6b", x"6a", x"6a", x"6a", x"68", x"66", x"6d", x"6b", x"6b", x"6b", x"6a", 
        x"69", x"6c", x"6a", x"67", x"66", x"69", x"6c", x"6c", x"6a", x"6c", x"6c", x"6b", x"6c", x"6e", x"6e", 
        x"6b", x"6a", x"6f", x"6d", x"6b", x"6f", x"6d", x"6b", x"6e", x"6c", x"6c", x"6d", x"6e", x"70", x"71", 
        x"71", x"6e", x"6d", x"70", x"6e", x"6f", x"6e", x"73", x"6d", x"69", x"62", x"86", x"bf", x"c6", x"91", 
        x"9f", x"ca", x"cb", x"cc", x"ce", x"cc", x"cf", x"cf", x"cc", x"cc", x"cd", x"ce", x"cf", x"cf", x"cd", 
        x"cd", x"ce", x"cf", x"cf", x"ce", x"ce", x"ce", x"cd", x"cc", x"cc", x"cc", x"cc", x"cb", x"cb", x"cc", 
        x"cc", x"cd", x"cc", x"ca", x"c9", x"cc", x"ce", x"ce", x"ce", x"cf", x"d0", x"d1", x"d1", x"d0", x"b3", 
        x"71", x"5c", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5d", x"5c", x"5d", x"60", 
        x"71", x"c0", x"f2", x"f6", x"f4", x"da", x"99", x"5e", x"5d", x"5e", x"5b", x"5d", x"5c", x"5c", x"5f", 
        x"5f", x"5d", x"5c", x"5e", x"5f", x"5d", x"5d", x"5e", x"5f", x"5e", x"5d", x"5d", x"5e", x"5f", x"5f", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"5f", x"5d", x"5a", x"5a", x"60", x"5e", x"65", x"76", 
        x"96", x"bc", x"d9", x"e9", x"de", x"be", x"8f", x"68", x"65", x"6e", x"74", x"75", x"74", x"74", x"74", 
        x"75", x"76", x"74", x"74", x"75", x"74", x"73", x"74", x"74", x"71", x"72", x"73", x"73", x"71", x"72", 
        x"74", x"75", x"74", x"73", x"73", x"74", x"76", x"77", x"73", x"72", x"73", x"74", x"74", x"72", x"6f", 
        x"71", x"72", x"72", x"71", x"71", x"72", x"72", x"74", x"73", x"70", x"71", x"72", x"72", x"72", x"73", 
        x"72", x"70", x"70", x"6e", x"6e", x"71", x"6f", x"6f", x"72", x"71", x"73", x"74", x"70", x"70", x"73", 
        x"71", x"70", x"71", x"73", x"75", x"75", x"74", x"74", x"74", x"71", x"73", x"76", x"73", x"73", x"73", 
        x"72", x"71", x"72", x"75", x"72", x"6f", x"70", x"72", x"71", x"70", x"6e", x"6f", x"71", x"71", x"70", 
        x"71", x"72", x"70", x"70", x"72", x"6f", x"72", x"70", x"73", x"72", x"6f", x"74", x"74", x"71", x"72", 
        x"72", x"6f", x"71", x"70", x"70", x"72", x"73", x"73", x"70", x"6f", x"6f", x"70", x"71", x"70", x"72", 
        x"6e", x"6e", x"72", x"71", x"72", x"70", x"72", x"72", x"72", x"72", x"6e", x"70", x"71", x"72", x"72", 
        x"72", x"71", x"71", x"72", x"72", x"70", x"6e", x"6d", x"6e", x"71", x"71", x"71", x"71", x"6e", x"6e", 
        x"70", x"71", x"6f", x"6f", x"71", x"71", x"6f", x"6e", x"70", x"70", x"6e", x"6f", x"6c", x"6e", x"71", 
        x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"6e", x"6e", x"6e", x"6f", x"71", x"72", x"70", 
        x"6f", x"70", x"6d", x"6f", x"6f", x"70", x"6f", x"6e", x"6f", x"70", x"6f", x"6e", x"6c", x"70", x"70", 
        x"70", x"70", x"6d", x"6e", x"6f", x"6e", x"6f", x"71", x"71", x"6e", x"6c", x"6d", x"70", x"6f", x"6d", 
        x"6d", x"6c", x"70", x"73", x"70", x"6f", x"71", x"6d", x"6b", x"6a", x"6c", x"6d", x"6d", x"70", x"6f", 
        x"69", x"6a", x"6d", x"6c", x"6e", x"71", x"6f", x"6c", x"6d", x"69", x"6d", x"6a", x"6a", x"6b", x"6c", 
        x"6d", x"6d", x"6c", x"6c", x"6e", x"6e", x"6b", x"6b", x"6f", x"6d", x"6b", x"6d", x"6c", x"6e", x"6d", 
        x"70", x"70", x"6e", x"6f", x"6d", x"6d", x"6c", x"6c", x"6e", x"6f", x"6f", x"70", x"71", x"71", x"70", 
        x"73", x"6f", x"6f", x"6c", x"6c", x"6d", x"6d", x"6e", x"6b", x"6d", x"6a", x"6e", x"6e", x"6c", x"6b", 
        x"67", x"69", x"6e", x"6a", x"68", x"6a", x"6a", x"68", x"69", x"6a", x"68", x"66", x"69", x"6c", x"6a", 
        x"67", x"67", x"6a", x"6c", x"6d", x"6a", x"69", x"6b", x"6a", x"68", x"6b", x"6b", x"67", x"67", x"69", 
        x"6a", x"69", x"69", x"6c", x"68", x"65", x"67", x"65", x"64", x"6b", x"67", x"6a", x"6b", x"69", x"69", 
        x"68", x"66", x"67", x"69", x"67", x"66", x"69", x"6a", x"67", x"68", x"68", x"69", x"68", x"67", x"64", 
        x"69", x"69", x"6a", x"6b", x"6a", x"68", x"66", x"66", x"67", x"6a", x"66", x"63", x"67", x"69", x"64", 
        x"6a", x"68", x"68", x"66", x"63", x"63", x"66", x"6a", x"66", x"69", x"69", x"68", x"67", x"64", x"66", 
        x"68", x"6b", x"69", x"67", x"68", x"65", x"67", x"67", x"64", x"64", x"64", x"64", x"64", x"64", x"64", 
        x"65", x"65", x"65", x"65", x"65", x"65", x"65", x"66", x"66", x"65", x"65", x"65", x"66", x"66", x"65", 
        x"66", x"65", x"65", x"66", x"69", x"68", x"65", x"63", x"62", x"63", x"65", x"65", x"62", x"65", x"64", 
        x"6c", x"65", x"67", x"66", x"64", x"69", x"66", x"67", x"69", x"68", x"67", x"64", x"64", x"66", x"67", 
        x"68", x"68", x"66", x"66", x"66", x"67", x"69", x"68", x"65", x"65", x"63", x"66", x"67", x"67", x"64", 
        x"66", x"67", x"65", x"67", x"6a", x"66", x"65", x"67", x"67", x"66", x"68", x"6a", x"68", x"66", x"64", 
        x"65", x"66", x"66", x"66", x"68", x"65", x"65", x"67", x"68", x"67", x"66", x"67", x"68", x"69", x"68", 
        x"65", x"64", x"65", x"65", x"66", x"69", x"66", x"65", x"6b", x"6a", x"66", x"68", x"69", x"6a", x"66", 
        x"66", x"67", x"66", x"69", x"69", x"6a", x"69", x"69", x"66", x"6a", x"6b", x"6b", x"6c", x"69", x"68", 
        x"6a", x"65", x"67", x"69", x"68", x"69", x"68", x"6a", x"69", x"68", x"69", x"6b", x"6a", x"68", x"67", 
        x"68", x"6b", x"6d", x"6c", x"6c", x"6a", x"69", x"6c", x"6b", x"69", x"6c", x"6c", x"6c", x"6a", x"6d", 
        x"6d", x"6d", x"6b", x"6b", x"6c", x"6e", x"6d", x"6c", x"6a", x"6b", x"6b", x"6b", x"6d", x"6e", x"6b", 
        x"65", x"67", x"6c", x"6c", x"6c", x"6c", x"6c", x"6b", x"6c", x"70", x"6f", x"6b", x"70", x"71", x"72", 
        x"70", x"70", x"71", x"70", x"6e", x"6d", x"6d", x"6d", x"6b", x"6e", x"99", x"c6", x"b3", x"8f", x"b0", 
        x"cc", x"d2", x"cd", x"cd", x"ce", x"cd", x"ce", x"ce", x"cd", x"cc", x"cd", x"ce", x"cf", x"cf", x"cd", 
        x"cd", x"cf", x"d0", x"cf", x"ce", x"ce", x"ce", x"cd", x"cd", x"cd", x"cd", x"cd", x"cb", x"ca", x"cc", 
        x"ce", x"cd", x"cb", x"cb", x"cc", x"cb", x"cd", x"d2", x"ce", x"d1", x"d0", x"d0", x"d0", x"ce", x"b5", 
        x"73", x"5d", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"5e", x"5d", x"67", 
        x"a3", x"ed", x"f8", x"f8", x"db", x"93", x"63", x"5d", x"5e", x"5c", x"5d", x"5f", x"5d", x"5d", x"5e", 
        x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", 
        x"5d", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5d", x"5c", x"5d", x"5f", x"60", x"5e", x"5e", 
        x"65", x"72", x"8a", x"ae", x"d2", x"e3", x"e2", x"c5", x"99", x"74", x"69", x"6f", x"74", x"75", x"75", 
        x"73", x"72", x"6f", x"6f", x"70", x"75", x"74", x"73", x"73", x"72", x"72", x"75", x"75", x"73", x"72", 
        x"75", x"75", x"74", x"73", x"73", x"73", x"73", x"74", x"72", x"72", x"74", x"76", x"75", x"72", x"73", 
        x"70", x"72", x"75", x"75", x"75", x"72", x"71", x"72", x"72", x"73", x"73", x"73", x"73", x"73", x"73", 
        x"71", x"73", x"70", x"70", x"72", x"71", x"72", x"71", x"6e", x"6f", x"73", x"72", x"71", x"72", x"72", 
        x"6e", x"72", x"72", x"71", x"73", x"74", x"71", x"70", x"6f", x"6f", x"71", x"72", x"73", x"72", x"72", 
        x"74", x"74", x"72", x"71", x"73", x"73", x"72", x"6f", x"6e", x"71", x"71", x"73", x"71", x"73", x"73", 
        x"72", x"72", x"72", x"72", x"72", x"6f", x"72", x"73", x"72", x"72", x"73", x"73", x"71", x"72", x"72", 
        x"71", x"71", x"70", x"71", x"75", x"71", x"73", x"76", x"6e", x"6f", x"71", x"6e", x"74", x"73", x"73", 
        x"72", x"71", x"71", x"71", x"73", x"73", x"74", x"73", x"73", x"71", x"6f", x"71", x"70", x"6f", x"6f", 
        x"71", x"71", x"71", x"6f", x"70", x"70", x"70", x"70", x"70", x"73", x"70", x"70", x"70", x"6d", x"6e", 
        x"71", x"72", x"71", x"72", x"72", x"72", x"70", x"6f", x"6f", x"70", x"70", x"6f", x"70", x"70", x"71", 
        x"6f", x"71", x"70", x"71", x"71", x"73", x"73", x"72", x"72", x"73", x"71", x"6e", x"6e", x"6f", x"6e", 
        x"6c", x"70", x"71", x"70", x"71", x"72", x"71", x"6f", x"6f", x"6d", x"6c", x"6d", x"6b", x"6e", x"6f", 
        x"6e", x"70", x"6f", x"70", x"71", x"6e", x"6d", x"70", x"72", x"71", x"70", x"70", x"70", x"6f", x"6d", 
        x"6d", x"6b", x"6e", x"6e", x"6f", x"74", x"71", x"72", x"73", x"6f", x"6e", x"70", x"71", x"6d", x"6c", 
        x"6c", x"6d", x"6d", x"6d", x"6d", x"6f", x"6f", x"6e", x"70", x"6e", x"6c", x"6d", x"6f", x"6f", x"6d", 
        x"6c", x"70", x"6e", x"6d", x"6e", x"6d", x"6f", x"6d", x"6d", x"6d", x"6d", x"71", x"6f", x"6f", x"6e", 
        x"6e", x"6f", x"70", x"6f", x"6e", x"6d", x"6d", x"6c", x"6c", x"6e", x"70", x"6f", x"6e", x"6d", x"6f", 
        x"6f", x"6e", x"6e", x"6b", x"6d", x"6d", x"6d", x"6d", x"6a", x"6b", x"6e", x"6f", x"6e", x"6c", x"6d", 
        x"68", x"69", x"6c", x"69", x"6a", x"6c", x"6d", x"6c", x"69", x"69", x"69", x"68", x"69", x"6a", x"6a", 
        x"6c", x"6b", x"68", x"66", x"69", x"6b", x"6b", x"6c", x"6b", x"68", x"6a", x"6b", x"67", x"6b", x"6e", 
        x"6a", x"67", x"6a", x"6e", x"6a", x"6a", x"69", x"69", x"6b", x"6a", x"67", x"6a", x"6a", x"6a", x"69", 
        x"67", x"69", x"69", x"6a", x"68", x"69", x"68", x"68", x"68", x"67", x"68", x"69", x"6a", x"66", x"66", 
        x"6b", x"69", x"6b", x"6b", x"68", x"65", x"67", x"6a", x"6b", x"69", x"68", x"69", x"6b", x"6c", x"6a", 
        x"69", x"67", x"66", x"67", x"67", x"65", x"66", x"6a", x"68", x"68", x"68", x"69", x"68", x"66", x"67", 
        x"67", x"67", x"67", x"66", x"66", x"65", x"67", x"67", x"66", x"67", x"67", x"66", x"65", x"66", x"66", 
        x"65", x"66", x"67", x"67", x"67", x"66", x"65", x"64", x"65", x"65", x"65", x"65", x"66", x"67", x"64", 
        x"65", x"64", x"64", x"67", x"66", x"63", x"64", x"64", x"64", x"64", x"68", x"6a", x"66", x"65", x"64", 
        x"6b", x"67", x"6a", x"6a", x"68", x"6b", x"67", x"66", x"67", x"68", x"65", x"64", x"64", x"66", x"67", 
        x"65", x"67", x"6c", x"66", x"65", x"68", x"67", x"65", x"63", x"64", x"65", x"68", x"67", x"67", x"66", 
        x"67", x"68", x"66", x"67", x"69", x"65", x"67", x"68", x"67", x"66", x"66", x"67", x"65", x"65", x"64", 
        x"65", x"66", x"66", x"66", x"68", x"66", x"65", x"65", x"66", x"67", x"68", x"69", x"67", x"66", x"68", 
        x"67", x"64", x"64", x"65", x"6a", x"6b", x"67", x"68", x"6a", x"6c", x"6d", x"6a", x"6a", x"6c", x"6a", 
        x"6a", x"68", x"66", x"68", x"6a", x"69", x"69", x"69", x"66", x"6a", x"6b", x"6b", x"6a", x"68", x"68", 
        x"6d", x"6b", x"6a", x"68", x"68", x"6a", x"69", x"69", x"67", x"67", x"6b", x"6c", x"6a", x"69", x"68", 
        x"69", x"6a", x"6c", x"6d", x"6f", x"6e", x"6b", x"6c", x"6c", x"6b", x"6c", x"6c", x"6c", x"69", x"6d", 
        x"6c", x"6b", x"6b", x"6b", x"6c", x"6c", x"6a", x"6a", x"6c", x"6d", x"6d", x"6d", x"6b", x"6a", x"69", 
        x"6c", x"6c", x"6c", x"6b", x"6b", x"6b", x"6c", x"6c", x"6c", x"6f", x"6d", x"6b", x"6f", x"6d", x"6d", 
        x"6d", x"6f", x"6d", x"74", x"70", x"6b", x"6b", x"67", x"7d", x"b1", x"ce", x"a1", x"92", x"be", x"d1", 
        x"cf", x"cd", x"cc", x"ca", x"cb", x"cc", x"cb", x"cd", x"cd", x"cd", x"cd", x"cf", x"cf", x"cf", x"ce", 
        x"ce", x"cf", x"cf", x"cf", x"ce", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"cc", x"ca", x"cd", 
        x"ce", x"cc", x"cb", x"cc", x"cd", x"ca", x"cb", x"d1", x"cd", x"d1", x"d1", x"d1", x"d2", x"ce", x"b6", 
        x"74", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5c", x"58", x"82", 
        x"d8", x"f9", x"f8", x"ef", x"9d", x"62", x"5a", x"61", x"61", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"60", x"5e", x"5d", 
        x"5f", x"62", x"5f", x"66", x"7e", x"9d", x"c4", x"e3", x"ea", x"da", x"a5", x"7b", x"6b", x"6d", x"6f", 
        x"72", x"75", x"75", x"77", x"6e", x"76", x"79", x"75", x"77", x"78", x"76", x"76", x"77", x"75", x"73", 
        x"75", x"75", x"74", x"73", x"72", x"72", x"73", x"74", x"76", x"74", x"73", x"73", x"73", x"73", x"76", 
        x"76", x"75", x"72", x"70", x"73", x"72", x"72", x"73", x"72", x"73", x"73", x"73", x"73", x"74", x"73", 
        x"72", x"74", x"70", x"71", x"73", x"71", x"71", x"72", x"6f", x"71", x"73", x"73", x"72", x"73", x"74", 
        x"71", x"74", x"73", x"73", x"74", x"76", x"74", x"75", x"75", x"74", x"73", x"73", x"76", x"73", x"70", 
        x"71", x"71", x"70", x"70", x"72", x"73", x"74", x"71", x"70", x"73", x"72", x"74", x"72", x"75", x"76", 
        x"75", x"72", x"6f", x"71", x"74", x"71", x"72", x"72", x"70", x"70", x"70", x"6e", x"6d", x"70", x"71", 
        x"70", x"70", x"6f", x"72", x"76", x"72", x"72", x"75", x"6f", x"71", x"72", x"6f", x"74", x"75", x"75", 
        x"73", x"73", x"73", x"72", x"70", x"72", x"70", x"6f", x"70", x"71", x"71", x"71", x"70", x"6e", x"6e", 
        x"70", x"71", x"70", x"6f", x"6f", x"71", x"72", x"72", x"72", x"73", x"70", x"70", x"72", x"71", x"72", 
        x"74", x"74", x"72", x"71", x"71", x"71", x"71", x"70", x"6f", x"71", x"71", x"70", x"70", x"6e", x"6e", 
        x"6b", x"6e", x"6f", x"70", x"70", x"72", x"74", x"73", x"72", x"70", x"71", x"71", x"72", x"71", x"70", 
        x"6f", x"72", x"71", x"70", x"70", x"70", x"70", x"6f", x"6e", x"6d", x"6e", x"70", x"6e", x"70", x"70", 
        x"6e", x"6f", x"6e", x"70", x"71", x"6f", x"6e", x"70", x"6f", x"6e", x"6e", x"6f", x"70", x"6f", x"6e", 
        x"6d", x"6e", x"70", x"6d", x"6c", x"70", x"70", x"70", x"70", x"6f", x"6d", x"6d", x"6d", x"6d", x"6e", 
        x"6f", x"6f", x"6f", x"6e", x"70", x"72", x"72", x"6f", x"6f", x"6e", x"6f", x"73", x"71", x"6e", x"6b", 
        x"6a", x"71", x"71", x"6e", x"6f", x"70", x"70", x"6d", x"6d", x"6c", x"6c", x"70", x"6e", x"6e", x"6d", 
        x"6d", x"6d", x"6e", x"6e", x"6d", x"6e", x"6f", x"70", x"6f", x"6f", x"6e", x"6b", x"6c", x"6d", x"6d", 
        x"6c", x"6d", x"6e", x"6c", x"6d", x"6c", x"6c", x"6d", x"6d", x"6c", x"6d", x"6e", x"70", x"6e", x"6e", 
        x"6b", x"6c", x"6c", x"6d", x"6a", x"69", x"69", x"6c", x"6e", x"6d", x"6a", x"69", x"6a", x"6b", x"6b", 
        x"6d", x"6c", x"67", x"68", x"6a", x"69", x"6b", x"6c", x"6b", x"6a", x"6b", x"6b", x"69", x"6c", x"6d", 
        x"6a", x"68", x"6a", x"6d", x"6b", x"6c", x"6b", x"6a", x"6a", x"66", x"67", x"6a", x"6a", x"6a", x"6a", 
        x"67", x"68", x"65", x"66", x"65", x"68", x"67", x"69", x"6a", x"68", x"69", x"67", x"6a", x"69", x"68", 
        x"68", x"65", x"66", x"68", x"67", x"66", x"67", x"68", x"69", x"69", x"68", x"68", x"69", x"6a", x"69", 
        x"68", x"6a", x"69", x"69", x"69", x"67", x"67", x"69", x"66", x"66", x"68", x"67", x"66", x"65", x"66", 
        x"68", x"69", x"69", x"68", x"67", x"67", x"68", x"66", x"64", x"64", x"65", x"66", x"66", x"67", x"68", 
        x"68", x"67", x"66", x"66", x"66", x"66", x"65", x"64", x"65", x"65", x"65", x"65", x"66", x"67", x"68", 
        x"66", x"65", x"65", x"64", x"63", x"63", x"63", x"63", x"62", x"64", x"68", x"6b", x"69", x"65", x"63", 
        x"69", x"66", x"69", x"6b", x"69", x"6b", x"67", x"67", x"67", x"66", x"65", x"64", x"65", x"65", x"65", 
        x"61", x"67", x"6c", x"67", x"67", x"69", x"66", x"66", x"63", x"66", x"68", x"6a", x"68", x"66", x"65", 
        x"66", x"68", x"67", x"68", x"6a", x"67", x"67", x"67", x"67", x"65", x"65", x"66", x"65", x"65", x"64", 
        x"65", x"66", x"65", x"65", x"68", x"65", x"63", x"67", x"69", x"6a", x"6a", x"68", x"65", x"65", x"67", 
        x"68", x"65", x"64", x"67", x"6a", x"67", x"66", x"67", x"67", x"6b", x"6d", x"65", x"68", x"6b", x"6a", 
        x"6a", x"69", x"67", x"69", x"6c", x"6a", x"69", x"6a", x"68", x"6b", x"6a", x"6a", x"68", x"69", x"69", 
        x"69", x"6b", x"6b", x"67", x"67", x"69", x"6a", x"69", x"67", x"69", x"6d", x"6c", x"6a", x"6a", x"6a", 
        x"6a", x"69", x"68", x"68", x"6d", x"6d", x"6b", x"6c", x"6d", x"6d", x"6c", x"6b", x"6b", x"69", x"6b", 
        x"6b", x"69", x"6e", x"6e", x"6e", x"6c", x"68", x"67", x"6c", x"6c", x"6b", x"6b", x"6a", x"69", x"6a", 
        x"6d", x"6d", x"6c", x"6b", x"6a", x"6b", x"6c", x"6c", x"6d", x"6e", x"6e", x"6e", x"70", x"6e", x"6c", 
        x"6e", x"72", x"72", x"70", x"70", x"68", x"67", x"90", x"c0", x"b6", x"96", x"a4", x"c9", x"d3", x"cb", 
        x"c9", x"cc", x"cd", x"ca", x"ca", x"cc", x"cb", x"cd", x"ce", x"ce", x"ce", x"cf", x"d0", x"cf", x"cf", 
        x"cf", x"cf", x"ce", x"cf", x"ce", x"cd", x"cc", x"cd", x"cc", x"cc", x"cc", x"cc", x"cc", x"cb", x"cc", 
        x"cd", x"cb", x"cb", x"cb", x"cc", x"ca", x"ca", x"cf", x"cb", x"d0", x"d1", x"d2", x"d3", x"cf", x"b7", 
        x"76", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5b", x"66", x"ad", 
        x"f3", x"f9", x"f5", x"c9", x"74", x"59", x"60", x"60", x"5f", x"60", x"5d", x"5d", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", 
        x"5e", x"60", x"60", x"5d", x"5f", x"67", x"78", x"94", x"b1", x"cb", x"e2", x"d7", x"b5", x"8d", x"72", 
        x"6d", x"70", x"72", x"76", x"74", x"75", x"74", x"74", x"76", x"74", x"74", x"75", x"75", x"74", x"73", 
        x"74", x"73", x"73", x"74", x"74", x"74", x"74", x"74", x"75", x"73", x"72", x"74", x"75", x"73", x"74", 
        x"72", x"73", x"71", x"6f", x"72", x"72", x"75", x"76", x"74", x"73", x"73", x"74", x"75", x"75", x"73", 
        x"71", x"73", x"71", x"71", x"73", x"72", x"72", x"70", x"70", x"72", x"72", x"71", x"71", x"73", x"74", 
        x"72", x"74", x"72", x"73", x"74", x"75", x"73", x"74", x"75", x"73", x"70", x"70", x"75", x"74", x"71", 
        x"70", x"70", x"71", x"72", x"74", x"74", x"74", x"73", x"72", x"72", x"71", x"71", x"70", x"71", x"72", 
        x"71", x"6f", x"6f", x"71", x"73", x"71", x"72", x"71", x"71", x"72", x"72", x"6f", x"6f", x"74", x"74", 
        x"72", x"72", x"70", x"72", x"75", x"73", x"73", x"74", x"72", x"73", x"73", x"71", x"71", x"72", x"72", 
        x"71", x"71", x"71", x"72", x"71", x"74", x"73", x"70", x"70", x"71", x"71", x"74", x"72", x"70", x"71", 
        x"72", x"72", x"72", x"70", x"70", x"71", x"72", x"73", x"73", x"72", x"6f", x"6f", x"72", x"73", x"74", 
        x"75", x"74", x"72", x"71", x"71", x"71", x"71", x"70", x"70", x"71", x"71", x"6f", x"71", x"70", x"70", 
        x"6e", x"70", x"70", x"6f", x"6f", x"71", x"73", x"73", x"71", x"6e", x"6f", x"71", x"71", x"6f", x"6d", 
        x"6d", x"72", x"73", x"72", x"71", x"70", x"71", x"70", x"6f", x"6d", x"6f", x"70", x"6f", x"6e", x"6f", 
        x"6f", x"6f", x"6f", x"71", x"71", x"6f", x"6e", x"6e", x"6e", x"6e", x"6f", x"70", x"72", x"72", x"70", 
        x"6f", x"6f", x"6f", x"6d", x"6c", x"6d", x"6d", x"6e", x"6e", x"6f", x"6f", x"6e", x"6d", x"70", x"70", 
        x"6f", x"6f", x"6e", x"6d", x"6d", x"6f", x"70", x"71", x"70", x"6e", x"6e", x"72", x"72", x"6f", x"6d", 
        x"6d", x"72", x"72", x"6d", x"6e", x"71", x"70", x"6d", x"6d", x"6c", x"6c", x"6e", x"6d", x"6d", x"6d", 
        x"6c", x"6d", x"6e", x"6d", x"6d", x"6d", x"6e", x"6d", x"6c", x"6e", x"70", x"6f", x"70", x"6f", x"6d", 
        x"6c", x"6d", x"6f", x"6d", x"6d", x"6d", x"6d", x"6c", x"6e", x"6e", x"6d", x"6e", x"70", x"6e", x"6d", 
        x"6c", x"6d", x"6c", x"6f", x"6c", x"6a", x"6a", x"6b", x"6d", x"6c", x"69", x"6b", x"6c", x"6c", x"6b", 
        x"6c", x"6c", x"68", x"6a", x"6b", x"69", x"6b", x"6d", x"6b", x"6a", x"6c", x"6c", x"6c", x"6b", x"6b", 
        x"69", x"69", x"6a", x"6c", x"6b", x"6c", x"6b", x"6b", x"69", x"66", x"67", x"6a", x"69", x"69", x"69", 
        x"67", x"68", x"6c", x"6d", x"6b", x"6c", x"6b", x"6b", x"6c", x"6a", x"6b", x"67", x"69", x"6c", x"69", 
        x"67", x"65", x"65", x"68", x"6b", x"6b", x"69", x"68", x"69", x"6a", x"69", x"68", x"68", x"68", x"67", 
        x"67", x"69", x"69", x"6a", x"6a", x"69", x"69", x"6a", x"66", x"68", x"6a", x"67", x"66", x"67", x"67", 
        x"67", x"68", x"68", x"67", x"67", x"67", x"69", x"68", x"66", x"65", x"66", x"67", x"68", x"67", x"68", 
        x"68", x"67", x"66", x"66", x"66", x"66", x"66", x"66", x"67", x"67", x"67", x"67", x"67", x"68", x"67", 
        x"66", x"67", x"67", x"65", x"64", x"64", x"63", x"63", x"63", x"64", x"67", x"68", x"66", x"64", x"63", 
        x"69", x"67", x"69", x"69", x"68", x"69", x"65", x"68", x"68", x"67", x"65", x"65", x"66", x"66", x"6a", 
        x"6f", x"71", x"6e", x"68", x"68", x"66", x"64", x"66", x"63", x"64", x"67", x"69", x"67", x"65", x"65", 
        x"66", x"67", x"68", x"69", x"69", x"68", x"65", x"65", x"66", x"66", x"67", x"68", x"68", x"66", x"65", 
        x"66", x"66", x"65", x"64", x"68", x"66", x"65", x"67", x"69", x"6b", x"6a", x"68", x"68", x"67", x"66", 
        x"67", x"67", x"66", x"68", x"68", x"66", x"69", x"68", x"68", x"6d", x"6a", x"64", x"67", x"69", x"68", 
        x"67", x"67", x"69", x"6b", x"6e", x"6b", x"6b", x"6b", x"6a", x"6c", x"6a", x"68", x"66", x"69", x"68", 
        x"64", x"6a", x"6d", x"6a", x"67", x"67", x"6a", x"6a", x"68", x"6a", x"6c", x"6c", x"6a", x"6a", x"6c", 
        x"6b", x"69", x"67", x"66", x"6a", x"6b", x"6b", x"6c", x"6c", x"6a", x"68", x"69", x"6a", x"6a", x"6d", 
        x"6e", x"6c", x"6e", x"6f", x"70", x"6f", x"6a", x"69", x"6f", x"6b", x"68", x"6a", x"6c", x"6d", x"6d", 
        x"6b", x"6c", x"6d", x"6c", x"6a", x"6b", x"6d", x"6d", x"6d", x"6e", x"6d", x"6e", x"6f", x"6e", x"6c", 
        x"6e", x"6a", x"6c", x"6d", x"69", x"74", x"99", x"c6", x"b0", x"94", x"aa", x"d1", x"d2", x"c8", x"ca", 
        x"cd", x"ce", x"ce", x"cc", x"cb", x"cb", x"cd", x"cf", x"cf", x"ce", x"ce", x"d0", x"d0", x"cf", x"ce", 
        x"ce", x"cd", x"ce", x"cf", x"d0", x"ce", x"cc", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"cc", 
        x"cc", x"cb", x"cb", x"cb", x"cc", x"ca", x"ca", x"cf", x"cb", x"cf", x"d0", x"d1", x"d2", x"cf", x"b8", 
        x"78", x"5e", x"5d", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5c", x"7f", x"d6", 
        x"fa", x"f9", x"ee", x"a0", x"62", x"5c", x"60", x"5c", x"5e", x"60", x"5f", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5d", x"5d", x"5e", x"5c", x"59", x"58", x"5e", x"77", x"a8", x"cc", x"e8", x"e0", x"ba", 
        x"95", x"74", x"6a", x"6e", x"74", x"71", x"74", x"79", x"76", x"77", x"78", x"77", x"74", x"72", x"73", 
        x"75", x"73", x"73", x"75", x"75", x"75", x"75", x"75", x"75", x"73", x"72", x"75", x"76", x"74", x"73", 
        x"70", x"73", x"75", x"73", x"73", x"71", x"73", x"76", x"74", x"73", x"73", x"75", x"76", x"75", x"72", 
        x"70", x"72", x"71", x"71", x"73", x"74", x"73", x"72", x"73", x"74", x"73", x"72", x"72", x"73", x"73", 
        x"71", x"73", x"72", x"74", x"73", x"73", x"71", x"72", x"72", x"70", x"6f", x"70", x"73", x"75", x"74", 
        x"72", x"71", x"73", x"74", x"75", x"74", x"72", x"73", x"74", x"75", x"75", x"75", x"75", x"75", x"73", 
        x"71", x"71", x"72", x"71", x"70", x"75", x"75", x"74", x"74", x"74", x"72", x"6f", x"6f", x"71", x"6f", 
        x"70", x"74", x"73", x"72", x"74", x"74", x"73", x"73", x"74", x"74", x"74", x"72", x"70", x"72", x"72", 
        x"71", x"71", x"72", x"72", x"6f", x"73", x"74", x"71", x"70", x"71", x"71", x"74", x"72", x"70", x"70", 
        x"71", x"72", x"72", x"70", x"6f", x"70", x"72", x"73", x"72", x"6f", x"6f", x"70", x"72", x"73", x"74", 
        x"73", x"71", x"71", x"71", x"71", x"72", x"71", x"70", x"70", x"70", x"71", x"71", x"72", x"74", x"72", 
        x"71", x"72", x"70", x"6f", x"6f", x"71", x"73", x"73", x"72", x"71", x"71", x"71", x"71", x"70", x"6e", 
        x"6c", x"71", x"73", x"73", x"73", x"71", x"71", x"70", x"70", x"70", x"71", x"70", x"6f", x"6e", x"6f", 
        x"70", x"71", x"71", x"71", x"70", x"6f", x"6e", x"6e", x"72", x"71", x"71", x"72", x"73", x"72", x"71", 
        x"70", x"6f", x"6c", x"6d", x"6e", x"6d", x"6c", x"70", x"70", x"70", x"71", x"71", x"6f", x"72", x"70", 
        x"6e", x"70", x"70", x"6d", x"6c", x"6d", x"6f", x"71", x"71", x"6f", x"6c", x"70", x"71", x"6f", x"6a", 
        x"6e", x"71", x"71", x"6f", x"70", x"73", x"71", x"6e", x"6f", x"6e", x"6e", x"70", x"6f", x"6e", x"6e", 
        x"6d", x"6e", x"6f", x"6f", x"6e", x"70", x"70", x"6e", x"6e", x"6e", x"6e", x"6d", x"6f", x"70", x"6e", 
        x"6d", x"6f", x"6f", x"6d", x"6c", x"6f", x"6e", x"6b", x"6f", x"70", x"6d", x"6f", x"6f", x"6d", x"6b", 
        x"6b", x"6d", x"6a", x"6f", x"6c", x"6b", x"6c", x"6c", x"6c", x"6b", x"6a", x"6c", x"6d", x"6d", x"6c", 
        x"6c", x"6b", x"68", x"69", x"6a", x"69", x"6b", x"6d", x"6c", x"69", x"68", x"6a", x"6c", x"69", x"69", 
        x"6c", x"6d", x"6c", x"6c", x"6b", x"6a", x"6b", x"6b", x"6a", x"68", x"69", x"6b", x"6a", x"6a", x"69", 
        x"68", x"6b", x"6f", x"6e", x"6c", x"6c", x"6c", x"6c", x"6b", x"6b", x"6d", x"69", x"69", x"6c", x"69", 
        x"67", x"68", x"66", x"69", x"6d", x"6f", x"6c", x"6a", x"6a", x"69", x"69", x"69", x"6a", x"69", x"69", 
        x"68", x"68", x"6a", x"6a", x"69", x"68", x"69", x"69", x"65", x"68", x"69", x"66", x"66", x"68", x"67", 
        x"66", x"66", x"67", x"67", x"67", x"67", x"69", x"6a", x"6a", x"68", x"68", x"6a", x"69", x"67", x"67", 
        x"67", x"67", x"67", x"67", x"68", x"68", x"68", x"67", x"67", x"67", x"67", x"66", x"67", x"67", x"64", 
        x"66", x"69", x"69", x"67", x"66", x"66", x"66", x"66", x"65", x"65", x"66", x"66", x"64", x"65", x"66", 
        x"67", x"66", x"67", x"68", x"69", x"6c", x"6b", x"6a", x"6a", x"68", x"66", x"65", x"67", x"68", x"68", 
        x"6b", x"6b", x"67", x"67", x"66", x"66", x"68", x"68", x"66", x"64", x"66", x"67", x"67", x"66", x"67", 
        x"67", x"67", x"6a", x"69", x"67", x"68", x"67", x"66", x"67", x"69", x"68", x"69", x"6a", x"67", x"65", 
        x"65", x"66", x"65", x"64", x"67", x"69", x"68", x"66", x"67", x"69", x"69", x"68", x"6a", x"69", x"65", 
        x"65", x"69", x"69", x"67", x"67", x"6a", x"6d", x"66", x"69", x"6e", x"69", x"68", x"69", x"68", x"67", 
        x"64", x"63", x"67", x"6a", x"6b", x"68", x"69", x"68", x"68", x"6a", x"69", x"6c", x"69", x"6a", x"68", 
        x"66", x"6b", x"6b", x"6b", x"68", x"65", x"68", x"6b", x"6c", x"6b", x"6b", x"6b", x"6a", x"6a", x"6c", 
        x"6b", x"6a", x"6a", x"6b", x"6c", x"6b", x"6c", x"6f", x"6e", x"6a", x"6a", x"6c", x"6b", x"6d", x"6d", 
        x"6d", x"6a", x"69", x"6b", x"6e", x"6d", x"6b", x"6b", x"6e", x"6d", x"6d", x"6e", x"6f", x"6d", x"6e", 
        x"6e", x"6f", x"6e", x"6c", x"6b", x"6c", x"6e", x"6e", x"6e", x"70", x"6d", x"6e", x"6c", x"6b", x"6c", 
        x"6c", x"6c", x"69", x"68", x"87", x"bc", x"c9", x"9c", x"a0", x"c2", x"d2", x"cb", x"ca", x"cc", x"cc", 
        x"d0", x"ce", x"cc", x"cc", x"ca", x"ca", x"cd", x"d0", x"cf", x"ce", x"ce", x"cf", x"cf", x"ce", x"cd", 
        x"cd", x"cd", x"ce", x"cf", x"d0", x"cf", x"cd", x"cb", x"cc", x"cc", x"cc", x"cc", x"cc", x"cd", x"cc", 
        x"cb", x"ca", x"cc", x"cc", x"cc", x"cc", x"cc", x"d1", x"cc", x"cf", x"d0", x"d0", x"d1", x"cf", x"b9", 
        x"7a", x"5e", x"5d", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5f", x"5f", x"65", x"a4", x"ed", 
        x"f9", x"f9", x"d9", x"7d", x"5c", x"5b", x"5d", x"5e", x"5d", x"5b", x"5c", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5d", x"5c", x"5e", x"5e", x"5c", x"5c", x"5e", x"5d", x"5d", x"62", x"75", x"a4", x"ca", x"d9", 
        x"e3", x"d0", x"ad", x"86", x"68", x"65", x"6f", x"75", x"76", x"76", x"77", x"77", x"77", x"77", x"75", 
        x"72", x"75", x"75", x"74", x"73", x"74", x"76", x"77", x"77", x"74", x"73", x"75", x"75", x"74", x"74", 
        x"72", x"73", x"74", x"74", x"76", x"75", x"75", x"77", x"75", x"74", x"74", x"75", x"76", x"76", x"73", 
        x"70", x"71", x"72", x"72", x"74", x"76", x"74", x"73", x"75", x"74", x"73", x"72", x"73", x"73", x"74", 
        x"74", x"74", x"73", x"77", x"74", x"73", x"73", x"72", x"71", x"71", x"73", x"74", x"73", x"74", x"74", 
        x"72", x"72", x"73", x"73", x"73", x"73", x"74", x"74", x"73", x"72", x"73", x"71", x"71", x"6e", x"71", 
        x"73", x"72", x"71", x"70", x"71", x"72", x"71", x"72", x"73", x"74", x"72", x"71", x"73", x"73", x"6f", 
        x"70", x"76", x"75", x"71", x"72", x"74", x"73", x"72", x"74", x"73", x"73", x"73", x"73", x"73", x"73", 
        x"73", x"74", x"74", x"73", x"6e", x"70", x"71", x"6f", x"6f", x"71", x"73", x"73", x"71", x"6f", x"6f", 
        x"70", x"70", x"70", x"6f", x"6f", x"70", x"71", x"72", x"71", x"6f", x"72", x"73", x"74", x"75", x"75", 
        x"73", x"72", x"73", x"74", x"73", x"73", x"71", x"70", x"6f", x"6f", x"70", x"70", x"72", x"73", x"70", 
        x"70", x"70", x"70", x"70", x"70", x"70", x"71", x"72", x"72", x"74", x"70", x"6e", x"70", x"73", x"73", 
        x"70", x"6f", x"6f", x"70", x"71", x"70", x"6f", x"6e", x"6f", x"70", x"6f", x"6d", x"6d", x"6c", x"6c", 
        x"6e", x"6f", x"70", x"70", x"6f", x"70", x"70", x"70", x"70", x"6f", x"70", x"72", x"73", x"73", x"71", 
        x"6f", x"6d", x"6d", x"6f", x"6e", x"6e", x"70", x"73", x"71", x"6f", x"71", x"72", x"71", x"70", x"6c", 
        x"6b", x"70", x"71", x"6f", x"6e", x"70", x"70", x"70", x"70", x"70", x"70", x"71", x"6f", x"6a", x"6c", 
        x"72", x"70", x"6f", x"71", x"70", x"70", x"71", x"6f", x"71", x"71", x"71", x"74", x"72", x"71", x"70", 
        x"6f", x"70", x"71", x"71", x"70", x"70", x"6f", x"6f", x"70", x"70", x"6e", x"6c", x"6f", x"71", x"6f", 
        x"6f", x"71", x"6f", x"6c", x"6a", x"6e", x"6e", x"6e", x"71", x"71", x"6d", x"6e", x"6f", x"6e", x"6d", 
        x"6d", x"6f", x"6c", x"70", x"6e", x"6b", x"6b", x"6d", x"6e", x"6d", x"6b", x"6a", x"6d", x"6d", x"6b", 
        x"6b", x"6b", x"69", x"69", x"6a", x"6a", x"68", x"6a", x"6c", x"6a", x"68", x"6a", x"6c", x"69", x"69", 
        x"6c", x"6d", x"6b", x"6a", x"6a", x"6a", x"6c", x"6c", x"6a", x"69", x"6a", x"6d", x"6a", x"6a", x"6a", 
        x"6a", x"6d", x"6a", x"67", x"67", x"68", x"6a", x"6a", x"69", x"6b", x"6c", x"6b", x"69", x"69", x"69", 
        x"69", x"6b", x"69", x"6a", x"6b", x"6b", x"6a", x"69", x"69", x"68", x"6a", x"6c", x"6c", x"6a", x"69", 
        x"69", x"69", x"6b", x"6b", x"68", x"67", x"67", x"66", x"68", x"6a", x"6b", x"6a", x"6b", x"6c", x"6b", 
        x"6a", x"6a", x"6a", x"6a", x"68", x"67", x"68", x"69", x"68", x"68", x"68", x"69", x"68", x"67", x"67", 
        x"66", x"67", x"69", x"6a", x"6a", x"6a", x"69", x"69", x"68", x"68", x"68", x"69", x"68", x"67", x"67", 
        x"6a", x"69", x"66", x"67", x"68", x"67", x"67", x"66", x"66", x"67", x"66", x"65", x"65", x"69", x"69", 
        x"6c", x"6a", x"68", x"68", x"68", x"69", x"68", x"68", x"69", x"69", x"67", x"66", x"66", x"67", x"68", 
        x"69", x"69", x"68", x"67", x"65", x"66", x"68", x"67", x"66", x"64", x"65", x"65", x"67", x"67", x"66", 
        x"67", x"67", x"6a", x"69", x"67", x"6b", x"69", x"67", x"68", x"69", x"68", x"68", x"69", x"69", x"65", 
        x"64", x"66", x"66", x"65", x"66", x"67", x"67", x"66", x"68", x"6a", x"69", x"67", x"68", x"6a", x"68", 
        x"67", x"6a", x"6a", x"67", x"65", x"69", x"6a", x"64", x"66", x"6b", x"69", x"69", x"69", x"68", x"68", 
        x"66", x"65", x"69", x"69", x"6c", x"6a", x"6c", x"6a", x"6b", x"6d", x"6d", x"6d", x"6a", x"6a", x"69", 
        x"69", x"6d", x"6a", x"6b", x"69", x"67", x"69", x"69", x"6c", x"6b", x"69", x"6a", x"6b", x"6b", x"6b", 
        x"6b", x"6c", x"6c", x"6c", x"6d", x"6c", x"6d", x"71", x"71", x"6e", x"6c", x"6e", x"6c", x"6e", x"6e", 
        x"6d", x"69", x"69", x"6d", x"6e", x"6b", x"6a", x"6b", x"69", x"6d", x"71", x"70", x"6e", x"6c", x"6c", 
        x"6f", x"70", x"6f", x"6d", x"6c", x"6e", x"6f", x"6e", x"6f", x"72", x"6f", x"6e", x"6d", x"6c", x"6e", 
        x"6a", x"69", x"6c", x"8f", x"c6", x"bd", x"95", x"9f", x"c6", x"ce", x"cd", x"cc", x"cc", x"ca", x"cc", 
        x"cf", x"cd", x"cb", x"cb", x"cb", x"cb", x"cd", x"cf", x"cf", x"ce", x"ce", x"cf", x"cf", x"ce", x"cd", 
        x"cd", x"ce", x"cf", x"cf", x"cf", x"cf", x"cd", x"ca", x"cc", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", 
        x"ca", x"cb", x"cc", x"cc", x"cc", x"cd", x"cd", x"d1", x"cd", x"d0", x"d0", x"d1", x"d1", x"cf", x"ba", 
        x"7b", x"5f", x"5c", x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5f", x"5f", x"71", x"c8", x"f6", 
        x"f9", x"f7", x"c0", x"6c", x"5b", x"5c", x"5b", x"5f", x"5e", x"5c", x"5f", x"5f", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5c", x"5d", x"5e", x"5c", x"5c", x"5e", x"5e", x"5e", x"5d", x"60", x"90", x"c6", x"c9", 
        x"ce", x"d9", x"e5", x"d3", x"b0", x"89", x"71", x"68", x"6e", x"72", x"75", x"76", x"74", x"75", x"78", 
        x"78", x"78", x"77", x"74", x"73", x"74", x"76", x"77", x"76", x"74", x"75", x"78", x"77", x"74", x"74", 
        x"75", x"77", x"75", x"74", x"77", x"77", x"75", x"75", x"74", x"74", x"74", x"75", x"74", x"75", x"74", 
        x"71", x"71", x"73", x"71", x"73", x"76", x"73", x"73", x"75", x"74", x"72", x"73", x"74", x"72", x"74", 
        x"73", x"72", x"6f", x"75", x"72", x"72", x"72", x"71", x"71", x"72", x"72", x"72", x"71", x"72", x"72", 
        x"72", x"73", x"74", x"74", x"72", x"73", x"77", x"75", x"74", x"73", x"74", x"72", x"71", x"70", x"74", 
        x"76", x"73", x"70", x"70", x"72", x"72", x"71", x"72", x"74", x"72", x"70", x"71", x"71", x"71", x"6e", 
        x"6f", x"74", x"74", x"72", x"73", x"73", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"71", x"71", 
        x"73", x"74", x"73", x"73", x"74", x"71", x"71", x"71", x"70", x"71", x"75", x"76", x"74", x"72", x"71", 
        x"72", x"72", x"72", x"71", x"71", x"72", x"72", x"72", x"71", x"71", x"73", x"75", x"74", x"75", x"76", 
        x"74", x"74", x"74", x"73", x"73", x"73", x"71", x"71", x"6f", x"6e", x"6f", x"6f", x"71", x"73", x"70", 
        x"70", x"70", x"71", x"72", x"72", x"71", x"70", x"71", x"73", x"72", x"6e", x"6c", x"6d", x"71", x"72", 
        x"71", x"6e", x"6e", x"6f", x"6f", x"6e", x"6e", x"6e", x"70", x"71", x"70", x"6e", x"70", x"6f", x"6e", 
        x"6f", x"6f", x"70", x"6f", x"6f", x"71", x"73", x"72", x"72", x"71", x"71", x"72", x"71", x"6f", x"6e", 
        x"6e", x"6c", x"6f", x"70", x"6d", x"6f", x"72", x"72", x"71", x"70", x"6f", x"6f", x"70", x"6f", x"6c", 
        x"6c", x"71", x"72", x"70", x"6f", x"72", x"72", x"70", x"71", x"71", x"72", x"73", x"6f", x"6a", x"6e", 
        x"72", x"70", x"70", x"72", x"71", x"71", x"71", x"6f", x"71", x"71", x"71", x"73", x"71", x"70", x"6f", 
        x"6f", x"70", x"71", x"71", x"70", x"72", x"6f", x"6d", x"6e", x"6f", x"6e", x"6e", x"70", x"71", x"6f", 
        x"70", x"70", x"6f", x"6f", x"6b", x"6c", x"6e", x"70", x"70", x"6f", x"6e", x"6d", x"6f", x"6e", x"6f", 
        x"6d", x"6e", x"6c", x"6d", x"6f", x"6d", x"6d", x"6e", x"6f", x"6d", x"6a", x"6a", x"6c", x"6c", x"6a", 
        x"6b", x"6b", x"6a", x"6a", x"6b", x"6a", x"6a", x"6b", x"6c", x"6b", x"6a", x"6b", x"6a", x"68", x"69", 
        x"6b", x"6b", x"69", x"6a", x"6b", x"6a", x"6c", x"6d", x"6a", x"6a", x"69", x"6b", x"6a", x"6a", x"6c", 
        x"6b", x"6d", x"6b", x"67", x"68", x"67", x"6b", x"6b", x"68", x"6b", x"6a", x"6c", x"6a", x"6b", x"6c", 
        x"6b", x"6c", x"6c", x"6c", x"6a", x"68", x"68", x"69", x"6a", x"6a", x"6b", x"6c", x"6a", x"68", x"67", 
        x"67", x"68", x"6b", x"6b", x"69", x"69", x"69", x"68", x"69", x"68", x"68", x"6a", x"6c", x"6b", x"6a", 
        x"6a", x"6c", x"6c", x"6b", x"6a", x"68", x"68", x"67", x"67", x"68", x"67", x"68", x"68", x"68", x"67", 
        x"66", x"67", x"69", x"69", x"6a", x"6a", x"6b", x"6a", x"68", x"67", x"68", x"69", x"68", x"68", x"6b", 
        x"6b", x"68", x"66", x"67", x"68", x"68", x"69", x"67", x"67", x"69", x"68", x"66", x"68", x"6a", x"69", 
        x"69", x"68", x"67", x"67", x"67", x"67", x"66", x"65", x"67", x"6b", x"69", x"67", x"64", x"64", x"65", 
        x"66", x"6a", x"6a", x"65", x"69", x"68", x"65", x"66", x"66", x"64", x"66", x"65", x"69", x"68", x"67", 
        x"67", x"67", x"6b", x"69", x"66", x"6b", x"69", x"66", x"67", x"69", x"68", x"67", x"69", x"6a", x"65", 
        x"63", x"66", x"67", x"65", x"65", x"68", x"67", x"64", x"65", x"68", x"69", x"69", x"67", x"68", x"6b", 
        x"6b", x"6b", x"6a", x"67", x"65", x"66", x"67", x"68", x"67", x"6b", x"6d", x"67", x"64", x"65", x"6b", 
        x"6b", x"6a", x"6c", x"6b", x"6a", x"68", x"6c", x"69", x"6a", x"6c", x"6d", x"68", x"69", x"6c", x"6a", 
        x"69", x"6a", x"67", x"69", x"6a", x"6b", x"6a", x"67", x"6a", x"6c", x"69", x"69", x"6a", x"6b", x"6a", 
        x"6b", x"6d", x"6e", x"6b", x"6e", x"6d", x"6b", x"6c", x"6f", x"6e", x"6c", x"6f", x"6d", x"70", x"6f", 
        x"6f", x"6b", x"6b", x"70", x"6f", x"6b", x"6c", x"6e", x"6a", x"6e", x"6f", x"6c", x"6b", x"6c", x"6c", 
        x"6a", x"6d", x"6f", x"6d", x"6d", x"70", x"71", x"6e", x"6d", x"6e", x"6b", x"6c", x"6d", x"6c", x"70", 
        x"64", x"6c", x"ab", x"d7", x"a1", x"8c", x"b3", x"ca", x"ce", x"cc", x"c9", x"cb", x"cd", x"cc", x"ca", 
        x"cc", x"cd", x"cc", x"cb", x"cd", x"cf", x"ce", x"ce", x"cf", x"ce", x"ce", x"ce", x"ce", x"cd", x"cc", 
        x"ce", x"d0", x"d0", x"ce", x"cd", x"cd", x"cc", x"c9", x"cc", x"ce", x"cd", x"cd", x"cd", x"cd", x"cd", 
        x"ca", x"cb", x"cd", x"cc", x"cc", x"cd", x"cd", x"d1", x"cd", x"d1", x"d2", x"d2", x"d2", x"cf", x"bb", 
        x"7c", x"5f", x"5c", x"5f", x"60", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"84", x"e5", x"f9", 
        x"fa", x"ed", x"9f", x"60", x"5d", x"5d", x"5e", x"5f", x"5f", x"5f", x"5d", x"5c", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"5f", x"5f", 
        x"5f", x"5f", x"5f", x"5e", x"5e", x"5f", x"5f", x"60", x"5f", x"5e", x"61", x"5e", x"90", x"df", x"ea", 
        x"dd", x"ca", x"c5", x"d2", x"e7", x"e0", x"c6", x"96", x"68", x"5d", x"6d", x"7a", x"76", x"73", x"76", 
        x"7a", x"77", x"77", x"77", x"76", x"76", x"75", x"75", x"76", x"75", x"75", x"76", x"74", x"73", x"76", 
        x"75", x"76", x"78", x"77", x"78", x"75", x"75", x"75", x"73", x"75", x"75", x"74", x"73", x"75", x"75", 
        x"74", x"73", x"74", x"72", x"72", x"74", x"70", x"74", x"75", x"74", x"72", x"74", x"74", x"71", x"78", 
        x"77", x"72", x"6f", x"75", x"74", x"75", x"73", x"72", x"75", x"74", x"71", x"6f", x"70", x"71", x"72", 
        x"74", x"76", x"77", x"77", x"75", x"76", x"77", x"73", x"72", x"72", x"75", x"72", x"72", x"73", x"73", 
        x"73", x"73", x"72", x"72", x"72", x"73", x"72", x"74", x"76", x"74", x"72", x"74", x"70", x"71", x"70", 
        x"70", x"71", x"71", x"73", x"75", x"72", x"71", x"72", x"70", x"70", x"71", x"71", x"74", x"72", x"72", 
        x"75", x"76", x"74", x"72", x"72", x"6f", x"71", x"73", x"71", x"70", x"75", x"76", x"75", x"73", x"72", 
        x"73", x"72", x"72", x"73", x"74", x"74", x"73", x"72", x"72", x"74", x"74", x"71", x"71", x"74", x"74", 
        x"72", x"73", x"74", x"73", x"72", x"72", x"72", x"71", x"70", x"71", x"73", x"72", x"74", x"75", x"6f", 
        x"6f", x"6e", x"72", x"74", x"74", x"71", x"6e", x"70", x"73", x"72", x"71", x"70", x"70", x"6f", x"70", 
        x"72", x"70", x"71", x"71", x"70", x"6f", x"70", x"73", x"71", x"70", x"6f", x"6f", x"73", x"72", x"70", 
        x"72", x"71", x"71", x"6f", x"6d", x"71", x"73", x"72", x"72", x"71", x"72", x"73", x"73", x"72", x"71", 
        x"71", x"6b", x"6f", x"71", x"6e", x"72", x"71", x"6e", x"71", x"73", x"6f", x"6e", x"6f", x"72", x"6f", 
        x"6e", x"70", x"6f", x"6b", x"6a", x"6e", x"70", x"72", x"74", x"72", x"6e", x"70", x"71", x"70", x"70", 
        x"72", x"70", x"72", x"72", x"6f", x"71", x"71", x"6f", x"70", x"70", x"70", x"71", x"6e", x"6e", x"6e", 
        x"6d", x"6e", x"6f", x"6f", x"6f", x"72", x"70", x"6f", x"70", x"70", x"6d", x"6d", x"6e", x"70", x"6e", 
        x"6f", x"6f", x"6f", x"72", x"6f", x"6d", x"6d", x"6f", x"6d", x"6c", x"6f", x"6e", x"6c", x"6c", x"6e", 
        x"6a", x"6b", x"6a", x"67", x"6b", x"6d", x"70", x"70", x"6e", x"6e", x"6f", x"6a", x"6b", x"6b", x"6a", 
        x"6a", x"6c", x"6a", x"6a", x"6a", x"6b", x"6f", x"6f", x"6c", x"69", x"6c", x"6d", x"6a", x"69", x"6a", 
        x"6b", x"68", x"67", x"6d", x"6c", x"68", x"6a", x"6b", x"6a", x"6b", x"65", x"69", x"6a", x"6c", x"6d", 
        x"6a", x"6b", x"6c", x"68", x"69", x"68", x"6c", x"6b", x"68", x"6c", x"67", x"69", x"6a", x"6d", x"70", 
        x"6a", x"68", x"6a", x"6c", x"6a", x"68", x"6b", x"6f", x"6d", x"66", x"68", x"69", x"68", x"68", x"6a", 
        x"6b", x"6b", x"6d", x"6d", x"6a", x"69", x"69", x"68", x"69", x"66", x"66", x"6a", x"6c", x"6b", x"69", 
        x"66", x"67", x"6a", x"6a", x"6a", x"69", x"6a", x"6a", x"6b", x"6b", x"6a", x"69", x"68", x"68", x"69", 
        x"69", x"68", x"68", x"68", x"69", x"6a", x"6b", x"6a", x"69", x"68", x"68", x"69", x"68", x"68", x"6b", 
        x"68", x"67", x"68", x"68", x"68", x"6a", x"6c", x"6a", x"6a", x"6b", x"68", x"67", x"68", x"6b", x"69", 
        x"6a", x"6a", x"6a", x"6b", x"67", x"67", x"67", x"68", x"64", x"66", x"64", x"66", x"69", x"68", x"67", 
        x"67", x"6a", x"69", x"67", x"67", x"67", x"65", x"64", x"66", x"67", x"68", x"68", x"67", x"66", x"64", 
        x"65", x"67", x"68", x"66", x"64", x"68", x"6a", x"66", x"67", x"67", x"67", x"6a", x"68", x"68", x"67", 
        x"67", x"68", x"68", x"67", x"67", x"68", x"67", x"67", x"6a", x"6a", x"69", x"6a", x"68", x"68", x"6c", 
        x"6c", x"69", x"68", x"69", x"6b", x"6b", x"6d", x"6d", x"6a", x"68", x"69", x"6a", x"6a", x"68", x"6b", 
        x"6a", x"69", x"6b", x"69", x"6d", x"68", x"6a", x"69", x"69", x"6a", x"6e", x"6d", x"6b", x"6c", x"6b", 
        x"69", x"6a", x"6d", x"6e", x"6b", x"6a", x"6b", x"69", x"6b", x"6c", x"6a", x"69", x"6c", x"6b", x"69", 
        x"6a", x"6a", x"6c", x"69", x"6b", x"6a", x"6c", x"6c", x"6a", x"6c", x"6d", x"6c", x"6a", x"6c", x"6f", 
        x"6d", x"6f", x"6d", x"6e", x"6e", x"6a", x"6b", x"6e", x"6d", x"6c", x"6c", x"6d", x"6f", x"6e", x"6d", 
        x"6f", x"70", x"6e", x"6c", x"6b", x"6b", x"6c", x"6d", x"6d", x"6f", x"6e", x"6e", x"6f", x"6b", x"63", 
        x"81", x"c0", x"c4", x"98", x"95", x"c5", x"d9", x"d1", x"cc", x"cb", x"c9", x"ca", x"cd", x"cd", x"cc", 
        x"cd", x"ce", x"cd", x"cd", x"cd", x"ce", x"ce", x"cd", x"cd", x"cc", x"cc", x"cc", x"cc", x"cd", x"cd", 
        x"cb", x"cb", x"ce", x"cb", x"cc", x"ce", x"cc", x"cb", x"cb", x"cc", x"cd", x"cd", x"cc", x"cc", x"cd", 
        x"cb", x"ca", x"ca", x"cb", x"cb", x"cb", x"ce", x"d3", x"cd", x"cf", x"d0", x"d2", x"d2", x"cf", x"ba", 
        x"7a", x"5f", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"5e", x"9a", x"f1", x"f9", 
        x"f9", x"e4", x"8e", x"5b", x"5e", x"5f", x"5f", x"5f", x"60", x"5e", x"5b", x"5c", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"5e", x"5e", x"5d", x"5e", x"5e", x"8e", x"df", x"ee", 
        x"ee", x"ea", x"e2", x"d3", x"c6", x"cc", x"de", x"e2", x"cf", x"a9", x"81", x"6b", x"71", x"76", x"77", 
        x"79", x"79", x"70", x"74", x"79", x"77", x"76", x"71", x"75", x"75", x"74", x"76", x"76", x"74", x"76", 
        x"78", x"77", x"77", x"77", x"77", x"77", x"76", x"76", x"75", x"75", x"77", x"77", x"78", x"78", x"77", 
        x"74", x"75", x"76", x"74", x"73", x"74", x"74", x"74", x"74", x"75", x"74", x"74", x"74", x"74", x"74", 
        x"75", x"76", x"78", x"79", x"76", x"72", x"74", x"76", x"75", x"75", x"74", x"74", x"73", x"73", x"73", 
        x"72", x"73", x"76", x"76", x"73", x"73", x"74", x"72", x"73", x"74", x"75", x"72", x"72", x"73", x"73", 
        x"74", x"73", x"73", x"73", x"74", x"74", x"72", x"72", x"76", x"74", x"6d", x"71", x"72", x"72", x"74", 
        x"73", x"72", x"72", x"73", x"73", x"73", x"71", x"71", x"71", x"71", x"71", x"71", x"74", x"75", x"74", 
        x"73", x"74", x"73", x"73", x"75", x"75", x"74", x"71", x"6f", x"71", x"73", x"71", x"72", x"73", x"73", 
        x"72", x"72", x"73", x"74", x"72", x"71", x"72", x"71", x"70", x"73", x"76", x"73", x"73", x"72", x"70", 
        x"72", x"72", x"71", x"73", x"71", x"70", x"72", x"73", x"73", x"74", x"74", x"73", x"72", x"6f", x"70", 
        x"72", x"70", x"74", x"73", x"72", x"71", x"71", x"72", x"72", x"71", x"70", x"70", x"70", x"70", x"70", 
        x"71", x"71", x"70", x"6f", x"70", x"72", x"73", x"72", x"6f", x"6e", x"6e", x"6e", x"6f", x"6f", x"6f", 
        x"70", x"73", x"72", x"6f", x"6e", x"70", x"71", x"6f", x"71", x"72", x"73", x"73", x"72", x"70", x"6f", 
        x"72", x"6e", x"71", x"73", x"70", x"72", x"71", x"70", x"70", x"70", x"70", x"73", x"75", x"70", x"6e", 
        x"6f", x"71", x"70", x"6f", x"70", x"70", x"6e", x"6c", x"70", x"6f", x"70", x"71", x"71", x"6f", x"6f", 
        x"6f", x"6f", x"71", x"72", x"71", x"72", x"6f", x"6f", x"71", x"6e", x"6e", x"71", x"6f", x"6f", x"6d", 
        x"6f", x"72", x"72", x"6f", x"6e", x"70", x"70", x"6c", x"6b", x"6d", x"70", x"6f", x"70", x"71", x"72", 
        x"71", x"71", x"71", x"6f", x"6f", x"6e", x"6c", x"6d", x"6d", x"6c", x"6e", x"70", x"6c", x"6e", x"6e", 
        x"6c", x"6d", x"6f", x"6e", x"70", x"6f", x"6c", x"6e", x"6e", x"69", x"6b", x"6d", x"6c", x"6b", x"6c", 
        x"6c", x"6c", x"6a", x"6a", x"6b", x"6b", x"6c", x"6f", x"6d", x"6b", x"6e", x"6d", x"69", x"6a", x"6c", 
        x"6b", x"69", x"6a", x"6c", x"6c", x"6b", x"6c", x"6d", x"6c", x"6c", x"6c", x"6c", x"6b", x"6b", x"69", 
        x"6a", x"6c", x"6b", x"6b", x"6d", x"6b", x"6b", x"6b", x"6d", x"6c", x"6a", x"6a", x"6c", x"6b", x"6a", 
        x"6c", x"6c", x"6b", x"6b", x"69", x"6a", x"6b", x"6a", x"6c", x"6a", x"68", x"6b", x"6b", x"6b", x"6c", 
        x"6c", x"6c", x"6a", x"69", x"6c", x"6b", x"6b", x"6c", x"6c", x"69", x"68", x"68", x"69", x"6a", x"6b", 
        x"6a", x"68", x"68", x"6a", x"68", x"66", x"69", x"6a", x"6a", x"69", x"68", x"68", x"69", x"6c", x"6a", 
        x"68", x"69", x"68", x"68", x"69", x"6a", x"6c", x"6c", x"69", x"68", x"69", x"6a", x"69", x"69", x"6c", 
        x"6a", x"67", x"6a", x"6b", x"6b", x"69", x"67", x"6b", x"6c", x"69", x"68", x"68", x"69", x"69", x"69", 
        x"6b", x"6b", x"6a", x"6c", x"68", x"67", x"68", x"69", x"64", x"67", x"67", x"69", x"6c", x"6b", x"68", 
        x"66", x"69", x"69", x"69", x"68", x"68", x"66", x"65", x"66", x"68", x"68", x"67", x"66", x"66", x"67", 
        x"67", x"69", x"69", x"67", x"67", x"6a", x"69", x"67", x"67", x"67", x"67", x"6a", x"69", x"68", x"68", 
        x"68", x"68", x"68", x"67", x"67", x"67", x"67", x"67", x"69", x"6a", x"6b", x"6c", x"6b", x"6b", x"6e", 
        x"6e", x"6b", x"6b", x"6d", x"6e", x"6b", x"6d", x"6b", x"69", x"67", x"6a", x"6c", x"68", x"66", x"69", 
        x"6b", x"6c", x"70", x"6e", x"6d", x"6a", x"6d", x"6d", x"6b", x"69", x"6a", x"6e", x"6e", x"6d", x"6d", 
        x"6c", x"6c", x"70", x"6e", x"6d", x"6f", x"6e", x"6b", x"6b", x"6e", x"6c", x"69", x"6c", x"6b", x"6a", 
        x"6c", x"6b", x"6e", x"6b", x"6c", x"6a", x"6b", x"6c", x"6c", x"6e", x"6e", x"6d", x"6c", x"6b", x"6d", 
        x"6b", x"6e", x"6d", x"6e", x"6e", x"6b", x"6a", x"6b", x"6b", x"6d", x"6c", x"6b", x"6d", x"6f", x"6e", 
        x"70", x"6f", x"6d", x"6d", x"6c", x"6c", x"6d", x"6e", x"6e", x"6c", x"6f", x"72", x"6d", x"6a", x"7e", 
        x"bc", x"bb", x"91", x"a2", x"c9", x"d0", x"d3", x"ce", x"ce", x"cd", x"cb", x"cc", x"cd", x"cd", x"cd", 
        x"cd", x"ce", x"cd", x"cd", x"cd", x"cd", x"ce", x"cd", x"cd", x"cc", x"cc", x"cc", x"cc", x"cc", x"cc", 
        x"ca", x"ca", x"cd", x"cb", x"cc", x"ce", x"cb", x"cc", x"cd", x"cc", x"cc", x"cc", x"cc", x"cd", x"cd", 
        x"cc", x"ca", x"ca", x"cc", x"cc", x"cc", x"d0", x"d4", x"ce", x"ce", x"ce", x"d0", x"cf", x"cf", x"ba", 
        x"79", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"60", x"ab", x"f3", x"f8", 
        x"fb", x"d9", x"85", x"5c", x"5c", x"5f", x"5f", x"5b", x"5c", x"5e", x"60", x"5f", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"8d", x"de", x"ec", 
        x"ef", x"ee", x"ed", x"ec", x"e5", x"d5", x"c8", x"ca", x"d9", x"e4", x"d9", x"b0", x"83", x"6c", x"6d", 
        x"6f", x"73", x"76", x"73", x"75", x"78", x"76", x"78", x"77", x"77", x"76", x"73", x"74", x"75", x"76", 
        x"77", x"77", x"76", x"75", x"77", x"78", x"78", x"76", x"75", x"76", x"77", x"78", x"78", x"78", x"77", 
        x"75", x"75", x"74", x"73", x"72", x"74", x"75", x"74", x"74", x"74", x"73", x"72", x"74", x"75", x"75", 
        x"75", x"76", x"77", x"78", x"77", x"74", x"75", x"76", x"76", x"75", x"73", x"73", x"75", x"76", x"74", 
        x"73", x"74", x"75", x"76", x"74", x"74", x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"74", 
        x"74", x"73", x"73", x"73", x"74", x"78", x"73", x"73", x"77", x"75", x"73", x"72", x"73", x"74", x"74", 
        x"73", x"74", x"75", x"76", x"74", x"71", x"70", x"72", x"74", x"75", x"77", x"76", x"75", x"75", x"75", 
        x"74", x"73", x"72", x"72", x"73", x"72", x"70", x"70", x"71", x"73", x"73", x"73", x"75", x"76", x"75", 
        x"74", x"73", x"74", x"76", x"74", x"72", x"73", x"73", x"73", x"75", x"75", x"73", x"73", x"73", x"71", 
        x"74", x"73", x"70", x"73", x"71", x"71", x"72", x"73", x"73", x"74", x"74", x"72", x"72", x"6f", x"71", 
        x"74", x"73", x"73", x"72", x"71", x"71", x"71", x"72", x"72", x"70", x"70", x"70", x"72", x"73", x"74", 
        x"74", x"75", x"73", x"71", x"71", x"71", x"70", x"6d", x"6f", x"71", x"70", x"70", x"71", x"71", x"71", 
        x"71", x"72", x"72", x"70", x"70", x"71", x"70", x"6f", x"72", x"73", x"73", x"73", x"71", x"70", x"6f", 
        x"71", x"70", x"72", x"72", x"71", x"71", x"71", x"73", x"73", x"71", x"6f", x"72", x"73", x"6d", x"6c", 
        x"6b", x"6f", x"6f", x"6e", x"70", x"70", x"70", x"70", x"72", x"72", x"71", x"72", x"70", x"6f", x"72", 
        x"6f", x"6d", x"6e", x"70", x"71", x"72", x"71", x"70", x"72", x"6e", x"6e", x"72", x"72", x"70", x"6e", 
        x"6f", x"72", x"72", x"6f", x"6f", x"70", x"70", x"6d", x"6b", x"6e", x"71", x"71", x"6f", x"6c", x"6e", 
        x"6f", x"71", x"74", x"72", x"72", x"6e", x"6c", x"6c", x"6c", x"6c", x"6e", x"70", x"70", x"6e", x"6e", 
        x"6f", x"6c", x"6b", x"6c", x"71", x"6e", x"6a", x"6c", x"6d", x"69", x"6d", x"6f", x"6d", x"6c", x"6c", 
        x"6c", x"6c", x"6b", x"6b", x"6c", x"6c", x"6c", x"70", x"6f", x"6d", x"6f", x"6d", x"68", x"69", x"6c", 
        x"6d", x"6d", x"6d", x"6d", x"6d", x"6c", x"6b", x"6a", x"69", x"69", x"6f", x"6e", x"6a", x"6b", x"6a", 
        x"6a", x"69", x"6b", x"6d", x"6f", x"6e", x"6b", x"6b", x"6e", x"6e", x"6d", x"6d", x"6c", x"6a", x"6a", 
        x"70", x"6d", x"68", x"6b", x"6c", x"6c", x"6a", x"6a", x"6b", x"69", x"66", x"6a", x"6b", x"6a", x"6b", 
        x"6b", x"6c", x"69", x"68", x"6a", x"6a", x"69", x"6b", x"66", x"66", x"67", x"69", x"6b", x"6a", x"6a", 
        x"6e", x"6a", x"67", x"6b", x"6b", x"68", x"68", x"69", x"69", x"6a", x"6b", x"6b", x"6a", x"69", x"67", 
        x"67", x"69", x"69", x"6a", x"6a", x"6a", x"6a", x"6a", x"69", x"6a", x"6a", x"6a", x"6a", x"69", x"6c", 
        x"6c", x"69", x"6b", x"6a", x"6b", x"69", x"64", x"68", x"6a", x"69", x"68", x"69", x"68", x"68", x"67", 
        x"6c", x"6d", x"6b", x"6c", x"67", x"65", x"66", x"6b", x"68", x"6b", x"6b", x"6a", x"69", x"69", x"6a", 
        x"6a", x"69", x"69", x"69", x"68", x"67", x"66", x"68", x"69", x"69", x"6a", x"6a", x"69", x"69", x"69", 
        x"69", x"6a", x"6a", x"69", x"69", x"6b", x"69", x"69", x"67", x"67", x"68", x"68", x"6a", x"69", x"69", 
        x"68", x"69", x"68", x"67", x"67", x"68", x"69", x"69", x"67", x"67", x"69", x"69", x"69", x"69", x"6a", 
        x"6a", x"69", x"6a", x"6b", x"6c", x"6b", x"6c", x"6c", x"6a", x"67", x"68", x"6a", x"6c", x"6a", x"6b", 
        x"6b", x"6b", x"6d", x"6b", x"6d", x"6c", x"6c", x"6d", x"6a", x"69", x"6a", x"69", x"68", x"68", x"69", 
        x"69", x"69", x"6b", x"6b", x"6b", x"69", x"68", x"6a", x"6a", x"69", x"6b", x"6b", x"6d", x"6c", x"6b", 
        x"6d", x"6b", x"6c", x"6b", x"6b", x"69", x"6a", x"6b", x"6a", x"6c", x"6a", x"6b", x"6e", x"6b", x"6c", 
        x"6e", x"6f", x"6b", x"6c", x"6c", x"6b", x"6d", x"6d", x"6b", x"6d", x"6d", x"6b", x"6d", x"6e", x"6f", 
        x"6f", x"6e", x"6e", x"6e", x"6e", x"6e", x"6f", x"6f", x"6f", x"6e", x"6f", x"6f", x"6c", x"6b", x"76", 
        x"9c", x"8c", x"b2", x"cf", x"cc", x"cf", x"d6", x"cc", x"ce", x"ce", x"cc", x"cd", x"ce", x"ce", x"cd", 
        x"cd", x"ce", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"ce", x"cd", x"cc", x"cb", x"cb", x"cb", x"cc", 
        x"cb", x"cb", x"cd", x"cb", x"cc", x"cd", x"cc", x"cd", x"ce", x"cd", x"cb", x"cb", x"cc", x"ce", x"ce", 
        x"cc", x"cb", x"cc", x"cd", x"ce", x"cd", x"cc", x"d1", x"cc", x"ce", x"d0", x"d2", x"d3", x"d0", x"bb", 
        x"78", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"60", x"af", x"f5", x"f7", 
        x"fc", x"d7", x"82", x"5e", x"5d", x"5e", x"61", x"5f", x"5d", x"5e", x"60", x"5f", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"8b", x"de", x"ed", 
        x"ee", x"ed", x"ed", x"ec", x"e9", x"e9", x"e7", x"d8", x"c6", x"ca", x"d7", x"e2", x"d4", x"b6", x"8c", 
        x"6f", x"6e", x"73", x"73", x"74", x"77", x"7b", x"7a", x"76", x"78", x"78", x"74", x"73", x"76", x"78", 
        x"79", x"7a", x"79", x"77", x"75", x"75", x"76", x"75", x"75", x"76", x"77", x"78", x"78", x"78", x"77", 
        x"76", x"76", x"74", x"73", x"72", x"74", x"75", x"75", x"75", x"74", x"72", x"72", x"73", x"76", x"76", 
        x"74", x"74", x"76", x"77", x"77", x"76", x"76", x"76", x"77", x"75", x"74", x"73", x"75", x"76", x"76", 
        x"75", x"75", x"75", x"77", x"76", x"75", x"75", x"75", x"74", x"73", x"73", x"74", x"74", x"73", x"73", 
        x"73", x"73", x"73", x"73", x"74", x"77", x"71", x"73", x"74", x"73", x"74", x"71", x"72", x"74", x"74", 
        x"75", x"75", x"75", x"73", x"72", x"73", x"72", x"73", x"73", x"73", x"76", x"76", x"76", x"75", x"75", 
        x"75", x"73", x"73", x"73", x"72", x"71", x"71", x"71", x"72", x"73", x"74", x"72", x"74", x"75", x"75", 
        x"74", x"73", x"72", x"75", x"73", x"71", x"72", x"72", x"72", x"73", x"74", x"72", x"73", x"73", x"72", 
        x"75", x"74", x"72", x"73", x"73", x"73", x"72", x"72", x"73", x"73", x"73", x"71", x"71", x"6f", x"6f", 
        x"71", x"71", x"72", x"72", x"72", x"71", x"71", x"72", x"73", x"71", x"70", x"71", x"72", x"72", x"72", 
        x"72", x"72", x"72", x"72", x"72", x"72", x"71", x"70", x"72", x"72", x"71", x"71", x"72", x"72", x"72", 
        x"71", x"72", x"73", x"72", x"71", x"72", x"70", x"6e", x"70", x"70", x"70", x"70", x"70", x"6f", x"6f", 
        x"70", x"72", x"71", x"71", x"72", x"71", x"71", x"73", x"73", x"70", x"6f", x"71", x"73", x"71", x"6f", 
        x"6d", x"70", x"6f", x"6e", x"6e", x"6e", x"6e", x"6f", x"70", x"70", x"70", x"70", x"70", x"6f", x"70", 
        x"6f", x"6f", x"70", x"72", x"71", x"70", x"6f", x"6e", x"71", x"70", x"71", x"73", x"74", x"71", x"71", 
        x"70", x"70", x"71", x"72", x"70", x"71", x"73", x"72", x"6f", x"6f", x"71", x"70", x"71", x"71", x"70", 
        x"6e", x"6e", x"6f", x"6d", x"6f", x"6f", x"6e", x"6c", x"6c", x"6d", x"6e", x"6e", x"6f", x"6c", x"6d", 
        x"6f", x"6e", x"6c", x"6b", x"6f", x"6d", x"6a", x"6c", x"6d", x"6c", x"70", x"70", x"6e", x"6d", x"6c", 
        x"6c", x"6d", x"6c", x"6b", x"6d", x"6e", x"6e", x"71", x"70", x"6f", x"6f", x"6a", x"69", x"6c", x"6f", 
        x"6e", x"6b", x"6a", x"6c", x"6b", x"6b", x"6b", x"6a", x"6a", x"6c", x"6d", x"6b", x"68", x"6c", x"6e", 
        x"6e", x"6b", x"6a", x"6c", x"6e", x"6e", x"6d", x"6d", x"70", x"6f", x"6e", x"6e", x"6e", x"6b", x"6b", 
        x"6e", x"6d", x"6b", x"6f", x"6e", x"6c", x"69", x"69", x"6c", x"6c", x"69", x"6b", x"6a", x"69", x"6a", 
        x"68", x"69", x"68", x"67", x"68", x"68", x"69", x"6c", x"6a", x"69", x"68", x"6a", x"6b", x"6b", x"6a", 
        x"6b", x"69", x"69", x"6c", x"6c", x"6a", x"6d", x"6e", x"6a", x"69", x"6a", x"6b", x"6b", x"69", x"68", 
        x"6a", x"6b", x"6b", x"6a", x"69", x"66", x"64", x"68", x"69", x"6b", x"6b", x"6b", x"6a", x"6a", x"6c", 
        x"6c", x"6a", x"6a", x"69", x"6a", x"6a", x"66", x"67", x"68", x"67", x"68", x"6a", x"6a", x"6a", x"69", 
        x"6b", x"6c", x"6b", x"6c", x"67", x"66", x"67", x"6b", x"67", x"69", x"6c", x"69", x"68", x"6b", x"6b", 
        x"69", x"67", x"67", x"69", x"6a", x"69", x"68", x"66", x"68", x"69", x"6a", x"69", x"6a", x"69", x"68", 
        x"67", x"69", x"6a", x"68", x"68", x"69", x"6a", x"6c", x"68", x"68", x"68", x"67", x"6b", x"6a", x"6a", 
        x"6b", x"6a", x"69", x"67", x"66", x"67", x"6a", x"6b", x"69", x"68", x"68", x"66", x"68", x"6b", x"6a", 
        x"6b", x"6c", x"6c", x"6b", x"6a", x"69", x"6c", x"6e", x"6d", x"6a", x"67", x"67", x"6c", x"6c", x"6c", 
        x"6b", x"6b", x"6a", x"69", x"6b", x"6c", x"69", x"6c", x"6a", x"6c", x"6d", x"6b", x"6a", x"6a", x"6c", 
        x"6c", x"6c", x"6d", x"6e", x"6f", x"6c", x"6b", x"6f", x"6e", x"6c", x"6d", x"6c", x"6d", x"6d", x"6c", 
        x"6e", x"6b", x"6b", x"6c", x"6d", x"6c", x"6e", x"6d", x"6a", x"6c", x"6d", x"6b", x"6f", x"6b", x"6c", 
        x"6f", x"6b", x"6c", x"6e", x"6d", x"6c", x"6d", x"6d", x"69", x"6a", x"6c", x"6f", x"70", x"6e", x"6d", 
        x"6d", x"6e", x"6f", x"6f", x"6f", x"6f", x"6f", x"6e", x"6d", x"6f", x"6e", x"6c", x"6f", x"71", x"66", 
        x"89", x"cf", x"d4", x"d2", x"cf", x"d5", x"d8", x"ce", x"cc", x"cb", x"cb", x"cc", x"ce", x"cf", x"cf", 
        x"ce", x"ce", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"ce", x"cd", x"cc", x"cb", x"cb", x"cb", x"cb", 
        x"cc", x"cc", x"cc", x"cc", x"cc", x"cc", x"cc", x"cd", x"ce", x"cd", x"cb", x"ca", x"cc", x"cf", x"ce", 
        x"cd", x"cb", x"cb", x"cc", x"cd", x"cd", x"ce", x"d4", x"cf", x"cf", x"ce", x"cf", x"d0", x"d0", x"bb", 
        x"78", x"5f", x"5f", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"60", x"ab", x"f3", x"f8", 
        x"fa", x"e6", x"99", x"5d", x"5e", x"5d", x"5c", x"5e", x"5d", x"5d", x"5f", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"60", x"87", x"dd", x"ee", 
        x"ee", x"ed", x"ec", x"ec", x"ed", x"ef", x"f0", x"ef", x"ee", x"e4", x"ce", x"c6", x"d7", x"e6", x"e2", 
        x"cd", x"9e", x"79", x"67", x"6f", x"77", x"74", x"71", x"74", x"77", x"79", x"78", x"75", x"72", x"75", 
        x"78", x"78", x"79", x"78", x"76", x"76", x"77", x"76", x"76", x"76", x"77", x"78", x"78", x"77", x"78", 
        x"78", x"78", x"77", x"77", x"76", x"76", x"76", x"76", x"76", x"75", x"74", x"73", x"74", x"76", x"75", 
        x"75", x"76", x"77", x"78", x"77", x"74", x"75", x"76", x"75", x"76", x"78", x"76", x"73", x"74", x"76", 
        x"76", x"74", x"74", x"76", x"76", x"76", x"73", x"76", x"75", x"73", x"74", x"76", x"75", x"73", x"73", 
        x"73", x"73", x"73", x"73", x"73", x"76", x"75", x"76", x"76", x"73", x"73", x"75", x"75", x"74", x"72", 
        x"72", x"73", x"72", x"70", x"72", x"75", x"74", x"73", x"71", x"6f", x"72", x"73", x"75", x"74", x"76", 
        x"76", x"75", x"74", x"76", x"75", x"77", x"77", x"74", x"71", x"72", x"75", x"71", x"72", x"74", x"75", 
        x"75", x"75", x"74", x"77", x"76", x"75", x"75", x"75", x"75", x"76", x"76", x"75", x"73", x"71", x"72", 
        x"75", x"76", x"74", x"74", x"75", x"75", x"73", x"72", x"73", x"74", x"75", x"73", x"74", x"73", x"72", 
        x"72", x"74", x"71", x"72", x"73", x"72", x"72", x"73", x"74", x"74", x"73", x"73", x"74", x"73", x"73", 
        x"73", x"72", x"73", x"74", x"73", x"72", x"71", x"71", x"72", x"70", x"6f", x"6f", x"71", x"71", x"70", 
        x"71", x"73", x"72", x"72", x"72", x"72", x"71", x"70", x"72", x"72", x"72", x"72", x"73", x"73", x"74", 
        x"71", x"74", x"71", x"70", x"72", x"71", x"71", x"74", x"74", x"72", x"70", x"6f", x"70", x"70", x"6f", 
        x"6d", x"71", x"71", x"71", x"73", x"73", x"73", x"71", x"71", x"71", x"70", x"6f", x"6e", x"6d", x"6d", 
        x"6e", x"6f", x"72", x"73", x"73", x"72", x"70", x"6f", x"73", x"72", x"70", x"6c", x"6f", x"71", x"73", 
        x"70", x"6e", x"70", x"74", x"71", x"70", x"72", x"73", x"71", x"70", x"71", x"6f", x"71", x"71", x"70", 
        x"6e", x"6e", x"6e", x"6b", x"6d", x"6e", x"6f", x"6d", x"6d", x"6f", x"70", x"6f", x"6f", x"71", x"6f", 
        x"6e", x"6e", x"6d", x"69", x"6d", x"6c", x"6d", x"6d", x"6d", x"6c", x"6f", x"70", x"6e", x"6d", x"6c", 
        x"6c", x"6d", x"6f", x"6c", x"6e", x"70", x"6f", x"70", x"6e", x"6e", x"6f", x"6b", x"6b", x"6c", x"6d", 
        x"6c", x"69", x"6a", x"6f", x"6e", x"6d", x"6d", x"6c", x"6b", x"6d", x"6d", x"6c", x"6a", x"6d", x"6d", 
        x"6c", x"6a", x"6a", x"6c", x"6d", x"6c", x"6b", x"6b", x"6c", x"6c", x"6c", x"6d", x"6f", x"6e", x"6b", 
        x"68", x"69", x"6c", x"6c", x"6b", x"6c", x"6b", x"6d", x"6e", x"6b", x"6a", x"6d", x"6d", x"6d", x"6e", 
        x"6b", x"69", x"69", x"6a", x"69", x"68", x"6a", x"6c", x"69", x"69", x"6b", x"6e", x"6e", x"6c", x"68", 
        x"69", x"69", x"6b", x"6d", x"6c", x"6b", x"6f", x"6f", x"6c", x"69", x"69", x"6b", x"6c", x"6a", x"69", 
        x"68", x"69", x"6c", x"6c", x"6b", x"69", x"65", x"69", x"6a", x"6b", x"6b", x"6b", x"6b", x"6c", x"6d", 
        x"6b", x"68", x"69", x"6a", x"6b", x"6a", x"6c", x"6a", x"68", x"68", x"6a", x"6b", x"6c", x"6c", x"6a", 
        x"68", x"69", x"69", x"6c", x"69", x"69", x"6b", x"6c", x"69", x"68", x"6b", x"67", x"66", x"6a", x"69", 
        x"69", x"69", x"6a", x"6a", x"69", x"67", x"67", x"6a", x"6a", x"6b", x"6b", x"6a", x"69", x"68", x"67", 
        x"67", x"69", x"6b", x"6a", x"68", x"69", x"6c", x"6d", x"6a", x"69", x"6a", x"68", x"6a", x"69", x"6a", 
        x"6c", x"6c", x"6a", x"69", x"66", x"67", x"69", x"6a", x"69", x"68", x"69", x"69", x"6b", x"6c", x"6b", 
        x"6c", x"6e", x"6e", x"6b", x"69", x"69", x"6a", x"6c", x"6c", x"6b", x"6a", x"69", x"6c", x"6c", x"6b", 
        x"6b", x"6a", x"69", x"6a", x"6a", x"6d", x"6b", x"6d", x"6b", x"6b", x"6b", x"6d", x"6c", x"6c", x"6d", 
        x"6d", x"6d", x"6e", x"6a", x"6c", x"6c", x"6a", x"6a", x"68", x"6a", x"6d", x"6b", x"6d", x"6d", x"6d", 
        x"6f", x"6c", x"6c", x"6c", x"6d", x"6c", x"6d", x"6d", x"6b", x"6d", x"6e", x"6a", x"6c", x"6b", x"70", 
        x"71", x"6c", x"6d", x"6f", x"6e", x"6d", x"6e", x"6f", x"6d", x"6c", x"6d", x"6f", x"6f", x"6e", x"6e", 
        x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6d", x"6c", x"6e", x"6d", x"6c", x"6e", x"6d", 
        x"9d", x"db", x"cf", x"d0", x"ce", x"d1", x"da", x"cc", x"cc", x"cb", x"ca", x"cb", x"cd", x"cd", x"cd", 
        x"cd", x"ce", x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"cd", x"cc", x"cb", x"cb", x"cb", x"cb", x"cb", 
        x"cc", x"cc", x"cb", x"cc", x"cc", x"cb", x"cc", x"cd", x"ce", x"cd", x"cb", x"ca", x"cd", x"cf", x"ce", 
        x"cd", x"cc", x"cb", x"ca", x"ca", x"cb", x"cc", x"d3", x"cf", x"cf", x"cf", x"d1", x"d2", x"d0", x"bb", 
        x"78", x"5f", x"5f", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"60", x"a8", x"f2", x"f9", 
        x"fb", x"f5", x"c9", x"78", x"60", x"5d", x"5e", x"5f", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"82", x"da", x"ed", 
        x"ee", x"ee", x"ed", x"ec", x"ee", x"ef", x"ec", x"ed", x"ef", x"ef", x"ee", x"e4", x"d5", x"cf", x"d5", 
        x"da", x"e1", x"d1", x"a8", x"88", x"76", x"69", x"6d", x"7b", x"7a", x"78", x"78", x"78", x"76", x"75", 
        x"76", x"78", x"79", x"79", x"77", x"76", x"74", x"75", x"76", x"77", x"77", x"78", x"77", x"77", x"77", 
        x"76", x"77", x"77", x"78", x"78", x"76", x"75", x"76", x"77", x"77", x"77", x"76", x"76", x"77", x"77", 
        x"76", x"76", x"76", x"76", x"76", x"74", x"74", x"75", x"77", x"79", x"79", x"76", x"73", x"73", x"75", 
        x"74", x"74", x"74", x"75", x"75", x"74", x"72", x"76", x"76", x"75", x"77", x"77", x"75", x"74", x"73", 
        x"73", x"73", x"74", x"74", x"73", x"75", x"74", x"71", x"73", x"74", x"70", x"74", x"76", x"74", x"71", 
        x"70", x"71", x"74", x"76", x"75", x"75", x"74", x"74", x"73", x"71", x"74", x"74", x"74", x"74", x"76", 
        x"76", x"76", x"76", x"77", x"76", x"77", x"76", x"74", x"73", x"73", x"74", x"75", x"75", x"76", x"77", 
        x"78", x"77", x"76", x"76", x"76", x"74", x"73", x"73", x"75", x"75", x"75", x"75", x"74", x"71", x"73", 
        x"75", x"75", x"73", x"74", x"75", x"75", x"73", x"72", x"73", x"74", x"76", x"75", x"74", x"74", x"72", 
        x"71", x"73", x"71", x"72", x"73", x"72", x"72", x"72", x"73", x"72", x"72", x"72", x"72", x"72", x"73", 
        x"73", x"72", x"73", x"74", x"74", x"73", x"72", x"73", x"73", x"71", x"70", x"70", x"71", x"71", x"70", 
        x"72", x"73", x"71", x"71", x"72", x"72", x"72", x"71", x"70", x"70", x"70", x"71", x"71", x"72", x"72", 
        x"70", x"73", x"71", x"70", x"72", x"71", x"71", x"71", x"71", x"71", x"72", x"71", x"72", x"72", x"72", 
        x"70", x"72", x"71", x"70", x"71", x"71", x"72", x"71", x"71", x"72", x"73", x"73", x"73", x"73", x"70", 
        x"6f", x"6f", x"70", x"72", x"73", x"72", x"6f", x"6f", x"71", x"71", x"71", x"6e", x"72", x"72", x"72", 
        x"70", x"6f", x"70", x"73", x"71", x"6d", x"6e", x"71", x"70", x"71", x"73", x"71", x"70", x"6e", x"6f", 
        x"6f", x"70", x"70", x"6c", x"6d", x"6f", x"70", x"6f", x"6f", x"71", x"71", x"6f", x"6e", x"70", x"71", 
        x"70", x"6e", x"6f", x"6f", x"6f", x"6d", x"6e", x"6f", x"6d", x"6d", x"6d", x"6e", x"6e", x"6e", x"6d", 
        x"6c", x"6e", x"70", x"6d", x"6e", x"70", x"6e", x"6e", x"6b", x"6c", x"6e", x"6d", x"6c", x"6a", x"6a", 
        x"6c", x"6d", x"6c", x"6c", x"6a", x"6b", x"6d", x"6c", x"6d", x"6f", x"6b", x"6d", x"6c", x"6e", x"6c", 
        x"6c", x"6c", x"6b", x"6c", x"6c", x"6b", x"6a", x"6a", x"6a", x"6b", x"6b", x"6b", x"6d", x"6f", x"6f", 
        x"6b", x"6b", x"6e", x"6a", x"69", x"6d", x"6d", x"6b", x"6b", x"6b", x"6a", x"6d", x"6c", x"6d", x"6d", 
        x"6a", x"6c", x"6d", x"6c", x"6a", x"69", x"6a", x"6a", x"68", x"68", x"68", x"69", x"6b", x"6c", x"6c", 
        x"6e", x"6b", x"69", x"6a", x"6d", x"6c", x"6b", x"6d", x"6d", x"6b", x"6b", x"6c", x"6b", x"68", x"68", 
        x"69", x"69", x"6d", x"6b", x"6b", x"6b", x"67", x"6a", x"6b", x"6a", x"6a", x"6a", x"6c", x"6d", x"6d", 
        x"6a", x"68", x"69", x"6d", x"6b", x"69", x"6c", x"6b", x"69", x"6a", x"6b", x"69", x"68", x"69", x"68", 
        x"6a", x"6b", x"6b", x"6d", x"69", x"69", x"6b", x"6b", x"69", x"67", x"6a", x"67", x"67", x"68", x"66", 
        x"68", x"6a", x"6b", x"6b", x"68", x"66", x"67", x"6a", x"6c", x"6c", x"6b", x"6a", x"69", x"68", x"68", 
        x"67", x"69", x"6c", x"6b", x"6b", x"6b", x"6b", x"6b", x"6a", x"6a", x"6a", x"69", x"69", x"6b", x"6b", 
        x"6d", x"6d", x"6c", x"6a", x"69", x"6a", x"6b", x"69", x"68", x"67", x"68", x"69", x"6c", x"6c", x"6a", 
        x"6a", x"6b", x"6c", x"6a", x"6a", x"6c", x"6b", x"6b", x"6b", x"6b", x"6b", x"6a", x"6b", x"6d", x"6b", 
        x"6b", x"6b", x"69", x"6c", x"6d", x"6e", x"6c", x"6a", x"6a", x"6b", x"6a", x"6f", x"6d", x"6c", x"6d", 
        x"6d", x"6d", x"6d", x"6d", x"6c", x"6b", x"6a", x"6c", x"6c", x"6c", x"6c", x"6c", x"6f", x"6e", x"6c", 
        x"6d", x"6a", x"6c", x"6d", x"6e", x"6b", x"6c", x"6d", x"6d", x"6f", x"6f", x"6c", x"6d", x"6c", x"71", 
        x"70", x"6f", x"6c", x"6e", x"6e", x"6d", x"6f", x"70", x"6e", x"6e", x"6f", x"6e", x"6c", x"6d", x"70", 
        x"71", x"6f", x"6e", x"6e", x"6e", x"6e", x"70", x"71", x"6f", x"6c", x"71", x"71", x"6f", x"6f", x"6c", 
        x"9c", x"d9", x"d3", x"ce", x"cd", x"d4", x"d8", x"cd", x"cd", x"cc", x"cb", x"cb", x"cc", x"cc", x"cc", 
        x"cd", x"ce", x"cd", x"cd", x"cd", x"cd", x"ce", x"cd", x"cc", x"cc", x"cb", x"cb", x"cb", x"cb", x"ca", 
        x"cc", x"cc", x"cb", x"cd", x"cd", x"cc", x"cd", x"cd", x"ce", x"cd", x"cc", x"cc", x"cd", x"ce", x"ce", 
        x"ce", x"cd", x"cb", x"ca", x"ca", x"cc", x"cb", x"d3", x"d1", x"d1", x"d0", x"d1", x"d2", x"d0", x"bb", 
        x"79", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"5e", x"98", x"ed", x"fa", 
        x"fa", x"f9", x"ee", x"b7", x"74", x"5d", x"5f", x"63", x"5e", x"5d", x"5e", x"5d", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"60", x"7c", x"d7", x"ed", 
        x"ee", x"ed", x"eb", x"ec", x"ed", x"ee", x"ee", x"ed", x"eb", x"ea", x"ed", x"f0", x"ee", x"e8", x"dc", 
        x"cf", x"d2", x"d9", x"e1", x"d6", x"b2", x"8a", x"75", x"6f", x"71", x"75", x"79", x"79", x"77", x"77", 
        x"77", x"78", x"79", x"79", x"79", x"77", x"75", x"75", x"76", x"77", x"78", x"78", x"77", x"77", x"76", 
        x"75", x"75", x"76", x"78", x"78", x"77", x"75", x"76", x"77", x"78", x"77", x"76", x"76", x"77", x"79", 
        x"77", x"75", x"74", x"75", x"75", x"75", x"75", x"76", x"79", x"7a", x"78", x"75", x"74", x"75", x"75", 
        x"74", x"74", x"75", x"75", x"75", x"73", x"73", x"76", x"75", x"74", x"77", x"77", x"75", x"75", x"73", 
        x"73", x"74", x"75", x"74", x"74", x"75", x"74", x"6f", x"72", x"75", x"72", x"73", x"74", x"73", x"73", 
        x"74", x"75", x"76", x"77", x"77", x"77", x"75", x"75", x"75", x"75", x"77", x"76", x"74", x"74", x"75", 
        x"75", x"75", x"76", x"76", x"74", x"75", x"73", x"72", x"74", x"75", x"72", x"76", x"76", x"75", x"75", 
        x"76", x"75", x"75", x"75", x"76", x"74", x"72", x"73", x"75", x"74", x"73", x"75", x"74", x"72", x"75", 
        x"76", x"73", x"72", x"73", x"73", x"74", x"74", x"73", x"72", x"74", x"78", x"79", x"74", x"73", x"70", 
        x"6e", x"6f", x"71", x"72", x"73", x"73", x"73", x"72", x"72", x"73", x"73", x"73", x"72", x"72", x"71", 
        x"71", x"72", x"73", x"74", x"74", x"73", x"72", x"73", x"73", x"72", x"72", x"72", x"71", x"71", x"72", 
        x"73", x"73", x"6f", x"70", x"73", x"72", x"72", x"73", x"71", x"72", x"73", x"73", x"73", x"73", x"72", 
        x"70", x"71", x"72", x"72", x"72", x"71", x"71", x"72", x"71", x"71", x"72", x"73", x"72", x"73", x"71", 
        x"6d", x"70", x"6f", x"6f", x"71", x"71", x"72", x"6f", x"6f", x"71", x"72", x"72", x"73", x"74", x"70", 
        x"70", x"71", x"73", x"72", x"71", x"6f", x"70", x"71", x"71", x"70", x"72", x"72", x"76", x"74", x"71", 
        x"70", x"70", x"71", x"72", x"71", x"6f", x"70", x"71", x"70", x"71", x"72", x"6f", x"6f", x"6f", x"70", 
        x"70", x"70", x"71", x"6e", x"70", x"71", x"71", x"70", x"70", x"6f", x"6e", x"6e", x"6e", x"6e", x"70", 
        x"71", x"6d", x"6e", x"71", x"70", x"6d", x"6f", x"6f", x"6e", x"6f", x"6c", x"6d", x"6e", x"6e", x"6e", 
        x"6d", x"6e", x"70", x"6d", x"6e", x"70", x"6e", x"6d", x"6b", x"6b", x"6c", x"6b", x"6d", x"6d", x"6d", 
        x"6e", x"6e", x"6c", x"6a", x"68", x"6a", x"6e", x"6c", x"6c", x"6e", x"6c", x"6e", x"6d", x"6e", x"6c", 
        x"6c", x"6b", x"6a", x"6a", x"6b", x"6c", x"6d", x"6e", x"6e", x"6c", x"6b", x"6b", x"6a", x"6c", x"6f", 
        x"6f", x"6d", x"6d", x"6a", x"69", x"6d", x"6d", x"6a", x"68", x"67", x"68", x"6b", x"6b", x"6e", x"6f", 
        x"6a", x"6b", x"6d", x"6d", x"6c", x"6c", x"6b", x"6a", x"6d", x"6d", x"6c", x"6b", x"6a", x"6b", x"6d", 
        x"6b", x"6b", x"6c", x"6b", x"6b", x"6c", x"6e", x"6f", x"6d", x"6a", x"69", x"6a", x"6b", x"6b", x"6c", 
        x"6a", x"6a", x"6e", x"6a", x"6b", x"6e", x"6a", x"6b", x"6b", x"6a", x"6a", x"6b", x"6c", x"6c", x"6c", 
        x"69", x"6a", x"6b", x"6d", x"6a", x"69", x"6b", x"6a", x"6a", x"6b", x"6c", x"69", x"67", x"69", x"68", 
        x"6c", x"6d", x"6c", x"6e", x"6a", x"69", x"6a", x"69", x"69", x"67", x"6c", x"6a", x"6b", x"69", x"66", 
        x"68", x"68", x"68", x"67", x"67", x"68", x"67", x"65", x"68", x"6b", x"6c", x"6b", x"6a", x"6a", x"69", 
        x"66", x"66", x"69", x"6b", x"6c", x"6d", x"68", x"66", x"69", x"6a", x"6a", x"6b", x"69", x"6c", x"6c", 
        x"6c", x"6c", x"6c", x"6c", x"6d", x"6b", x"69", x"69", x"6a", x"69", x"68", x"69", x"6e", x"6f", x"6b", 
        x"68", x"6a", x"6c", x"6d", x"6d", x"6c", x"6b", x"6b", x"6c", x"6c", x"6c", x"6b", x"6a", x"6d", x"6c", 
        x"6d", x"6d", x"6c", x"6e", x"6b", x"6c", x"6d", x"6a", x"6c", x"6c", x"69", x"70", x"6e", x"6a", x"6a", 
        x"6b", x"6a", x"6b", x"6c", x"6a", x"6a", x"6b", x"69", x"6b", x"6c", x"6a", x"6b", x"6f", x"6f", x"6c", 
        x"6b", x"68", x"6b", x"6c", x"6e", x"6c", x"6f", x"70", x"6e", x"70", x"6f", x"70", x"70", x"6e", x"6f", 
        x"6c", x"73", x"6a", x"6c", x"6f", x"6e", x"6f", x"6f", x"6d", x"6b", x"6f", x"72", x"6f", x"6c", x"6f", 
        x"73", x"73", x"71", x"70", x"6f", x"6f", x"70", x"71", x"70", x"6f", x"71", x"72", x"73", x"71", x"6a", 
        x"9a", x"d8", x"cf", x"d0", x"cf", x"d0", x"d6", x"cd", x"cd", x"cc", x"cb", x"cc", x"cd", x"ce", x"ce", 
        x"cd", x"ce", x"cd", x"cd", x"cd", x"cd", x"ce", x"cd", x"cb", x"cb", x"cb", x"cb", x"cb", x"cc", x"cb", 
        x"cb", x"cb", x"c9", x"cd", x"cd", x"cc", x"ce", x"cd", x"ce", x"ce", x"ce", x"cd", x"ce", x"cd", x"cd", 
        x"ce", x"cd", x"cc", x"cb", x"cd", x"ce", x"cd", x"d5", x"d3", x"d2", x"d0", x"d1", x"d2", x"cf", x"ba", 
        x"79", x"60", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"5b", x"7e", x"e3", x"f9", 
        x"f9", x"fa", x"f8", x"ed", x"ba", x"80", x"5d", x"5d", x"5d", x"5c", x"5f", x"5f", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"60", x"5f", x"78", x"d3", x"ec", 
        x"ee", x"ef", x"ed", x"eb", x"ed", x"ee", x"ec", x"ed", x"ef", x"ec", x"ed", x"ee", x"ec", x"ec", x"ef", 
        x"eb", x"df", x"d3", x"cd", x"d4", x"e3", x"e3", x"c7", x"9e", x"7a", x"66", x"6c", x"7a", x"7c", x"78", 
        x"77", x"77", x"77", x"78", x"79", x"7a", x"78", x"77", x"77", x"77", x"78", x"78", x"77", x"77", x"76", 
        x"76", x"75", x"76", x"78", x"7a", x"79", x"78", x"77", x"76", x"76", x"75", x"75", x"76", x"78", x"78", 
        x"76", x"74", x"73", x"75", x"76", x"77", x"77", x"77", x"77", x"77", x"77", x"76", x"75", x"76", x"76", 
        x"75", x"76", x"78", x"78", x"76", x"74", x"77", x"78", x"74", x"72", x"76", x"76", x"73", x"76", x"74", 
        x"73", x"74", x"76", x"75", x"75", x"77", x"76", x"75", x"74", x"74", x"77", x"76", x"73", x"73", x"75", 
        x"75", x"74", x"72", x"72", x"73", x"75", x"72", x"73", x"75", x"76", x"77", x"76", x"76", x"77", x"75", 
        x"74", x"74", x"74", x"72", x"74", x"7a", x"76", x"72", x"75", x"77", x"74", x"77", x"76", x"74", x"75", 
        x"76", x"78", x"77", x"75", x"76", x"74", x"72", x"72", x"75", x"74", x"72", x"75", x"73", x"70", x"75", 
        x"76", x"74", x"73", x"71", x"71", x"72", x"74", x"74", x"72", x"71", x"75", x"77", x"72", x"72", x"72", 
        x"6f", x"70", x"73", x"73", x"73", x"74", x"74", x"72", x"71", x"73", x"74", x"73", x"73", x"72", x"72", 
        x"71", x"71", x"71", x"73", x"74", x"73", x"74", x"73", x"72", x"71", x"73", x"72", x"70", x"6f", x"71", 
        x"73", x"71", x"6f", x"71", x"74", x"72", x"71", x"71", x"6f", x"71", x"72", x"73", x"72", x"71", x"70", 
        x"70", x"6f", x"73", x"75", x"72", x"71", x"70", x"76", x"74", x"71", x"72", x"72", x"70", x"72", x"71", 
        x"6e", x"70", x"6f", x"6e", x"6f", x"6f", x"71", x"71", x"70", x"71", x"73", x"71", x"72", x"73", x"6f", 
        x"70", x"71", x"73", x"73", x"72", x"70", x"70", x"73", x"71", x"6f", x"72", x"70", x"72", x"73", x"70", 
        x"6f", x"71", x"71", x"70", x"71", x"71", x"72", x"71", x"70", x"71", x"72", x"6e", x"6f", x"70", x"71", 
        x"6f", x"70", x"73", x"71", x"71", x"6e", x"6d", x"6f", x"6f", x"6d", x"6d", x"6e", x"6f", x"6e", x"6d", 
        x"6e", x"6e", x"6e", x"6d", x"6f", x"6c", x"6d", x"6e", x"6e", x"71", x"6d", x"6d", x"6e", x"6f", x"6f", 
        x"6f", x"6f", x"70", x"6c", x"6e", x"6f", x"6e", x"6e", x"6c", x"6c", x"6c", x"6b", x"6f", x"6f", x"6e", 
        x"6f", x"6c", x"6b", x"6d", x"6b", x"6d", x"70", x"6c", x"6b", x"6e", x"70", x"6e", x"6c", x"6e", x"6d", 
        x"6c", x"69", x"6d", x"6e", x"6e", x"6f", x"6f", x"70", x"6f", x"6a", x"6c", x"6f", x"6c", x"68", x"69", 
        x"6b", x"6b", x"6b", x"6a", x"69", x"6a", x"6a", x"6b", x"6b", x"69", x"6b", x"6d", x"6c", x"6f", x"70", 
        x"6a", x"6a", x"6c", x"6d", x"6d", x"6e", x"6c", x"67", x"6b", x"6f", x"6f", x"6d", x"6a", x"69", x"6b", 
        x"6c", x"6c", x"6d", x"6c", x"6c", x"6e", x"6f", x"6e", x"6c", x"6c", x"6b", x"6b", x"6b", x"6b", x"6c", 
        x"6b", x"6b", x"6f", x"69", x"6c", x"71", x"6d", x"6c", x"6b", x"6b", x"6c", x"6c", x"6b", x"69", x"68", 
        x"6a", x"6f", x"6c", x"6a", x"68", x"6a", x"6f", x"6c", x"6a", x"6b", x"6b", x"6a", x"6c", x"6a", x"68", 
        x"6d", x"6b", x"69", x"6a", x"6c", x"6d", x"6e", x"6b", x"6c", x"6c", x"6e", x"6b", x"6a", x"6a", x"67", 
        x"68", x"66", x"65", x"67", x"67", x"67", x"68", x"66", x"68", x"6a", x"68", x"6a", x"6b", x"6a", x"67", 
        x"67", x"69", x"69", x"6a", x"6c", x"6b", x"68", x"67", x"68", x"67", x"69", x"6b", x"69", x"69", x"6e", 
        x"6d", x"6b", x"6b", x"6b", x"6e", x"6d", x"69", x"6b", x"6d", x"6b", x"6a", x"6d", x"6d", x"6c", x"6a", 
        x"6a", x"6a", x"6c", x"6a", x"6c", x"6d", x"6e", x"6e", x"6e", x"6d", x"6c", x"6b", x"6c", x"6d", x"6c", 
        x"6d", x"6e", x"6d", x"6d", x"6a", x"6a", x"6c", x"6c", x"6d", x"6d", x"6b", x"6e", x"6d", x"6e", x"6b", 
        x"6c", x"6d", x"6d", x"6d", x"6c", x"6c", x"6c", x"6b", x"6b", x"6d", x"6a", x"69", x"6c", x"6e", x"6d", 
        x"6f", x"6e", x"6d", x"6a", x"6e", x"6e", x"6e", x"6f", x"6f", x"6f", x"6d", x"6f", x"6f", x"6f", x"70", 
        x"6e", x"70", x"6a", x"70", x"6f", x"6c", x"71", x"70", x"6e", x"6c", x"6e", x"70", x"6e", x"6e", x"71", 
        x"73", x"71", x"71", x"71", x"6f", x"6e", x"6f", x"70", x"6f", x"6f", x"6f", x"71", x"73", x"6e", x"69", 
        x"9a", x"db", x"d2", x"cf", x"cd", x"d0", x"d9", x"ce", x"cf", x"ce", x"cc", x"cd", x"ce", x"d0", x"d0", 
        x"cf", x"ce", x"cc", x"cb", x"cb", x"ce", x"cf", x"cf", x"cb", x"c9", x"cb", x"cd", x"cb", x"cb", x"cb", 
        x"cb", x"cc", x"cb", x"cd", x"cd", x"cd", x"cf", x"cf", x"cf", x"cf", x"ce", x"cd", x"cc", x"cb", x"cc", 
        x"cc", x"cc", x"cb", x"cb", x"ce", x"cf", x"ce", x"d5", x"d1", x"d3", x"d2", x"d1", x"d1", x"d0", x"ba", 
        x"7c", x"5f", x"5c", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5d", x"5e", x"5e", x"5c", x"6d", x"c6", x"f3", 
        x"f7", x"f9", x"f8", x"f7", x"f0", x"cf", x"98", x"6a", x"5a", x"5e", x"5e", x"5c", x"5d", x"5e", x"5d", 
        x"5c", x"5e", x"5e", x"5d", x"5c", x"5c", x"5c", x"5d", x"5d", x"5d", x"5f", x"5e", x"5c", x"5c", x"60", 
        x"60", x"5d", x"5d", x"5d", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"60", x"5f", x"76", x"d3", x"ec", 
        x"ee", x"ef", x"ee", x"ed", x"ee", x"ee", x"ed", x"ed", x"ee", x"f0", x"ef", x"ef", x"ed", x"ed", x"ed", 
        x"ed", x"ec", x"ea", x"e2", x"da", x"d6", x"d9", x"dd", x"e1", x"cd", x"ab", x"88", x"6e", x"6a", x"72", 
        x"78", x"78", x"76", x"76", x"79", x"77", x"73", x"75", x"77", x"78", x"7a", x"79", x"75", x"76", x"76", 
        x"77", x"77", x"77", x"77", x"78", x"78", x"78", x"77", x"76", x"77", x"77", x"76", x"76", x"76", x"77", 
        x"78", x"77", x"78", x"76", x"76", x"75", x"76", x"77", x"76", x"76", x"76", x"76", x"76", x"76", x"75", 
        x"75", x"76", x"78", x"79", x"79", x"78", x"78", x"77", x"75", x"73", x"76", x"76", x"75", x"74", x"75", 
        x"76", x"77", x"77", x"76", x"75", x"75", x"74", x"77", x"74", x"75", x"76", x"74", x"73", x"74", x"75", 
        x"74", x"74", x"74", x"74", x"75", x"76", x"75", x"75", x"76", x"76", x"75", x"75", x"77", x"75", x"75", 
        x"76", x"74", x"74", x"74", x"74", x"79", x"76", x"75", x"78", x"78", x"74", x"74", x"76", x"75", x"77", 
        x"78", x"75", x"75", x"74", x"72", x"72", x"73", x"75", x"75", x"74", x"73", x"75", x"74", x"72", x"74", 
        x"74", x"76", x"74", x"73", x"73", x"71", x"74", x"72", x"71", x"73", x"75", x"72", x"71", x"74", x"72", 
        x"72", x"75", x"75", x"72", x"75", x"75", x"75", x"75", x"73", x"73", x"72", x"72", x"72", x"73", x"74", 
        x"74", x"71", x"70", x"74", x"74", x"73", x"72", x"72", x"71", x"71", x"73", x"71", x"70", x"6f", x"70", 
        x"73", x"73", x"72", x"72", x"73", x"72", x"73", x"73", x"72", x"73", x"72", x"73", x"73", x"72", x"73", 
        x"72", x"71", x"72", x"73", x"72", x"73", x"72", x"73", x"73", x"73", x"74", x"74", x"72", x"72", x"71", 
        x"6e", x"6f", x"71", x"71", x"73", x"73", x"72", x"72", x"71", x"71", x"72", x"73", x"72", x"73", x"72", 
        x"72", x"72", x"71", x"71", x"72", x"73", x"71", x"73", x"74", x"73", x"71", x"6f", x"72", x"72", x"72", 
        x"72", x"71", x"71", x"72", x"71", x"70", x"70", x"72", x"73", x"74", x"72", x"6f", x"70", x"73", x"70", 
        x"6f", x"73", x"72", x"71", x"72", x"6e", x"6e", x"71", x"70", x"6d", x"6e", x"71", x"6f", x"6e", x"71", 
        x"70", x"70", x"72", x"70", x"71", x"70", x"6f", x"6e", x"70", x"70", x"6f", x"70", x"71", x"6f", x"6c", 
        x"6c", x"6e", x"70", x"6e", x"6e", x"6f", x"6d", x"6f", x"6d", x"6e", x"6f", x"6f", x"6e", x"6d", x"6e", 
        x"6f", x"6d", x"6b", x"6c", x"6a", x"6d", x"70", x"6e", x"6c", x"6d", x"70", x"6d", x"6d", x"6f", x"6e", 
        x"6c", x"6a", x"71", x"6f", x"6c", x"6d", x"6d", x"6a", x"6f", x"6e", x"6d", x"6e", x"6d", x"6c", x"6c", 
        x"6a", x"6c", x"6d", x"6b", x"6a", x"6b", x"6c", x"6d", x"6d", x"6a", x"6d", x"6e", x"6e", x"6e", x"6d", 
        x"6b", x"6b", x"6b", x"6d", x"6b", x"6c", x"6d", x"69", x"6b", x"6d", x"6d", x"6c", x"6a", x"6b", x"6c", 
        x"6d", x"6c", x"6d", x"6e", x"6c", x"6d", x"6b", x"6a", x"6c", x"6d", x"6c", x"6e", x"6e", x"6b", x"6c", 
        x"6d", x"6c", x"6d", x"6b", x"6a", x"6c", x"6c", x"6d", x"6c", x"6b", x"6c", x"6b", x"6b", x"69", x"6a", 
        x"6d", x"6f", x"6d", x"6a", x"6a", x"6c", x"6b", x"6b", x"6b", x"6b", x"6c", x"6a", x"6c", x"6d", x"6c", 
        x"6b", x"6a", x"6c", x"6d", x"6b", x"6a", x"6f", x"6b", x"6b", x"6d", x"6c", x"69", x"68", x"69", x"67", 
        x"65", x"65", x"66", x"66", x"66", x"66", x"68", x"68", x"68", x"6a", x"68", x"68", x"6b", x"6a", x"67", 
        x"67", x"69", x"68", x"69", x"6e", x"6d", x"6c", x"6d", x"6d", x"6b", x"6b", x"6b", x"68", x"66", x"6d", 
        x"6e", x"6b", x"6b", x"6c", x"6e", x"6e", x"69", x"6b", x"6e", x"6b", x"6c", x"6e", x"6b", x"6c", x"6c", 
        x"6d", x"68", x"69", x"69", x"6c", x"6c", x"6c", x"6c", x"6c", x"6c", x"6c", x"6c", x"6c", x"6c", x"6d", 
        x"6d", x"6d", x"6c", x"6b", x"6c", x"6c", x"6b", x"6b", x"6c", x"6d", x"6d", x"6c", x"6c", x"6e", x"6b", 
        x"6c", x"6d", x"6d", x"6f", x"6f", x"6f", x"6e", x"6d", x"6d", x"6d", x"6b", x"6b", x"6a", x"6d", x"6c", 
        x"6e", x"6d", x"6c", x"69", x"6e", x"70", x"6e", x"6e", x"6f", x"6f", x"6e", x"6f", x"70", x"72", x"72", 
        x"6f", x"6d", x"6d", x"74", x"71", x"6c", x"70", x"70", x"6d", x"6e", x"70", x"71", x"6f", x"6f", x"71", 
        x"72", x"70", x"70", x"72", x"6f", x"6e", x"6f", x"6f", x"6d", x"6c", x"6d", x"71", x"74", x"6f", x"6a", 
        x"99", x"db", x"d1", x"ce", x"cf", x"d2", x"d9", x"d0", x"d1", x"d0", x"ce", x"ce", x"cf", x"d0", x"d0", 
        x"ce", x"ce", x"cc", x"cb", x"cc", x"cf", x"cf", x"cf", x"cc", x"ca", x"cd", x"cf", x"ca", x"cb", x"cc", 
        x"cc", x"cc", x"cd", x"cd", x"cd", x"cd", x"cd", x"cf", x"cf", x"cf", x"ce", x"cd", x"cb", x"cb", x"cc", 
        x"cc", x"cb", x"ca", x"ca", x"cc", x"ce", x"d0", x"d8", x"cf", x"d2", x"d2", x"d1", x"d1", x"d1", x"bb", 
        x"7e", x"5f", x"5d", x"5f", x"60", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5d", x"64", x"9f", x"ea", 
        x"f8", x"f9", x"fb", x"f9", x"f9", x"f6", x"df", x"ab", x"6d", x"5c", x"61", x"5f", x"5d", x"5e", x"5e", 
        x"5b", x"5e", x"5f", x"5c", x"5b", x"5b", x"5c", x"5d", x"5a", x"5a", x"5c", x"5e", x"5d", x"5c", x"5d", 
        x"5c", x"5d", x"61", x"5f", x"5e", x"5f", x"5d", x"5d", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"5f", x"75", x"d2", x"ed", 
        x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ed", x"ee", x"ef", x"e9", x"dd", x"d3", x"cf", x"dd", x"e6", x"d7", x"b2", x"8d", x"71", 
        x"69", x"6f", x"77", x"7b", x"79", x"78", x"77", x"76", x"78", x"78", x"76", x"78", x"78", x"7c", x"77", 
        x"78", x"79", x"79", x"78", x"76", x"77", x"78", x"77", x"77", x"77", x"77", x"77", x"76", x"76", x"78", 
        x"7a", x"78", x"7a", x"76", x"77", x"76", x"76", x"76", x"75", x"76", x"76", x"77", x"77", x"77", x"78", 
        x"77", x"77", x"77", x"77", x"78", x"77", x"77", x"76", x"76", x"76", x"76", x"77", x"76", x"73", x"74", 
        x"75", x"76", x"76", x"75", x"75", x"76", x"76", x"78", x"75", x"77", x"76", x"75", x"75", x"75", x"75", 
        x"74", x"74", x"74", x"74", x"74", x"74", x"74", x"75", x"76", x"75", x"73", x"75", x"76", x"73", x"74", 
        x"76", x"74", x"76", x"79", x"75", x"76", x"73", x"74", x"77", x"76", x"73", x"72", x"75", x"74", x"74", 
        x"74", x"71", x"71", x"74", x"73", x"73", x"76", x"77", x"76", x"75", x"74", x"75", x"75", x"75", x"73", 
        x"73", x"74", x"73", x"75", x"74", x"73", x"76", x"73", x"73", x"75", x"76", x"73", x"74", x"74", x"72", 
        x"73", x"75", x"74", x"70", x"74", x"74", x"74", x"76", x"74", x"74", x"73", x"72", x"73", x"74", x"74", 
        x"73", x"71", x"71", x"75", x"73", x"72", x"71", x"70", x"71", x"73", x"74", x"72", x"72", x"70", x"72", 
        x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"74", x"72", x"72", x"73", x"72", x"75", 
        x"73", x"72", x"72", x"72", x"73", x"73", x"73", x"73", x"74", x"76", x"75", x"74", x"72", x"71", x"72", 
        x"70", x"71", x"72", x"71", x"72", x"73", x"72", x"72", x"72", x"72", x"73", x"74", x"72", x"71", x"71", 
        x"71", x"71", x"70", x"6f", x"71", x"72", x"70", x"72", x"74", x"73", x"71", x"72", x"73", x"6f", x"71", 
        x"72", x"6f", x"6f", x"71", x"70", x"70", x"73", x"74", x"73", x"73", x"71", x"6e", x"6e", x"74", x"72", 
        x"6f", x"74", x"73", x"70", x"73", x"71", x"72", x"73", x"70", x"6d", x"6e", x"70", x"71", x"70", x"73", 
        x"71", x"6f", x"71", x"70", x"70", x"71", x"6e", x"6d", x"6f", x"6e", x"6f", x"70", x"70", x"6e", x"6b", 
        x"6c", x"70", x"71", x"71", x"70", x"70", x"6f", x"70", x"6f", x"70", x"70", x"70", x"6e", x"6e", x"70", 
        x"70", x"6d", x"6c", x"6c", x"6a", x"6c", x"6e", x"6e", x"6d", x"6d", x"6f", x"6b", x"6c", x"71", x"6e", 
        x"6a", x"6c", x"72", x"6e", x"69", x"6b", x"6c", x"69", x"70", x"71", x"6e", x"6d", x"6e", x"6f", x"6e", 
        x"6c", x"6d", x"6e", x"6b", x"6a", x"6a", x"6b", x"6b", x"6c", x"6d", x"6f", x"70", x"6f", x"6d", x"6c", 
        x"6d", x"6e", x"6c", x"6e", x"6b", x"69", x"6c", x"69", x"6b", x"6b", x"6c", x"6d", x"6d", x"6d", x"6c", 
        x"6b", x"6b", x"6d", x"6d", x"6a", x"6b", x"6b", x"6a", x"6d", x"6d", x"6c", x"6e", x"6f", x"6d", x"6b", 
        x"6b", x"6b", x"6b", x"6c", x"6d", x"6f", x"6f", x"6f", x"6e", x"6c", x"6c", x"6a", x"6b", x"6a", x"6d", 
        x"6f", x"6d", x"6d", x"6a", x"6c", x"6c", x"6c", x"6e", x"6c", x"6a", x"6b", x"69", x"6a", x"6c", x"6e", 
        x"69", x"6a", x"6f", x"70", x"69", x"67", x"6d", x"6a", x"69", x"6a", x"6a", x"69", x"68", x"68", x"69", 
        x"68", x"6b", x"6c", x"67", x"68", x"69", x"68", x"66", x"66", x"6b", x"6c", x"6b", x"6d", x"6d", x"69", 
        x"68", x"69", x"69", x"6a", x"6e", x"6d", x"6d", x"6e", x"6f", x"6d", x"6c", x"6b", x"69", x"68", x"6d", 
        x"6e", x"6c", x"6c", x"6b", x"6b", x"6e", x"6b", x"6a", x"6c", x"6b", x"6b", x"6a", x"6b", x"6d", x"6e", 
        x"6e", x"68", x"69", x"6b", x"6d", x"6a", x"6a", x"6b", x"6b", x"6c", x"6d", x"6d", x"6b", x"6c", x"6e", 
        x"6e", x"6d", x"6c", x"6b", x"6e", x"6e", x"6c", x"6b", x"6b", x"6d", x"6e", x"70", x"6e", x"6e", x"6d", 
        x"6d", x"6c", x"6b", x"6e", x"6f", x"6f", x"6e", x"6d", x"6d", x"6d", x"6d", x"6e", x"6c", x"6c", x"6c", 
        x"6c", x"6b", x"6a", x"69", x"6d", x"6f", x"6f", x"6d", x"6d", x"6f", x"6c", x"6d", x"70", x"70", x"70", 
        x"6f", x"6e", x"6e", x"72", x"72", x"6e", x"70", x"70", x"6d", x"6e", x"72", x"73", x"71", x"70", x"71", 
        x"71", x"6f", x"6f", x"70", x"6f", x"6e", x"6f", x"71", x"71", x"6f", x"6f", x"73", x"72", x"6f", x"6a", 
        x"96", x"d8", x"d0", x"d0", x"d1", x"d2", x"d9", x"d0", x"cf", x"cf", x"ce", x"cf", x"cf", x"d0", x"cf", 
        x"cd", x"ce", x"cc", x"cc", x"ce", x"d0", x"ce", x"cd", x"cc", x"cc", x"cf", x"cd", x"c9", x"cb", x"ce", 
        x"ce", x"cd", x"cd", x"cd", x"cc", x"cc", x"cc", x"ce", x"cf", x"cf", x"ce", x"cd", x"cd", x"cd", x"ce", 
        x"cd", x"cc", x"cb", x"cc", x"cc", x"cd", x"d0", x"d8", x"ce", x"d0", x"d1", x"d2", x"d3", x"d2", x"bd", 
        x"7f", x"5f", x"5e", x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5d", x"5e", x"77", x"d2", 
        x"fa", x"f9", x"fa", x"fa", x"f9", x"f4", x"f6", x"e4", x"9d", x"63", x"5b", x"5e", x"5b", x"5d", x"60", 
        x"60", x"60", x"5d", x"5d", x"5f", x"5c", x"5d", x"5e", x"5d", x"5e", x"5f", x"5d", x"5b", x"59", x"5b", 
        x"5d", x"5c", x"5c", x"5c", x"5f", x"5d", x"5c", x"5e", x"5f", x"5f", x"5e", x"5e", x"5d", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"73", x"cf", x"ee", 
        x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"f0", x"f0", x"ed", x"eb", x"ed", x"ef", x"ea", x"e2", x"d1", x"c7", x"cf", x"e2", x"dc", x"c5", 
        x"98", x"72", x"65", x"71", x"78", x"7a", x"7b", x"79", x"77", x"79", x"7a", x"7b", x"77", x"77", x"76", 
        x"78", x"7a", x"7a", x"79", x"77", x"77", x"77", x"78", x"78", x"76", x"76", x"77", x"77", x"77", x"78", 
        x"7a", x"79", x"7a", x"77", x"78", x"79", x"77", x"75", x"75", x"76", x"77", x"78", x"78", x"79", x"79", 
        x"78", x"77", x"76", x"75", x"75", x"75", x"78", x"77", x"78", x"78", x"78", x"77", x"77", x"78", x"77", 
        x"76", x"75", x"76", x"78", x"79", x"78", x"76", x"76", x"74", x"76", x"76", x"76", x"79", x"76", x"75", 
        x"74", x"73", x"71", x"73", x"74", x"73", x"73", x"74", x"75", x"75", x"74", x"75", x"76", x"73", x"74", 
        x"75", x"74", x"77", x"7a", x"77", x"78", x"74", x"72", x"73", x"72", x"73", x"75", x"76", x"74", x"74", 
        x"74", x"73", x"74", x"75", x"75", x"75", x"76", x"76", x"77", x"75", x"75", x"75", x"75", x"75", x"73", 
        x"73", x"74", x"72", x"72", x"72", x"73", x"76", x"74", x"74", x"74", x"74", x"76", x"76", x"74", x"73", 
        x"74", x"74", x"74", x"72", x"74", x"73", x"73", x"73", x"71", x"75", x"75", x"74", x"74", x"74", x"74", 
        x"73", x"71", x"71", x"74", x"73", x"73", x"73", x"72", x"71", x"72", x"74", x"73", x"74", x"72", x"73", 
        x"74", x"71", x"72", x"73", x"74", x"74", x"73", x"73", x"73", x"74", x"72", x"73", x"74", x"72", x"74", 
        x"73", x"73", x"73", x"73", x"73", x"73", x"72", x"73", x"74", x"74", x"74", x"74", x"74", x"73", x"72", 
        x"71", x"74", x"74", x"70", x"70", x"73", x"73", x"71", x"71", x"73", x"74", x"74", x"71", x"70", x"70", 
        x"72", x"73", x"73", x"73", x"73", x"72", x"6f", x"72", x"72", x"72", x"73", x"75", x"73", x"6f", x"70", 
        x"71", x"71", x"71", x"71", x"6f", x"70", x"74", x"73", x"71", x"71", x"72", x"71", x"6f", x"75", x"75", 
        x"6f", x"72", x"72", x"70", x"71", x"6f", x"73", x"72", x"70", x"70", x"71", x"71", x"72", x"71", x"72", 
        x"6f", x"6f", x"71", x"70", x"70", x"71", x"6e", x"6d", x"6f", x"6e", x"71", x"70", x"70", x"70", x"6e", 
        x"6e", x"6f", x"6e", x"6d", x"6d", x"6f", x"6e", x"70", x"6d", x"6e", x"6e", x"70", x"70", x"70", x"6f", 
        x"70", x"6e", x"6e", x"6d", x"6c", x"6c", x"6e", x"6e", x"6e", x"6f", x"70", x"6b", x"6d", x"71", x"6c", 
        x"67", x"6b", x"72", x"70", x"6b", x"6c", x"6d", x"6c", x"70", x"70", x"6e", x"6e", x"6e", x"6f", x"6e", 
        x"6d", x"6c", x"6b", x"6b", x"6a", x"6a", x"6b", x"6d", x"6d", x"6a", x"6b", x"6d", x"6e", x"6f", x"6f", 
        x"6f", x"6e", x"6d", x"6e", x"6c", x"6b", x"6c", x"6a", x"6c", x"6c", x"6c", x"6d", x"6d", x"6d", x"6e", 
        x"6b", x"6c", x"6c", x"6b", x"6b", x"6b", x"6c", x"6d", x"6d", x"6d", x"6d", x"6e", x"6f", x"6e", x"6c", 
        x"6f", x"70", x"6d", x"6c", x"6e", x"6f", x"6d", x"6c", x"6c", x"6b", x"6b", x"6d", x"6e", x"6f", x"6e", 
        x"6d", x"6b", x"6c", x"6a", x"6c", x"6b", x"6b", x"6d", x"6c", x"6c", x"6e", x"6b", x"6b", x"6b", x"6b", 
        x"6d", x"6d", x"6b", x"6a", x"6c", x"6c", x"6a", x"69", x"69", x"6a", x"6b", x"6c", x"6d", x"6d", x"6c", 
        x"6c", x"6e", x"6e", x"69", x"69", x"6b", x"6c", x"6a", x"68", x"6d", x"6c", x"68", x"68", x"69", x"6d", 
        x"6b", x"6a", x"6b", x"6a", x"6b", x"69", x"6a", x"6b", x"6a", x"68", x"69", x"6b", x"6b", x"6a", x"6c", 
        x"6c", x"6a", x"6b", x"6b", x"6a", x"6b", x"6a", x"69", x"6b", x"6c", x"6f", x"70", x"6f", x"6d", x"6d", 
        x"6e", x"6c", x"6c", x"6c", x"6b", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6c", x"69", x"6a", x"6c", 
        x"6d", x"6d", x"6e", x"6e", x"6e", x"6d", x"6c", x"6b", x"6c", x"6d", x"6e", x"6f", x"6c", x"6c", x"6f", 
        x"70", x"6e", x"6f", x"6e", x"6d", x"6d", x"6d", x"6d", x"6d", x"6e", x"6e", x"6f", x"6d", x"6d", x"6e", 
        x"6f", x"6f", x"6e", x"6c", x"6d", x"6f", x"6f", x"6c", x"6c", x"6e", x"6d", x"6f", x"70", x"70", x"6f", 
        x"70", x"71", x"6d", x"6e", x"71", x"70", x"70", x"73", x"70", x"71", x"72", x"70", x"6e", x"71", x"73", 
        x"70", x"6d", x"6e", x"70", x"70", x"70", x"70", x"71", x"71", x"6e", x"6e", x"72", x"72", x"6f", x"6d", 
        x"96", x"d9", x"d2", x"d1", x"d0", x"d0", x"d6", x"cd", x"cd", x"ce", x"cf", x"cf", x"cf", x"cf", x"ce", 
        x"ce", x"ce", x"cd", x"cd", x"cf", x"d1", x"cf", x"ce", x"cd", x"cc", x"cf", x"ce", x"cb", x"cc", x"cd", 
        x"cc", x"cc", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"ce", x"cf", x"ce", x"ce", x"cf", x"cf", x"cf", 
        x"cd", x"cc", x"cc", x"cd", x"cd", x"cc", x"cf", x"d7", x"cf", x"d2", x"d2", x"d1", x"d1", x"d1", x"bf", 
        x"81", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5d", x"5d", x"66", x"a4", 
        x"ef", x"f7", x"f8", x"fb", x"f9", x"f8", x"f7", x"f6", x"e0", x"b1", x"82", x"69", x"5f", x"5d", x"5e", 
        x"5c", x"5d", x"5e", x"5c", x"5a", x"5c", x"5f", x"5e", x"5f", x"60", x"5d", x"5b", x"5c", x"5e", x"5d", 
        x"5d", x"5f", x"63", x"6c", x"71", x"73", x"69", x"60", x"5e", x"5d", x"5d", x"5e", x"5d", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"6f", x"cc", x"ee", 
        x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ef", x"ee", x"eb", x"ed", x"f1", x"ef", x"ed", x"ee", x"e7", x"d6", x"c6", x"cc", x"dd", 
        x"e3", x"d2", x"ad", x"81", x"71", x"73", x"75", x"77", x"79", x"7a", x"7c", x"7e", x"79", x"79", x"78", 
        x"79", x"79", x"79", x"78", x"79", x"79", x"78", x"79", x"78", x"76", x"75", x"76", x"77", x"78", x"77", 
        x"7a", x"7a", x"7b", x"77", x"78", x"77", x"77", x"76", x"75", x"76", x"78", x"79", x"78", x"77", x"77", 
        x"77", x"77", x"76", x"77", x"77", x"76", x"77", x"78", x"79", x"79", x"78", x"77", x"77", x"78", x"77", 
        x"76", x"75", x"76", x"77", x"78", x"77", x"76", x"76", x"75", x"76", x"76", x"76", x"76", x"75", x"74", 
        x"75", x"74", x"74", x"77", x"78", x"77", x"75", x"75", x"76", x"75", x"74", x"74", x"76", x"75", x"76", 
        x"77", x"74", x"74", x"75", x"76", x"77", x"76", x"75", x"74", x"74", x"76", x"76", x"75", x"73", x"75", 
        x"76", x"77", x"78", x"75", x"75", x"75", x"74", x"74", x"76", x"74", x"75", x"76", x"76", x"75", x"74", 
        x"74", x"74", x"72", x"71", x"72", x"74", x"76", x"74", x"74", x"73", x"75", x"76", x"76", x"74", x"73", 
        x"74", x"74", x"74", x"73", x"73", x"74", x"73", x"72", x"71", x"75", x"74", x"73", x"73", x"74", x"74", 
        x"73", x"73", x"72", x"73", x"73", x"74", x"74", x"73", x"71", x"72", x"73", x"72", x"73", x"72", x"72", 
        x"74", x"72", x"72", x"73", x"73", x"73", x"73", x"72", x"73", x"74", x"72", x"74", x"74", x"72", x"74", 
        x"72", x"72", x"72", x"73", x"74", x"74", x"73", x"73", x"73", x"73", x"74", x"76", x"75", x"73", x"72", 
        x"71", x"73", x"73", x"72", x"72", x"74", x"73", x"71", x"71", x"72", x"73", x"73", x"71", x"70", x"6f", 
        x"71", x"72", x"72", x"72", x"71", x"71", x"72", x"73", x"72", x"72", x"73", x"73", x"71", x"71", x"71", 
        x"71", x"72", x"73", x"73", x"71", x"70", x"74", x"74", x"70", x"71", x"74", x"72", x"70", x"74", x"75", 
        x"70", x"70", x"70", x"6f", x"71", x"72", x"74", x"73", x"71", x"70", x"70", x"70", x"71", x"71", x"71", 
        x"70", x"6f", x"6f", x"70", x"73", x"73", x"70", x"6e", x"70", x"70", x"72", x"6e", x"6d", x"6e", x"6f", 
        x"70", x"70", x"70", x"6c", x"6b", x"6d", x"6d", x"6d", x"6c", x"6d", x"6e", x"6f", x"6f", x"6e", x"6d", 
        x"6e", x"6f", x"70", x"6f", x"6d", x"6d", x"6d", x"6e", x"6e", x"6f", x"70", x"6d", x"6f", x"72", x"6d", 
        x"68", x"68", x"6f", x"6f", x"6c", x"6c", x"6e", x"6d", x"6d", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", 
        x"6c", x"6b", x"6b", x"6b", x"6b", x"69", x"6a", x"6c", x"6e", x"70", x"6e", x"6d", x"6e", x"6f", x"6f", 
        x"6d", x"6b", x"6b", x"6d", x"6e", x"6d", x"6e", x"6d", x"6f", x"6e", x"6c", x"6c", x"6c", x"6c", x"6c", 
        x"6b", x"6e", x"6d", x"6c", x"6d", x"6b", x"6c", x"6e", x"6b", x"6c", x"6e", x"6d", x"6f", x"6f", x"6c", 
        x"6e", x"6f", x"6d", x"6d", x"6f", x"6f", x"6f", x"6e", x"6d", x"6c", x"6a", x"6d", x"6b", x"6e", x"6e", 
        x"6d", x"69", x"6a", x"6a", x"6c", x"6b", x"6d", x"6d", x"6d", x"6d", x"6d", x"6a", x"67", x"6a", x"6b", 
        x"70", x"6e", x"6a", x"69", x"6e", x"6f", x"6a", x"69", x"6a", x"6a", x"6b", x"6c", x"6e", x"6e", x"6a", 
        x"6b", x"6b", x"69", x"69", x"68", x"69", x"6d", x"6a", x"68", x"6d", x"6c", x"67", x"66", x"68", x"6f", 
        x"6c", x"68", x"69", x"69", x"6b", x"6b", x"6b", x"6c", x"6b", x"69", x"6b", x"6c", x"6b", x"6a", x"6a", 
        x"6a", x"6a", x"6b", x"6f", x"6e", x"6d", x"6e", x"6c", x"6b", x"6b", x"6e", x"70", x"70", x"6a", x"6b", 
        x"6d", x"6b", x"6c", x"6e", x"6b", x"6d", x"6d", x"6d", x"6d", x"6e", x"6e", x"6d", x"6b", x"6a", x"6a", 
        x"6b", x"6c", x"6e", x"6e", x"6b", x"6b", x"6b", x"6c", x"6d", x"6d", x"6d", x"6f", x"6d", x"6c", x"6f", 
        x"70", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6f", x"6f", x"6f", x"6d", x"6c", x"6e", 
        x"70", x"70", x"6f", x"6f", x"6e", x"6f", x"6f", x"6d", x"6c", x"6d", x"6e", x"6f", x"6f", x"6e", x"6e", 
        x"70", x"73", x"6e", x"6d", x"71", x"71", x"70", x"73", x"71", x"71", x"71", x"6e", x"6c", x"6f", x"72", 
        x"71", x"70", x"71", x"72", x"72", x"71", x"6f", x"6e", x"6f", x"6e", x"6e", x"72", x"71", x"6f", x"6b", 
        x"93", x"d9", x"d1", x"d0", x"ce", x"cf", x"d6", x"ce", x"cd", x"ce", x"cf", x"d0", x"cf", x"ce", x"ce", 
        x"ce", x"ce", x"cd", x"cc", x"ce", x"d0", x"cf", x"d0", x"ce", x"cb", x"cd", x"d0", x"ce", x"cd", x"cb", 
        x"cb", x"cb", x"cc", x"cd", x"cd", x"ce", x"ce", x"ce", x"ce", x"cf", x"cf", x"cf", x"cf", x"cf", x"ce", 
        x"cc", x"cb", x"cc", x"cc", x"cc", x"cb", x"cd", x"d7", x"d0", x"d3", x"d3", x"d1", x"d0", x"d0", x"c1", 
        x"83", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5d", x"5c", x"5e", x"78", 
        x"cb", x"f6", x"f8", x"f8", x"f9", x"fa", x"f9", x"f8", x"f7", x"ee", x"d9", x"bb", x"9a", x"75", x"60", 
        x"5b", x"60", x"5e", x"5c", x"5e", x"5d", x"5f", x"5c", x"5e", x"5f", x"5c", x"5d", x"5f", x"68", x"71", 
        x"83", x"9f", x"b6", x"be", x"bc", x"ba", x"8e", x"64", x"5f", x"5f", x"5e", x"5f", x"5e", x"5f", x"5f", 
        x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5e", x"5e", x"6b", x"c6", x"ed", 
        x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ed", x"ec", x"ec", x"f0", x"ef", x"e8", x"da", x"cd", 
        x"cf", x"db", x"e2", x"d5", x"b2", x"89", x"6d", x"6d", x"74", x"78", x"77", x"79", x"7a", x"79", x"77", 
        x"79", x"78", x"78", x"78", x"79", x"7a", x"7a", x"7a", x"78", x"77", x"76", x"76", x"78", x"79", x"78", 
        x"7a", x"79", x"79", x"76", x"77", x"76", x"78", x"78", x"77", x"77", x"78", x"78", x"77", x"77", x"77", 
        x"77", x"77", x"77", x"77", x"78", x"77", x"76", x"77", x"78", x"78", x"77", x"76", x"76", x"78", x"78", 
        x"78", x"77", x"77", x"77", x"77", x"76", x"77", x"77", x"77", x"77", x"76", x"75", x"73", x"74", x"75", 
        x"75", x"75", x"77", x"77", x"76", x"76", x"75", x"75", x"75", x"76", x"74", x"75", x"76", x"76", x"76", 
        x"77", x"76", x"75", x"74", x"72", x"75", x"76", x"77", x"77", x"76", x"77", x"75", x"73", x"73", x"75", 
        x"76", x"77", x"75", x"73", x"75", x"75", x"73", x"73", x"75", x"74", x"76", x"76", x"75", x"75", x"75", 
        x"75", x"75", x"74", x"75", x"75", x"77", x"77", x"75", x"76", x"75", x"77", x"74", x"74", x"74", x"74", 
        x"74", x"74", x"73", x"73", x"73", x"75", x"76", x"75", x"75", x"75", x"74", x"73", x"74", x"75", x"76", 
        x"76", x"75", x"74", x"74", x"74", x"73", x"73", x"73", x"73", x"75", x"75", x"74", x"75", x"73", x"72", 
        x"75", x"75", x"73", x"73", x"73", x"73", x"73", x"73", x"74", x"75", x"73", x"74", x"74", x"73", x"74", 
        x"71", x"71", x"72", x"73", x"75", x"75", x"74", x"73", x"73", x"74", x"76", x"77", x"75", x"73", x"72", 
        x"72", x"71", x"72", x"74", x"75", x"74", x"75", x"74", x"73", x"73", x"74", x"75", x"74", x"73", x"72", 
        x"72", x"72", x"72", x"72", x"70", x"71", x"75", x"73", x"72", x"74", x"74", x"71", x"71", x"72", x"70", 
        x"6f", x"71", x"72", x"71", x"71", x"71", x"75", x"76", x"71", x"72", x"73", x"70", x"6f", x"73", x"73", 
        x"71", x"71", x"6e", x"6e", x"72", x"72", x"72", x"73", x"73", x"70", x"70", x"71", x"71", x"73", x"72", 
        x"71", x"6f", x"6d", x"6e", x"72", x"73", x"70", x"6f", x"70", x"6f", x"71", x"72", x"71", x"70", x"70", 
        x"6e", x"6d", x"6d", x"6d", x"6e", x"6f", x"6f", x"6d", x"6f", x"70", x"6e", x"6c", x"6f", x"6f", x"6e", 
        x"6d", x"6e", x"6f", x"6f", x"6f", x"6e", x"6d", x"6e", x"6e", x"6f", x"6e", x"6f", x"70", x"71", x"71", 
        x"6d", x"6a", x"6d", x"6d", x"6e", x"6d", x"6e", x"6d", x"6b", x"6c", x"6e", x"6e", x"6e", x"6e", x"6d", 
        x"6c", x"6b", x"6b", x"6c", x"6c", x"6c", x"6d", x"6f", x"70", x"70", x"6d", x"6c", x"6d", x"6e", x"6f", 
        x"6e", x"6d", x"6d", x"6e", x"6e", x"6e", x"6d", x"6d", x"6f", x"6e", x"6c", x"6c", x"6d", x"6d", x"6c", 
        x"6a", x"6d", x"6d", x"6e", x"6f", x"6d", x"6d", x"6f", x"6a", x"6b", x"6d", x"6c", x"6d", x"6e", x"6c", 
        x"6c", x"6b", x"6d", x"6e", x"6e", x"6f", x"70", x"6b", x"6a", x"6b", x"6a", x"6e", x"6e", x"71", x"6e", 
        x"6d", x"6a", x"6b", x"6b", x"6b", x"6a", x"6b", x"69", x"68", x"69", x"6b", x"6c", x"6d", x"6d", x"6a", 
        x"6f", x"6d", x"6d", x"6d", x"6d", x"6c", x"6c", x"6b", x"6b", x"6b", x"69", x"69", x"6a", x"6b", x"69", 
        x"6b", x"6b", x"69", x"6c", x"6a", x"6a", x"6d", x"67", x"68", x"6c", x"6b", x"69", x"69", x"69", x"6b", 
        x"6b", x"69", x"6b", x"6b", x"6a", x"6c", x"6e", x"6f", x"6f", x"6d", x"6d", x"6d", x"6b", x"6b", x"6c", 
        x"6c", x"6b", x"6b", x"70", x"6e", x"6f", x"73", x"71", x"6c", x"6b", x"6b", x"6d", x"6e", x"69", x"6c", 
        x"6c", x"68", x"69", x"71", x"6e", x"6a", x"6b", x"6d", x"6d", x"6e", x"6d", x"6d", x"6e", x"6b", x"69", 
        x"6a", x"6b", x"6c", x"6c", x"6a", x"6a", x"6b", x"6c", x"6d", x"6e", x"6d", x"6d", x"6e", x"6d", x"6e", 
        x"6e", x"6e", x"6f", x"70", x"71", x"71", x"70", x"6f", x"6e", x"6e", x"6f", x"6e", x"6d", x"6b", x"6d", 
        x"6c", x"6e", x"6e", x"70", x"70", x"6f", x"6f", x"6e", x"6e", x"6e", x"6e", x"6e", x"6d", x"6d", x"6e", 
        x"6f", x"71", x"70", x"6f", x"71", x"72", x"70", x"71", x"70", x"6f", x"71", x"70", x"6e", x"6d", x"6f", 
        x"71", x"72", x"72", x"72", x"73", x"72", x"6f", x"70", x"72", x"71", x"70", x"72", x"71", x"70", x"6a", 
        x"92", x"d7", x"d0", x"cf", x"cf", x"d1", x"d8", x"cf", x"cd", x"cf", x"d0", x"d0", x"cf", x"cf", x"ce", 
        x"cd", x"cf", x"cf", x"cc", x"cd", x"cf", x"d0", x"d0", x"cf", x"cc", x"cd", x"d0", x"d0", x"cd", x"cb", 
        x"cb", x"cb", x"cc", x"cd", x"cd", x"ce", x"ce", x"ce", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"cc", 
        x"cc", x"cc", x"cc", x"cc", x"cc", x"cc", x"cf", x"d8", x"cf", x"d2", x"d2", x"d1", x"d1", x"d1", x"c4", 
        x"85", x"5f", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5d", x"5c", x"5b", x"60", 
        x"99", x"e6", x"f9", x"f9", x"f9", x"f7", x"f8", x"fa", x"fa", x"f7", x"f8", x"f3", x"e5", x"c6", x"9c", 
        x"77", x"65", x"61", x"5d", x"5a", x"5d", x"60", x"58", x"59", x"67", x"71", x"7d", x"94", x"b3", x"ca", 
        x"db", x"ec", x"f4", x"eb", x"cf", x"b4", x"86", x"62", x"5d", x"5d", x"5e", x"5f", x"5e", x"5f", x"5f", 
        x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"5e", x"67", x"c1", x"ed", 
        x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ec", x"ec", x"ef", x"f0", x"eb", x"ea", x"ed", x"f0", x"ee", x"ea", 
        x"de", x"d0", x"cc", x"d6", x"e3", x"e0", x"be", x"8f", x"77", x"6f", x"6b", x"71", x"77", x"7c", x"7d", 
        x"7a", x"79", x"78", x"79", x"79", x"7a", x"7a", x"7a", x"79", x"78", x"78", x"77", x"78", x"79", x"7a", 
        x"7a", x"77", x"77", x"75", x"78", x"78", x"78", x"78", x"79", x"79", x"78", x"78", x"78", x"78", x"78", 
        x"78", x"77", x"77", x"78", x"78", x"77", x"77", x"77", x"78", x"77", x"77", x"77", x"77", x"78", x"78", 
        x"79", x"79", x"79", x"78", x"78", x"77", x"78", x"77", x"78", x"78", x"77", x"75", x"74", x"76", x"77", 
        x"76", x"75", x"77", x"75", x"73", x"73", x"72", x"73", x"75", x"76", x"76", x"77", x"76", x"76", x"75", 
        x"76", x"77", x"78", x"77", x"74", x"77", x"76", x"76", x"77", x"74", x"74", x"77", x"75", x"76", x"77", 
        x"77", x"77", x"73", x"74", x"75", x"75", x"74", x"73", x"74", x"75", x"76", x"76", x"75", x"75", x"76", 
        x"76", x"76", x"76", x"76", x"76", x"77", x"76", x"73", x"74", x"74", x"78", x"75", x"74", x"74", x"75", 
        x"75", x"75", x"74", x"74", x"73", x"75", x"77", x"74", x"74", x"76", x"75", x"74", x"75", x"77", x"78", 
        x"77", x"75", x"75", x"73", x"73", x"72", x"72", x"74", x"75", x"78", x"77", x"76", x"77", x"76", x"74", 
        x"76", x"76", x"74", x"73", x"73", x"73", x"73", x"74", x"74", x"75", x"73", x"74", x"75", x"73", x"75", 
        x"72", x"71", x"72", x"73", x"75", x"75", x"75", x"74", x"74", x"76", x"77", x"77", x"75", x"72", x"73", 
        x"74", x"71", x"71", x"76", x"76", x"73", x"74", x"74", x"73", x"73", x"73", x"74", x"74", x"74", x"74", 
        x"73", x"73", x"73", x"73", x"72", x"72", x"74", x"72", x"72", x"75", x"74", x"73", x"73", x"74", x"72", 
        x"72", x"73", x"72", x"72", x"73", x"71", x"73", x"75", x"74", x"74", x"74", x"70", x"71", x"73", x"72", 
        x"72", x"72", x"6f", x"70", x"72", x"72", x"72", x"74", x"75", x"72", x"72", x"73", x"70", x"72", x"72", 
        x"71", x"71", x"6e", x"6f", x"6f", x"71", x"6f", x"6e", x"70", x"6e", x"6f", x"71", x"6f", x"6f", x"70", 
        x"6f", x"6f", x"70", x"6e", x"6f", x"6f", x"70", x"6d", x"6f", x"71", x"6e", x"6a", x"6d", x"71", x"71", 
        x"6f", x"6d", x"6d", x"6f", x"6f", x"6e", x"6d", x"6e", x"6e", x"6e", x"6e", x"70", x"71", x"70", x"71", 
        x"6f", x"6a", x"6c", x"6c", x"6f", x"70", x"6d", x"6c", x"6c", x"6d", x"6d", x"6d", x"6d", x"6e", x"6d", 
        x"6c", x"6b", x"6c", x"6d", x"6e", x"6f", x"71", x"71", x"70", x"6c", x"6b", x"6b", x"6d", x"6e", x"70", 
        x"6f", x"6e", x"6f", x"6d", x"6e", x"6f", x"6d", x"6e", x"6e", x"6c", x"6b", x"6c", x"6f", x"6f", x"6d", 
        x"6a", x"6b", x"6e", x"6f", x"6f", x"6f", x"6f", x"6f", x"6c", x"6b", x"6c", x"6d", x"6d", x"6e", x"6f", 
        x"6e", x"6c", x"6d", x"6d", x"6c", x"6d", x"6e", x"6d", x"6c", x"6c", x"6a", x"6c", x"6c", x"6d", x"6c", 
        x"6d", x"6c", x"6d", x"6b", x"6b", x"6a", x"6c", x"6a", x"6b", x"6b", x"69", x"6a", x"6a", x"6c", x"6a", 
        x"6b", x"6e", x"6e", x"6b", x"6a", x"6c", x"6c", x"6a", x"6a", x"6b", x"69", x"68", x"69", x"6c", x"6c", 
        x"6b", x"6c", x"6d", x"6c", x"6c", x"6d", x"6c", x"6a", x"6b", x"6e", x"6b", x"69", x"6a", x"68", x"69", 
        x"6c", x"6a", x"6c", x"6b", x"69", x"6b", x"6c", x"6d", x"6d", x"6b", x"6c", x"6c", x"6b", x"6d", x"6d", 
        x"70", x"6d", x"6b", x"6f", x"6c", x"6b", x"70", x"6e", x"6c", x"6e", x"6d", x"6c", x"6e", x"6b", x"6e", 
        x"6e", x"6a", x"6b", x"72", x"6e", x"6c", x"6d", x"6f", x"6f", x"6e", x"6c", x"6c", x"6d", x"6a", x"68", 
        x"6b", x"6d", x"6c", x"6a", x"6e", x"6e", x"6d", x"6d", x"6e", x"6f", x"6f", x"6c", x"6e", x"6d", x"6d", 
        x"6d", x"6f", x"71", x"6e", x"6e", x"6e", x"6e", x"6d", x"6c", x"6c", x"6e", x"6f", x"70", x"6d", x"6d", 
        x"6c", x"6f", x"6f", x"6f", x"70", x"6f", x"6f", x"70", x"71", x"70", x"6f", x"6f", x"6f", x"70", x"71", 
        x"70", x"6f", x"6f", x"6e", x"70", x"71", x"71", x"71", x"72", x"70", x"72", x"73", x"71", x"6f", x"70", 
        x"6f", x"71", x"73", x"71", x"72", x"71", x"71", x"75", x"75", x"71", x"72", x"71", x"74", x"73", x"6c", 
        x"95", x"d7", x"cf", x"ce", x"d0", x"d2", x"d8", x"cc", x"ce", x"d0", x"d1", x"d0", x"cf", x"cf", x"cf", 
        x"cb", x"ce", x"d1", x"cf", x"cd", x"ce", x"cf", x"cf", x"d0", x"cf", x"ce", x"cf", x"cf", x"ce", x"cc", 
        x"cc", x"cc", x"cd", x"cd", x"cd", x"cd", x"cd", x"cf", x"cf", x"cf", x"cf", x"ce", x"cf", x"ce", x"cb", 
        x"cb", x"cc", x"cc", x"cc", x"cc", x"cd", x"cf", x"d8", x"cf", x"d1", x"d2", x"d1", x"d1", x"d1", x"c5", 
        x"86", x"5f", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5f", x"5e", x"5d", 
        x"6b", x"b7", x"ef", x"f9", x"f7", x"fa", x"fa", x"f9", x"fc", x"fa", x"f9", x"f7", x"f9", x"f9", x"ed", 
        x"d5", x"b8", x"9a", x"82", x"6a", x"58", x"65", x"7a", x"95", x"b4", x"cd", x"e4", x"ee", x"f7", x"f8", 
        x"f7", x"f4", x"e2", x"c4", x"93", x"6a", x"5e", x"5e", x"5f", x"5f", x"60", x"5f", x"5f", x"5f", x"5f", 
        x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"5e", x"62", x"be", x"ed", 
        x"ef", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ed", x"ec", x"ed", x"ed", x"ee", x"ef", x"ef", 
        x"f0", x"ee", x"ed", x"ee", x"ef", x"ef", x"ed", x"ed", x"ed", x"ec", x"ed", x"ee", x"ec", x"eb", x"ee", 
        x"ef", x"ec", x"e5", x"d7", x"cf", x"d7", x"e0", x"e4", x"cf", x"a5", x"7a", x"6d", x"6e", x"72", x"77", 
        x"7c", x"7b", x"7a", x"7b", x"7a", x"78", x"77", x"7a", x"7a", x"7a", x"79", x"7a", x"79", x"79", x"7b", 
        x"7a", x"76", x"78", x"79", x"7c", x"7a", x"78", x"78", x"7a", x"79", x"78", x"77", x"7a", x"7a", x"79", 
        x"78", x"78", x"78", x"78", x"79", x"79", x"79", x"78", x"78", x"77", x"78", x"79", x"78", x"76", x"77", 
        x"78", x"78", x"78", x"78", x"78", x"77", x"78", x"76", x"77", x"76", x"76", x"77", x"76", x"77", x"78", 
        x"79", x"78", x"76", x"75", x"76", x"76", x"75", x"74", x"76", x"78", x"78", x"77", x"77", x"77", x"76", 
        x"77", x"78", x"78", x"77", x"77", x"79", x"76", x"75", x"78", x"77", x"75", x"79", x"76", x"78", x"79", 
        x"79", x"79", x"75", x"77", x"77", x"77", x"77", x"74", x"74", x"76", x"77", x"74", x"73", x"74", x"77", 
        x"78", x"78", x"77", x"76", x"75", x"77", x"74", x"73", x"75", x"72", x"76", x"78", x"75", x"72", x"75", 
        x"76", x"74", x"74", x"76", x"72", x"74", x"75", x"72", x"72", x"77", x"77", x"76", x"76", x"77", x"77", 
        x"77", x"73", x"74", x"73", x"73", x"71", x"71", x"76", x"74", x"75", x"74", x"74", x"76", x"75", x"74", 
        x"75", x"74", x"74", x"74", x"75", x"75", x"75", x"74", x"75", x"75", x"73", x"73", x"74", x"73", x"76", 
        x"75", x"74", x"73", x"73", x"73", x"74", x"74", x"74", x"76", x"77", x"76", x"75", x"73", x"73", x"74", 
        x"77", x"75", x"73", x"75", x"72", x"71", x"74", x"73", x"73", x"74", x"75", x"75", x"73", x"73", x"74", 
        x"72", x"71", x"72", x"74", x"74", x"73", x"73", x"73", x"73", x"73", x"74", x"74", x"73", x"72", x"71", 
        x"73", x"74", x"73", x"70", x"72", x"72", x"72", x"74", x"74", x"74", x"73", x"71", x"72", x"75", x"74", 
        x"73", x"73", x"74", x"74", x"73", x"75", x"75", x"75", x"73", x"73", x"72", x"70", x"70", x"73", x"70", 
        x"71", x"72", x"70", x"72", x"6d", x"6f", x"6e", x"70", x"72", x"70", x"70", x"72", x"6f", x"6f", x"71", 
        x"6f", x"6e", x"6f", x"6e", x"6f", x"71", x"73", x"6f", x"71", x"72", x"70", x"6c", x"6e", x"6f", x"70", 
        x"70", x"6f", x"6e", x"6d", x"70", x"70", x"6d", x"6d", x"6d", x"6d", x"6f", x"6e", x"6e", x"6f", x"6f", 
        x"6e", x"6d", x"6f", x"6d", x"70", x"70", x"6b", x"6d", x"70", x"6f", x"6e", x"6d", x"6e", x"6f", x"6e", 
        x"6c", x"6d", x"6f", x"6e", x"6e", x"6e", x"6d", x"6c", x"6d", x"70", x"70", x"6f", x"6d", x"6c", x"6d", 
        x"6d", x"6d", x"6e", x"6c", x"6e", x"6f", x"6e", x"70", x"6f", x"6c", x"6c", x"6d", x"6f", x"6f", x"6d", 
        x"6e", x"6d", x"6f", x"6f", x"6d", x"6d", x"6e", x"6f", x"6f", x"6c", x"6d", x"70", x"6e", x"6e", x"70", 
        x"6d", x"6d", x"6d", x"6d", x"6e", x"6f", x"6e", x"6b", x"6b", x"6b", x"6d", x"6b", x"6d", x"6c", x"6b", 
        x"6e", x"6e", x"6f", x"6c", x"6b", x"6a", x"6b", x"6a", x"6d", x"6c", x"69", x"6c", x"6d", x"6e", x"6a", 
        x"6c", x"6e", x"6d", x"6b", x"69", x"6d", x"69", x"68", x"69", x"6a", x"69", x"69", x"6b", x"6e", x"6d", 
        x"6a", x"6b", x"6c", x"6b", x"6b", x"69", x"68", x"6a", x"6c", x"6c", x"6c", x"6b", x"6a", x"6a", x"69", 
        x"6b", x"6b", x"6c", x"6d", x"6d", x"6e", x"6b", x"6a", x"69", x"6a", x"6b", x"6c", x"6b", x"6c", x"6d", 
        x"6f", x"6d", x"6c", x"6e", x"6b", x"6c", x"6e", x"6d", x"6c", x"6e", x"6d", x"6a", x"6e", x"6d", x"6e", 
        x"6f", x"6e", x"6e", x"70", x"6c", x"6d", x"6d", x"6e", x"70", x"6e", x"6d", x"6c", x"6c", x"6a", x"6a", 
        x"6c", x"6d", x"6d", x"6d", x"6e", x"70", x"6f", x"6d", x"6e", x"6f", x"6e", x"6d", x"70", x"6e", x"6a", 
        x"68", x"6a", x"6c", x"6a", x"6c", x"6d", x"6d", x"6c", x"6c", x"6d", x"6d", x"6d", x"6f", x"6f", x"70", 
        x"6e", x"71", x"71", x"71", x"70", x"70", x"70", x"71", x"71", x"6e", x"6f", x"6f", x"70", x"6f", x"6e", 
        x"6f", x"6f", x"71", x"71", x"71", x"70", x"70", x"70", x"72", x"72", x"72", x"71", x"72", x"72", x"70", 
        x"6e", x"71", x"73", x"71", x"71", x"72", x"70", x"73", x"74", x"73", x"74", x"72", x"73", x"73", x"6b", 
        x"92", x"d8", x"d1", x"cf", x"d0", x"d1", x"d7", x"cf", x"cd", x"cf", x"d0", x"cf", x"ce", x"ce", x"cf", 
        x"cd", x"ce", x"d0", x"cf", x"ce", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"ce", x"cf", x"cf", x"cd", 
        x"cc", x"cc", x"cc", x"ce", x"ce", x"ce", x"cd", x"ce", x"ce", x"cf", x"cf", x"cf", x"cf", x"ce", x"cc", 
        x"cc", x"cd", x"cd", x"cc", x"cc", x"cd", x"cf", x"d9", x"cc", x"d1", x"d3", x"d1", x"cf", x"d1", x"c4", 
        x"85", x"5d", x"5e", x"5e", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", 
        x"5b", x"80", x"c0", x"ee", x"f6", x"f9", x"f9", x"f7", x"f9", x"fb", x"f9", x"fb", x"fc", x"fb", x"f9", 
        x"f8", x"f3", x"e4", x"ca", x"9d", x"89", x"a7", x"cd", x"e7", x"f4", x"f8", x"fa", x"f8", x"f4", x"e6", 
        x"d1", x"b7", x"98", x"76", x"63", x"5c", x"5f", x"60", x"5e", x"5d", x"5f", x"5e", x"61", x"60", x"5f", 
        x"5f", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"5e", x"60", x"bd", x"ec", 
        x"ee", x"ed", x"ec", x"ed", x"ed", x"ed", x"ee", x"ed", x"ed", x"ec", x"ed", x"ed", x"ee", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ef", x"ec", x"eb", x"ec", 
        x"ec", x"f0", x"f2", x"ed", x"e5", x"d9", x"d0", x"d1", x"d8", x"df", x"cf", x"af", x"8d", x"73", x"6c", 
        x"72", x"7a", x"7a", x"7a", x"7a", x"78", x"78", x"79", x"79", x"79", x"7a", x"7a", x"79", x"78", x"7c", 
        x"79", x"76", x"7a", x"7b", x"7b", x"7a", x"79", x"79", x"7a", x"79", x"78", x"78", x"79", x"79", x"78", 
        x"78", x"78", x"78", x"78", x"79", x"7a", x"7b", x"79", x"78", x"78", x"76", x"76", x"77", x"77", x"77", 
        x"78", x"78", x"7a", x"7a", x"7a", x"78", x"77", x"76", x"76", x"76", x"77", x"77", x"79", x"78", x"76", 
        x"78", x"78", x"77", x"79", x"7a", x"79", x"77", x"78", x"78", x"78", x"78", x"77", x"78", x"79", x"79", 
        x"79", x"79", x"78", x"75", x"78", x"7a", x"77", x"77", x"7a", x"7a", x"77", x"76", x"75", x"77", x"77", 
        x"76", x"76", x"75", x"76", x"77", x"78", x"78", x"75", x"76", x"77", x"76", x"75", x"75", x"76", x"78", 
        x"78", x"77", x"77", x"77", x"74", x"75", x"75", x"75", x"76", x"74", x"75", x"77", x"74", x"72", x"75", 
        x"76", x"73", x"73", x"74", x"71", x"74", x"78", x"74", x"73", x"76", x"77", x"76", x"76", x"76", x"77", 
        x"77", x"74", x"75", x"74", x"74", x"72", x"73", x"78", x"75", x"73", x"74", x"73", x"74", x"74", x"74", 
        x"75", x"73", x"74", x"76", x"76", x"77", x"75", x"75", x"76", x"74", x"73", x"74", x"75", x"75", x"73", 
        x"76", x"76", x"74", x"74", x"76", x"74", x"72", x"72", x"73", x"74", x"74", x"74", x"74", x"76", x"75", 
        x"76", x"76", x"74", x"74", x"72", x"73", x"75", x"75", x"73", x"74", x"75", x"75", x"74", x"73", x"73", 
        x"73", x"73", x"72", x"75", x"77", x"75", x"73", x"73", x"74", x"74", x"75", x"74", x"70", x"71", x"71", 
        x"72", x"72", x"71", x"70", x"72", x"73", x"73", x"73", x"75", x"75", x"73", x"73", x"73", x"76", x"74", 
        x"72", x"76", x"76", x"73", x"73", x"73", x"74", x"73", x"73", x"74", x"75", x"73", x"71", x"72", x"70", 
        x"72", x"72", x"70", x"71", x"70", x"71", x"70", x"71", x"72", x"70", x"70", x"70", x"6f", x"70", x"72", 
        x"71", x"70", x"70", x"6f", x"71", x"73", x"74", x"71", x"71", x"71", x"71", x"6e", x"6e", x"6f", x"6f", 
        x"6f", x"6f", x"6f", x"6e", x"70", x"70", x"6f", x"6e", x"6d", x"6c", x"6e", x"6e", x"6d", x"6f", x"70", 
        x"6d", x"6e", x"72", x"70", x"6f", x"70", x"6e", x"6d", x"71", x"70", x"6d", x"6b", x"6b", x"6c", x"6d", 
        x"6a", x"6c", x"70", x"6e", x"6c", x"6f", x"71", x"6d", x"6d", x"6f", x"6e", x"6d", x"6c", x"6d", x"6c", 
        x"6c", x"6e", x"6f", x"6f", x"6f", x"70", x"6e", x"70", x"6e", x"6c", x"6c", x"6f", x"71", x"6f", x"6c", 
        x"6d", x"6f", x"71", x"6f", x"6c", x"6d", x"6e", x"70", x"70", x"6d", x"6d", x"6f", x"6e", x"6c", x"6d", 
        x"6d", x"6f", x"6e", x"6d", x"6f", x"6d", x"6e", x"6d", x"6d", x"6b", x"6d", x"6d", x"6e", x"6d", x"6d", 
        x"6e", x"6e", x"6e", x"6c", x"6d", x"6d", x"6e", x"6d", x"6d", x"6d", x"6b", x"6c", x"6c", x"6d", x"6c", 
        x"71", x"6d", x"6e", x"70", x"6b", x"6e", x"6a", x"69", x"6a", x"6a", x"69", x"69", x"6b", x"6e", x"6e", 
        x"6c", x"6c", x"6d", x"6d", x"6c", x"6a", x"69", x"6b", x"6a", x"68", x"6b", x"6b", x"6a", x"6c", x"6b", 
        x"6b", x"6d", x"6f", x"71", x"71", x"6f", x"6d", x"6b", x"6b", x"6d", x"6c", x"6b", x"6b", x"6d", x"6f", 
        x"6e", x"6c", x"6e", x"6f", x"6b", x"6c", x"6c", x"6b", x"6c", x"6e", x"6e", x"6c", x"6c", x"6d", x"6c", 
        x"6e", x"70", x"6e", x"6f", x"6e", x"6c", x"6a", x"6b", x"6e", x"6c", x"6e", x"6d", x"6d", x"6c", x"6d", 
        x"6d", x"6c", x"6d", x"70", x"6d", x"71", x"71", x"6e", x"6e", x"70", x"6e", x"6c", x"6e", x"6d", x"69", 
        x"69", x"6d", x"6e", x"6c", x"6e", x"70", x"6f", x"6d", x"6d", x"6f", x"6e", x"6c", x"6f", x"72", x"71", 
        x"6f", x"70", x"72", x"71", x"6f", x"71", x"70", x"70", x"71", x"6e", x"70", x"71", x"73", x"70", x"6e", 
        x"71", x"72", x"73", x"73", x"72", x"70", x"6e", x"6f", x"71", x"72", x"6f", x"6e", x"72", x"72", x"6f", 
        x"6e", x"71", x"70", x"70", x"71", x"72", x"70", x"71", x"71", x"72", x"74", x"72", x"72", x"74", x"6c", 
        x"8f", x"d8", x"d3", x"ce", x"ce", x"cf", x"d8", x"d3", x"cc", x"cd", x"cf", x"ce", x"ce", x"ce", x"ce", 
        x"d0", x"d0", x"ce", x"cf", x"d0", x"d1", x"d0", x"d0", x"cd", x"ce", x"cf", x"ce", x"cf", x"ce", x"cc", 
        x"cd", x"cc", x"cd", x"cf", x"d1", x"d0", x"ce", x"cd", x"cd", x"ce", x"d0", x"cf", x"cf", x"ce", x"cf", 
        x"cf", x"cf", x"cf", x"ce", x"ce", x"cd", x"ca", x"d9", x"cc", x"d0", x"d2", x"d2", x"d1", x"d3", x"c3", 
        x"84", x"5e", x"5e", x"5c", x"5c", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"60", x"5f", 
        x"5d", x"5d", x"7b", x"bc", x"ec", x"f9", x"fa", x"f8", x"fb", x"fc", x"fb", x"fa", x"fc", x"fc", x"f9", 
        x"fb", x"fb", x"f9", x"f0", x"dc", x"db", x"ef", x"fa", x"fc", x"fd", x"fa", x"f3", x"da", x"b8", x"94", 
        x"7d", x"6a", x"5c", x"5a", x"5d", x"60", x"61", x"5f", x"5e", x"5d", x"5b", x"5a", x"5d", x"5c", x"5e", 
        x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5f", x"bd", x"ec", 
        x"ee", x"ec", x"ec", x"ec", x"ec", x"ec", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ee", x"ed", x"ef", x"ef", x"e8", x"d9", x"cd", x"cb", x"d8", x"e5", x"de", x"ba", x"98", 
        x"78", x"68", x"6e", x"79", x"7a", x"79", x"79", x"7c", x"79", x"77", x"7a", x"7d", x"7c", x"79", x"7b", 
        x"78", x"77", x"7a", x"7b", x"79", x"7a", x"7c", x"7b", x"7a", x"79", x"78", x"78", x"79", x"78", x"79", 
        x"7b", x"7b", x"7a", x"79", x"7a", x"7a", x"79", x"77", x"78", x"7a", x"75", x"76", x"76", x"78", x"77", 
        x"76", x"78", x"79", x"7a", x"7a", x"78", x"78", x"78", x"78", x"78", x"79", x"79", x"7b", x"78", x"77", 
        x"79", x"79", x"78", x"79", x"79", x"79", x"78", x"78", x"78", x"77", x"75", x"74", x"76", x"78", x"78", 
        x"77", x"79", x"78", x"76", x"78", x"78", x"78", x"77", x"77", x"77", x"77", x"76", x"77", x"78", x"76", 
        x"74", x"73", x"75", x"74", x"75", x"76", x"77", x"73", x"76", x"75", x"73", x"75", x"75", x"76", x"77", 
        x"78", x"78", x"76", x"76", x"74", x"72", x"77", x"77", x"74", x"75", x"76", x"75", x"73", x"73", x"76", 
        x"75", x"73", x"74", x"76", x"72", x"74", x"79", x"76", x"75", x"78", x"77", x"76", x"74", x"74", x"76", 
        x"78", x"77", x"77", x"77", x"76", x"76", x"76", x"77", x"76", x"74", x"74", x"74", x"75", x"75", x"74", 
        x"75", x"75", x"76", x"76", x"75", x"76", x"74", x"76", x"76", x"71", x"73", x"74", x"74", x"74", x"6f", 
        x"73", x"76", x"73", x"74", x"77", x"75", x"72", x"71", x"71", x"71", x"72", x"73", x"75", x"76", x"76", 
        x"74", x"73", x"73", x"73", x"73", x"72", x"74", x"76", x"73", x"74", x"75", x"73", x"76", x"74", x"73", 
        x"74", x"74", x"72", x"74", x"78", x"76", x"74", x"73", x"73", x"75", x"74", x"71", x"6e", x"72", x"73", 
        x"72", x"72", x"72", x"72", x"74", x"75", x"73", x"73", x"75", x"75", x"73", x"74", x"74", x"74", x"73", 
        x"70", x"76", x"73", x"70", x"73", x"73", x"75", x"75", x"75", x"75", x"74", x"73", x"70", x"70", x"72", 
        x"73", x"74", x"73", x"71", x"73", x"73", x"73", x"71", x"70", x"6f", x"6e", x"71", x"72", x"72", x"72", 
        x"72", x"71", x"6f", x"6f", x"70", x"72", x"71", x"6f", x"6e", x"6f", x"6f", x"6f", x"6f", x"6f", x"6e", 
        x"6e", x"6e", x"6e", x"70", x"71", x"70", x"71", x"6f", x"6e", x"6c", x"6d", x"6f", x"6d", x"70", x"72", 
        x"70", x"70", x"74", x"73", x"6d", x"6e", x"71", x"6f", x"70", x"70", x"6b", x"68", x"68", x"69", x"69", 
        x"68", x"6c", x"72", x"6e", x"6a", x"70", x"72", x"6c", x"6c", x"6f", x"6d", x"6d", x"6d", x"70", x"6c", 
        x"6c", x"6d", x"6e", x"70", x"6e", x"6f", x"6f", x"70", x"6f", x"6c", x"6c", x"71", x"72", x"6e", x"6c", 
        x"6b", x"6e", x"70", x"6d", x"6b", x"6d", x"6f", x"70", x"6e", x"6d", x"6d", x"6e", x"6e", x"6b", x"6a", 
        x"69", x"6c", x"6d", x"6b", x"6d", x"6a", x"6e", x"6e", x"6d", x"6c", x"6d", x"6f", x"6f", x"6f", x"6e", 
        x"6d", x"6c", x"6c", x"6c", x"6e", x"6e", x"6d", x"6f", x"6e", x"6e", x"70", x"6d", x"6b", x"6a", x"6a", 
        x"71", x"6c", x"6c", x"6c", x"69", x"6c", x"69", x"69", x"6c", x"6c", x"6a", x"68", x"69", x"6c", x"6b", 
        x"69", x"69", x"68", x"69", x"6a", x"6b", x"6c", x"6e", x"6e", x"6d", x"6f", x"70", x"70", x"70", x"6d", 
        x"6d", x"6d", x"6d", x"6d", x"6e", x"6d", x"6a", x"6d", x"6f", x"6e", x"6c", x"6b", x"6c", x"6c", x"6e", 
        x"6e", x"6b", x"6b", x"6b", x"6b", x"6c", x"6d", x"6d", x"6e", x"6e", x"6f", x"6e", x"6d", x"6b", x"6b", 
        x"6c", x"6d", x"6e", x"70", x"72", x"70", x"6e", x"6f", x"70", x"6d", x"70", x"70", x"6e", x"6c", x"6c", 
        x"6d", x"6d", x"6e", x"70", x"6f", x"6f", x"6d", x"6c", x"6d", x"6f", x"6e", x"6d", x"6f", x"70", x"6e", 
        x"6e", x"6e", x"6e", x"6d", x"6e", x"6f", x"6f", x"6e", x"6e", x"6f", x"6f", x"6e", x"6e", x"6f", x"6e", 
        x"6b", x"6c", x"6f", x"73", x"70", x"70", x"6f", x"70", x"71", x"6e", x"6c", x"6d", x"72", x"72", x"6f", 
        x"70", x"6f", x"6f", x"70", x"72", x"72", x"72", x"71", x"72", x"72", x"71", x"72", x"74", x"74", x"72", 
        x"73", x"73", x"71", x"70", x"73", x"74", x"73", x"73", x"73", x"72", x"73", x"70", x"72", x"74", x"6b", 
        x"8e", x"d8", x"d2", x"ce", x"ce", x"cf", x"d8", x"d3", x"cc", x"cd", x"cf", x"ce", x"ce", x"ce", x"ce", 
        x"d0", x"d0", x"cf", x"cf", x"d1", x"d1", x"d0", x"d0", x"cd", x"cd", x"ce", x"ce", x"ce", x"cd", x"cc", 
        x"cd", x"cd", x"cd", x"cf", x"d0", x"d0", x"cf", x"ce", x"ce", x"cf", x"d0", x"cf", x"ce", x"cd", x"ce", 
        x"cf", x"cf", x"cf", x"ce", x"ce", x"cd", x"cd", x"d5", x"cb", x"d3", x"d2", x"d2", x"d1", x"d4", x"c2", 
        x"84", x"5e", x"5c", x"5d", x"5d", x"5c", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"5f", x"5e", 
        x"60", x"5a", x"5b", x"70", x"b5", x"e4", x"f7", x"f9", x"f6", x"f9", x"fa", x"fa", x"fa", x"fc", x"fa", 
        x"fa", x"fc", x"fb", x"fa", x"f9", x"fa", x"fa", x"f5", x"f8", x"fc", x"fa", x"f3", x"d0", x"9c", x"6a", 
        x"5b", x"5b", x"5b", x"5c", x"5e", x"5c", x"59", x"5c", x"5e", x"5c", x"6a", x"73", x"6f", x"6a", x"6d", 
        x"71", x"63", x"5c", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"b8", x"eb", 
        x"ee", x"ec", x"ec", x"ec", x"ed", x"ed", x"ed", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"ee", x"ed", x"ee", x"ef", x"ed", x"ee", x"ed", x"e9", x"e5", x"d6", x"ca", x"cb", x"de", x"e7", 
        x"d0", x"a9", x"80", x"6a", x"6d", x"78", x"7b", x"7b", x"7b", x"7a", x"79", x"79", x"7a", x"7c", x"7a", 
        x"79", x"7a", x"7a", x"7a", x"7c", x"7d", x"7b", x"7a", x"7a", x"79", x"79", x"7a", x"7c", x"7a", x"7a", 
        x"7b", x"7b", x"7a", x"7a", x"7a", x"7b", x"7b", x"7a", x"7a", x"7c", x"77", x"78", x"77", x"79", x"78", 
        x"78", x"78", x"79", x"79", x"78", x"79", x"79", x"7b", x"7c", x"7b", x"7a", x"79", x"78", x"78", x"79", 
        x"7b", x"7a", x"77", x"76", x"76", x"76", x"76", x"76", x"77", x"77", x"78", x"78", x"78", x"7a", x"7a", 
        x"79", x"7a", x"79", x"77", x"76", x"77", x"78", x"77", x"77", x"78", x"79", x"78", x"79", x"79", x"78", 
        x"76", x"76", x"77", x"76", x"77", x"76", x"78", x"77", x"79", x"75", x"76", x"78", x"77", x"77", x"77", 
        x"78", x"78", x"76", x"76", x"75", x"75", x"78", x"78", x"76", x"77", x"77", x"75", x"75", x"76", x"76", 
        x"76", x"76", x"75", x"77", x"75", x"74", x"74", x"73", x"76", x"75", x"74", x"75", x"76", x"76", x"77", 
        x"77", x"75", x"74", x"74", x"74", x"74", x"74", x"74", x"76", x"76", x"74", x"75", x"77", x"77", x"75", 
        x"74", x"74", x"75", x"75", x"74", x"76", x"76", x"78", x"77", x"73", x"74", x"74", x"75", x"75", x"72", 
        x"71", x"74", x"71", x"71", x"74", x"74", x"73", x"72", x"73", x"75", x"74", x"74", x"74", x"75", x"76", 
        x"75", x"75", x"74", x"74", x"74", x"73", x"73", x"75", x"74", x"75", x"76", x"75", x"77", x"75", x"76", 
        x"75", x"74", x"74", x"74", x"74", x"75", x"73", x"74", x"75", x"73", x"72", x"72", x"72", x"73", x"74", 
        x"73", x"74", x"74", x"74", x"74", x"76", x"76", x"75", x"74", x"73", x"70", x"70", x"72", x"73", x"74", 
        x"73", x"74", x"73", x"72", x"73", x"73", x"75", x"75", x"75", x"74", x"74", x"74", x"70", x"70", x"72", 
        x"73", x"74", x"72", x"71", x"74", x"74", x"74", x"73", x"72", x"71", x"71", x"70", x"70", x"70", x"71", 
        x"73", x"73", x"72", x"70", x"6f", x"6f", x"70", x"70", x"71", x"71", x"70", x"6f", x"70", x"6d", x"6c", 
        x"6f", x"70", x"6f", x"70", x"71", x"70", x"70", x"6e", x"6f", x"6f", x"71", x"6f", x"6e", x"6e", x"6f", 
        x"70", x"6f", x"70", x"6e", x"6b", x"6d", x"70", x"6e", x"6f", x"70", x"6f", x"6e", x"6d", x"6e", x"6e", 
        x"6e", x"6f", x"71", x"6d", x"6c", x"71", x"73", x"6f", x"6c", x"6d", x"6e", x"6f", x"6f", x"70", x"6c", 
        x"6c", x"6f", x"6e", x"6e", x"6d", x"6f", x"6f", x"71", x"73", x"70", x"6e", x"6f", x"6f", x"6d", x"6c", 
        x"6d", x"70", x"70", x"6e", x"6d", x"6d", x"6e", x"6f", x"70", x"6f", x"6f", x"6f", x"6e", x"6c", x"6d", 
        x"6c", x"6d", x"6d", x"6c", x"6e", x"6b", x"6e", x"6f", x"6f", x"6f", x"6e", x"6d", x"6c", x"6c", x"6d", 
        x"6d", x"6d", x"6d", x"6e", x"6f", x"6f", x"6f", x"6f", x"6c", x"6c", x"6e", x"6c", x"6b", x"6a", x"6c", 
        x"72", x"6e", x"6e", x"6e", x"6c", x"6e", x"6a", x"6a", x"6c", x"6d", x"6a", x"68", x"69", x"6c", x"6c", 
        x"6b", x"6d", x"6d", x"6d", x"6d", x"6e", x"6d", x"6b", x"6c", x"6c", x"6e", x"6d", x"6b", x"6b", x"6a", 
        x"6b", x"6b", x"6a", x"6a", x"6c", x"6c", x"6a", x"6d", x"6f", x"6d", x"6d", x"6e", x"6d", x"6c", x"6e", 
        x"6e", x"6c", x"6a", x"6a", x"69", x"6b", x"6d", x"6d", x"6e", x"6f", x"6e", x"6d", x"6d", x"6e", x"6d", 
        x"6d", x"6c", x"6c", x"6e", x"6e", x"6c", x"6c", x"6e", x"6d", x"6a", x"6a", x"6d", x"6f", x"6c", x"6c", 
        x"6d", x"6d", x"6e", x"70", x"71", x"6e", x"6c", x"6d", x"6e", x"6e", x"6f", x"6e", x"6f", x"70", x"6f", 
        x"6c", x"6c", x"6b", x"6d", x"6f", x"6e", x"6f", x"6f", x"70", x"6f", x"6f", x"6f", x"70", x"71", x"72", 
        x"6e", x"6d", x"6f", x"71", x"6f", x"70", x"70", x"70", x"71", x"70", x"6e", x"6e", x"73", x"73", x"72", 
        x"72", x"6f", x"70", x"72", x"72", x"72", x"71", x"71", x"73", x"72", x"72", x"74", x"74", x"72", x"71", 
        x"72", x"72", x"71", x"72", x"73", x"74", x"73", x"74", x"73", x"72", x"71", x"6f", x"72", x"74", x"6b", 
        x"8d", x"d7", x"d2", x"ce", x"cf", x"d0", x"d8", x"d2", x"cc", x"ce", x"cf", x"cf", x"ce", x"ce", x"cf", 
        x"ce", x"cd", x"cc", x"cd", x"ce", x"cf", x"cf", x"cf", x"ce", x"ce", x"ce", x"d0", x"cf", x"ce", x"cd", 
        x"ce", x"ce", x"ce", x"cf", x"cf", x"d0", x"d0", x"ce", x"cf", x"cf", x"d0", x"cf", x"cd", x"cd", x"ce", 
        x"cf", x"cf", x"cf", x"ce", x"ce", x"ce", x"cf", x"d7", x"cb", x"d3", x"d3", x"d1", x"d2", x"d1", x"c0", 
        x"86", x"5f", x"5b", x"5e", x"5e", x"5c", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"5c", x"5f", 
        x"60", x"5e", x"60", x"5d", x"6d", x"9e", x"d4", x"f0", x"f5", x"f7", x"f7", x"fa", x"fc", x"fb", x"fb", 
        x"fa", x"fb", x"fc", x"fb", x"fa", x"fa", x"f9", x"f7", x"fa", x"fc", x"fb", x"f9", x"f0", x"da", x"b3", 
        x"94", x"87", x"89", x"87", x"82", x"7b", x"7e", x"8b", x"99", x"a0", x"bc", x"c8", x"c7", x"c3", x"c5", 
        x"c0", x"88", x"61", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"b4", x"ea", 
        x"ed", x"ed", x"ed", x"ec", x"ed", x"ed", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ee", x"f0", x"ee", x"eb", x"ec", x"ee", x"ee", x"ee", x"ea", x"e3", x"d9", x"ce", x"cb", 
        x"d5", x"df", x"d1", x"b4", x"8c", x"71", x"6e", x"78", x"7b", x"7b", x"7b", x"7a", x"7b", x"7a", x"7a", 
        x"7b", x"7b", x"79", x"7a", x"7c", x"7d", x"7c", x"7b", x"7a", x"79", x"79", x"7a", x"7b", x"7a", x"7a", 
        x"79", x"79", x"78", x"79", x"79", x"79", x"79", x"79", x"7a", x"7c", x"7a", x"7b", x"7b", x"7a", x"79", 
        x"78", x"79", x"7a", x"79", x"77", x"78", x"79", x"7a", x"7a", x"7a", x"79", x"78", x"79", x"79", x"79", 
        x"7a", x"78", x"76", x"79", x"79", x"78", x"78", x"78", x"77", x"77", x"78", x"78", x"76", x"78", x"78", 
        x"77", x"77", x"76", x"75", x"76", x"78", x"79", x"78", x"77", x"78", x"7a", x"79", x"78", x"78", x"79", 
        x"79", x"77", x"76", x"78", x"79", x"77", x"77", x"78", x"79", x"77", x"75", x"76", x"77", x"78", x"78", 
        x"77", x"77", x"76", x"76", x"76", x"74", x"75", x"74", x"75", x"77", x"76", x"74", x"75", x"77", x"77", 
        x"78", x"78", x"75", x"75", x"77", x"77", x"74", x"73", x"77", x"77", x"76", x"75", x"76", x"78", x"78", 
        x"77", x"77", x"75", x"73", x"73", x"75", x"75", x"76", x"75", x"75", x"75", x"75", x"74", x"74", x"75", 
        x"76", x"75", x"77", x"77", x"76", x"75", x"72", x"74", x"76", x"74", x"74", x"74", x"75", x"75", x"75", 
        x"72", x"75", x"73", x"73", x"76", x"75", x"75", x"75", x"75", x"75", x"74", x"73", x"74", x"77", x"76", 
        x"74", x"75", x"75", x"76", x"77", x"76", x"75", x"73", x"74", x"76", x"75", x"74", x"76", x"75", x"76", 
        x"75", x"73", x"76", x"76", x"73", x"75", x"73", x"74", x"75", x"74", x"73", x"74", x"74", x"74", x"74", 
        x"75", x"75", x"75", x"74", x"74", x"75", x"74", x"74", x"73", x"72", x"71", x"71", x"72", x"73", x"76", 
        x"77", x"74", x"75", x"75", x"74", x"75", x"75", x"74", x"72", x"73", x"75", x"76", x"72", x"72", x"72", 
        x"73", x"74", x"72", x"71", x"72", x"73", x"73", x"72", x"72", x"72", x"71", x"6f", x"6f", x"70", x"71", 
        x"73", x"74", x"74", x"73", x"71", x"70", x"70", x"71", x"71", x"6f", x"6e", x"6f", x"71", x"6e", x"6d", 
        x"71", x"72", x"70", x"70", x"71", x"70", x"6f", x"6e", x"6f", x"70", x"6f", x"6d", x"6f", x"70", x"70", 
        x"72", x"71", x"71", x"70", x"6e", x"70", x"71", x"70", x"70", x"6f", x"70", x"70", x"70", x"70", x"70", 
        x"71", x"71", x"6f", x"6b", x"6b", x"70", x"71", x"6f", x"6c", x"6c", x"6f", x"70", x"6f", x"6f", x"6d", 
        x"6d", x"70", x"6f", x"70", x"70", x"71", x"6f", x"6f", x"71", x"6f", x"6d", x"6f", x"6f", x"6f", x"6e", 
        x"6f", x"6f", x"6f", x"6f", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6f", x"70", x"72", 
        x"72", x"70", x"6f", x"6f", x"70", x"6f", x"6f", x"6e", x"6f", x"70", x"6f", x"6c", x"6c", x"6c", x"6c", 
        x"6d", x"6d", x"6d", x"6e", x"6e", x"6f", x"6e", x"6e", x"6b", x"6b", x"6e", x"6c", x"6c", x"6b", x"6d", 
        x"6e", x"6c", x"6c", x"6c", x"6b", x"6b", x"68", x"69", x"6c", x"6d", x"6b", x"69", x"6a", x"6e", x"6b", 
        x"6a", x"6d", x"6d", x"6b", x"6a", x"6b", x"6d", x"6e", x"6d", x"6d", x"6c", x"6c", x"6d", x"6c", x"6a", 
        x"6b", x"6b", x"69", x"6a", x"6c", x"6e", x"6e", x"6e", x"6d", x"6c", x"6e", x"6e", x"6b", x"68", x"6a", 
        x"6c", x"6c", x"6b", x"6a", x"6a", x"6a", x"6b", x"6d", x"6e", x"6e", x"6c", x"6b", x"6c", x"70", x"70", 
        x"6f", x"6d", x"6c", x"6c", x"6e", x"6f", x"6f", x"70", x"6e", x"6c", x"6c", x"6f", x"6f", x"6c", x"6d", 
        x"6d", x"6c", x"6d", x"6f", x"70", x"6d", x"6e", x"70", x"6f", x"6e", x"6e", x"6d", x"6d", x"6d", x"6d", 
        x"6b", x"6b", x"6c", x"6f", x"6f", x"6e", x"6f", x"70", x"71", x"70", x"6d", x"6b", x"6b", x"6e", x"70", 
        x"6e", x"6d", x"6e", x"6e", x"6f", x"70", x"71", x"71", x"72", x"72", x"73", x"72", x"75", x"74", x"73", 
        x"74", x"71", x"71", x"72", x"73", x"72", x"71", x"72", x"74", x"70", x"71", x"74", x"72", x"70", x"6f", 
        x"71", x"72", x"71", x"72", x"72", x"72", x"72", x"72", x"72", x"73", x"72", x"72", x"75", x"77", x"6d", 
        x"90", x"d8", x"d3", x"ce", x"d0", x"d2", x"d9", x"d2", x"cd", x"ce", x"d0", x"cf", x"ce", x"ce", x"cf", 
        x"ce", x"cd", x"cc", x"cc", x"ce", x"cf", x"cf", x"cf", x"d0", x"cf", x"cf", x"d1", x"d1", x"cf", x"ce", 
        x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"d0", x"ce", x"cf", x"cf", x"d0", x"cf", x"cd", x"cd", x"ce", 
        x"cf", x"cf", x"cf", x"ce", x"ce", x"cd", x"cb", x"db", x"cd", x"d3", x"d5", x"d2", x"d0", x"d1", x"c4", 
        x"88", x"5b", x"5b", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"61", x"5d", 
        x"5e", x"61", x"5f", x"5f", x"5a", x"63", x"83", x"ba", x"e4", x"f5", x"fa", x"fb", x"fd", x"fb", x"fc", 
        x"fb", x"fa", x"fc", x"fc", x"fd", x"f9", x"f8", x"fb", x"fb", x"f9", x"f9", x"f7", x"f8", x"f8", x"f2", 
        x"e7", x"e1", x"e3", x"e2", x"dc", x"d8", x"da", x"e2", x"ea", x"ee", x"f5", x"f8", x"f8", x"f5", x"f1", 
        x"e1", x"99", x"65", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5d", x"5e", x"ad", x"e9", 
        x"ed", x"ed", x"ec", x"ed", x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ed", x"ee", x"ee", x"ed", x"ee", x"f0", x"ed", x"e7", x"de", 
        x"cf", x"c2", x"d3", x"e5", x"de", x"b8", x"8f", x"6b", x"6c", x"75", x"7b", x"7c", x"79", x"78", x"78", 
        x"78", x"79", x"7b", x"7b", x"7a", x"78", x"7b", x"7b", x"7a", x"79", x"79", x"7a", x"7b", x"7b", x"7b", 
        x"7a", x"7a", x"7a", x"7b", x"7b", x"7b", x"7c", x"7b", x"7b", x"7b", x"78", x"78", x"77", x"7a", x"79", 
        x"79", x"7a", x"7a", x"78", x"77", x"78", x"79", x"79", x"78", x"78", x"77", x"77", x"7a", x"7a", x"79", 
        x"78", x"78", x"78", x"7d", x"7a", x"77", x"78", x"79", x"78", x"77", x"78", x"78", x"78", x"7a", x"7b", 
        x"7a", x"79", x"79", x"78", x"75", x"77", x"77", x"76", x"75", x"76", x"77", x"79", x"78", x"77", x"78", 
        x"79", x"78", x"76", x"77", x"79", x"78", x"75", x"75", x"77", x"77", x"75", x"75", x"76", x"78", x"79", 
        x"78", x"77", x"76", x"77", x"76", x"75", x"72", x"72", x"75", x"76", x"75", x"73", x"75", x"76", x"75", 
        x"76", x"77", x"75", x"73", x"77", x"78", x"76", x"74", x"75", x"79", x"77", x"76", x"76", x"78", x"78", 
        x"78", x"78", x"77", x"75", x"75", x"77", x"78", x"77", x"75", x"74", x"75", x"75", x"72", x"72", x"74", 
        x"75", x"73", x"75", x"76", x"76", x"77", x"75", x"75", x"73", x"73", x"72", x"72", x"72", x"72", x"74", 
        x"73", x"77", x"76", x"75", x"76", x"75", x"74", x"75", x"75", x"75", x"74", x"73", x"75", x"79", x"76", 
        x"73", x"73", x"73", x"74", x"76", x"76", x"75", x"75", x"77", x"78", x"77", x"77", x"77", x"77", x"76", 
        x"74", x"72", x"77", x"76", x"73", x"77", x"78", x"75", x"74", x"75", x"75", x"72", x"70", x"73", x"75", 
        x"76", x"76", x"76", x"75", x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"72", x"74", 
        x"77", x"73", x"74", x"76", x"73", x"73", x"75", x"76", x"75", x"75", x"75", x"74", x"72", x"72", x"72", 
        x"73", x"74", x"72", x"71", x"71", x"72", x"72", x"72", x"72", x"72", x"72", x"71", x"72", x"72", x"72", 
        x"72", x"71", x"71", x"74", x"74", x"72", x"71", x"71", x"70", x"6e", x"6d", x"6f", x"72", x"6f", x"6f", 
        x"73", x"72", x"6f", x"70", x"71", x"70", x"6f", x"6e", x"70", x"70", x"6c", x"6b", x"71", x"73", x"72", 
        x"73", x"71", x"72", x"72", x"71", x"71", x"71", x"71", x"70", x"6d", x"6e", x"70", x"6f", x"6f", x"6f", 
        x"71", x"73", x"72", x"6e", x"6e", x"70", x"70", x"6e", x"6b", x"6e", x"6f", x"70", x"6f", x"6d", x"6e", 
        x"6e", x"6c", x"6c", x"6e", x"6d", x"6e", x"6c", x"6d", x"6d", x"6e", x"6e", x"6f", x"71", x"71", x"70", 
        x"6f", x"6e", x"6e", x"6f", x"6f", x"6f", x"6f", x"71", x"71", x"70", x"6e", x"6b", x"6b", x"6d", x"72", 
        x"74", x"71", x"6f", x"6f", x"6f", x"6f", x"6d", x"6c", x"6d", x"6f", x"6f", x"6e", x"6e", x"6e", x"6c", 
        x"6c", x"6d", x"6d", x"6e", x"6e", x"6e", x"6e", x"6f", x"6c", x"6c", x"6f", x"6c", x"6b", x"6b", x"6c", 
        x"71", x"6f", x"70", x"6f", x"70", x"6e", x"6b", x"6a", x"6b", x"6d", x"6c", x"6a", x"6a", x"6d", x"6f", 
        x"6e", x"6e", x"6d", x"6c", x"6c", x"6d", x"6c", x"6a", x"6a", x"6c", x"6a", x"6b", x"6c", x"6d", x"70", 
        x"6f", x"6e", x"6d", x"6d", x"6e", x"70", x"6f", x"6d", x"6b", x"6c", x"6f", x"6f", x"6b", x"69", x"68", 
        x"69", x"6c", x"6b", x"69", x"6a", x"6a", x"6a", x"6d", x"6e", x"6d", x"6b", x"6a", x"6b", x"6e", x"71", 
        x"70", x"6e", x"6e", x"6f", x"70", x"6f", x"6e", x"6d", x"6c", x"6d", x"6b", x"6f", x"6e", x"6e", x"6e", 
        x"6e", x"6b", x"6c", x"6f", x"6d", x"6b", x"6e", x"71", x"6f", x"6d", x"6d", x"6f", x"6f", x"6e", x"6e", 
        x"6d", x"6c", x"6f", x"70", x"6f", x"6e", x"6f", x"70", x"71", x"70", x"6f", x"6e", x"6e", x"70", x"71", 
        x"71", x"72", x"73", x"70", x"72", x"72", x"72", x"71", x"6f", x"71", x"74", x"73", x"75", x"73", x"71", 
        x"72", x"71", x"6f", x"71", x"73", x"74", x"74", x"74", x"75", x"6f", x"6f", x"73", x"72", x"71", x"72", 
        x"74", x"73", x"72", x"73", x"71", x"71", x"72", x"71", x"71", x"73", x"72", x"73", x"77", x"77", x"6c", 
        x"91", x"d8", x"d3", x"ce", x"d1", x"d3", x"d9", x"d2", x"cd", x"ce", x"d0", x"cf", x"cf", x"cf", x"cf", 
        x"cf", x"ce", x"cd", x"ce", x"d0", x"d0", x"cf", x"d0", x"d1", x"cf", x"ce", x"d2", x"d0", x"ce", x"cf", 
        x"d0", x"cf", x"cf", x"d0", x"d0", x"d0", x"cf", x"ce", x"cf", x"cf", x"d0", x"cf", x"ce", x"cd", x"ce", 
        x"cf", x"cf", x"cf", x"ce", x"ce", x"cd", x"cc", x"db", x"ce", x"d3", x"d1", x"d0", x"d4", x"d6", x"b7", 
        x"7b", x"61", x"60", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"60", x"61", 
        x"5d", x"5c", x"5f", x"5e", x"5d", x"5e", x"60", x"69", x"8a", x"b2", x"db", x"eb", x"f7", x"fb", x"fc", 
        x"fb", x"f9", x"fb", x"fa", x"fb", x"fc", x"fb", x"fc", x"fd", x"fb", x"fa", x"fb", x"fa", x"fa", x"fb", 
        x"fa", x"f9", x"f9", x"f9", x"f9", x"f9", x"f9", x"fa", x"f9", x"fa", x"f7", x"f5", x"ed", x"e2", x"ce", 
        x"a7", x"72", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"a7", x"e9", 
        x"ed", x"ed", x"ec", x"ed", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ed", x"ee", x"ed", x"ec", x"ee", x"ef", x"ef", x"ed", x"ed", x"ec", x"ec", x"ee", x"ef", x"ee", x"ec", 
        x"ea", x"e4", x"d3", x"ca", x"d6", x"e1", x"df", x"cd", x"a4", x"7d", x"6b", x"72", x"79", x"7a", x"7e", 
        x"7e", x"7d", x"7d", x"7b", x"7a", x"79", x"7a", x"7b", x"7a", x"7a", x"7a", x"7b", x"7c", x"7b", x"7b", 
        x"7a", x"7a", x"7a", x"7b", x"7a", x"79", x"79", x"7a", x"7a", x"7b", x"7a", x"7b", x"79", x"7a", x"7a", 
        x"7a", x"7b", x"7a", x"78", x"77", x"7a", x"7a", x"7a", x"79", x"79", x"78", x"78", x"79", x"78", x"79", 
        x"7b", x"7a", x"79", x"7c", x"76", x"71", x"74", x"78", x"79", x"7a", x"7a", x"79", x"76", x"77", x"7a", 
        x"79", x"76", x"76", x"78", x"77", x"77", x"77", x"77", x"78", x"78", x"78", x"7b", x"78", x"76", x"76", 
        x"77", x"79", x"78", x"77", x"7a", x"7a", x"76", x"76", x"76", x"77", x"79", x"77", x"77", x"76", x"76", 
        x"76", x"76", x"77", x"78", x"79", x"79", x"76", x"75", x"77", x"76", x"76", x"77", x"77", x"76", x"74", 
        x"73", x"75", x"77", x"74", x"77", x"77", x"76", x"73", x"70", x"71", x"74", x"76", x"78", x"79", x"78", 
        x"76", x"75", x"75", x"76", x"78", x"78", x"76", x"74", x"75", x"76", x"73", x"72", x"74", x"75", x"75", 
        x"77", x"77", x"77", x"76", x"73", x"74", x"72", x"73", x"73", x"75", x"74", x"75", x"75", x"74", x"76", 
        x"74", x"77", x"76", x"75", x"77", x"74", x"72", x"74", x"75", x"75", x"75", x"76", x"76", x"76", x"76", 
        x"76", x"75", x"75", x"75", x"75", x"74", x"74", x"74", x"77", x"77", x"75", x"75", x"74", x"77", x"77", 
        x"75", x"74", x"76", x"76", x"75", x"78", x"77", x"74", x"74", x"76", x"77", x"74", x"71", x"74", x"76", 
        x"76", x"76", x"76", x"76", x"75", x"74", x"74", x"74", x"73", x"73", x"74", x"73", x"72", x"70", x"72", 
        x"74", x"71", x"73", x"75", x"74", x"74", x"75", x"74", x"75", x"76", x"75", x"74", x"73", x"72", x"72", 
        x"72", x"73", x"72", x"72", x"73", x"73", x"74", x"73", x"74", x"73", x"73", x"71", x"72", x"73", x"72", 
        x"70", x"70", x"70", x"71", x"72", x"71", x"71", x"72", x"71", x"71", x"6f", x"6f", x"72", x"70", x"70", 
        x"72", x"71", x"6f", x"70", x"70", x"71", x"70", x"70", x"70", x"70", x"6e", x"70", x"73", x"73", x"71", 
        x"70", x"6e", x"70", x"70", x"70", x"6e", x"6c", x"6e", x"6d", x"6c", x"6e", x"70", x"70", x"6f", x"6f", 
        x"70", x"73", x"72", x"6f", x"70", x"71", x"70", x"6f", x"6d", x"6f", x"6f", x"6e", x"6e", x"6d", x"70", 
        x"71", x"6f", x"6f", x"6f", x"6c", x"6c", x"6b", x"6e", x"6f", x"70", x"70", x"6f", x"70", x"71", x"6f", 
        x"6e", x"6d", x"6e", x"6f", x"6f", x"6e", x"70", x"6f", x"6d", x"6d", x"6d", x"6c", x"6d", x"70", x"72", 
        x"73", x"71", x"70", x"70", x"6e", x"70", x"6e", x"6c", x"6d", x"6f", x"6f", x"70", x"70", x"71", x"6e", 
        x"6e", x"6d", x"6e", x"6e", x"6f", x"6f", x"70", x"71", x"70", x"6e", x"6e", x"6a", x"6a", x"6e", x"6f", 
        x"71", x"6e", x"6f", x"6d", x"6e", x"6c", x"6a", x"6c", x"6d", x"6d", x"6c", x"6a", x"6a", x"6b", x"6d", 
        x"6e", x"6d", x"6d", x"6d", x"6d", x"6c", x"6c", x"6b", x"6d", x"70", x"6d", x"6d", x"6e", x"6c", x"6f", 
        x"6e", x"6d", x"6d", x"6e", x"6e", x"6f", x"6c", x"6b", x"6c", x"6e", x"6e", x"6e", x"6e", x"70", x"6d", 
        x"6c", x"6d", x"6d", x"6c", x"6d", x"6c", x"6c", x"6d", x"6d", x"6c", x"6c", x"6d", x"6c", x"6e", x"71", 
        x"6f", x"6d", x"6f", x"72", x"72", x"6f", x"6f", x"71", x"71", x"72", x"6d", x"6e", x"6d", x"6e", x"71", 
        x"6f", x"6b", x"6b", x"6e", x"6d", x"6e", x"71", x"72", x"70", x"6e", x"6f", x"72", x"71", x"70", x"70", 
        x"6e", x"6c", x"6f", x"70", x"6f", x"6f", x"6f", x"70", x"71", x"70", x"70", x"6f", x"6e", x"6f", x"6e", 
        x"6d", x"70", x"71", x"6f", x"72", x"70", x"72", x"72", x"71", x"74", x"73", x"73", x"75", x"73", x"71", 
        x"73", x"74", x"72", x"72", x"73", x"73", x"73", x"74", x"76", x"6f", x"6e", x"71", x"70", x"70", x"72", 
        x"72", x"72", x"73", x"73", x"71", x"72", x"74", x"74", x"73", x"74", x"75", x"76", x"78", x"75", x"69", 
        x"8e", x"d8", x"d2", x"ce", x"d2", x"d4", x"d9", x"d1", x"cd", x"ce", x"d0", x"d0", x"cf", x"cf", x"cf", 
        x"cf", x"cf", x"cd", x"ce", x"cf", x"d0", x"cf", x"cf", x"d0", x"cd", x"cc", x"d1", x"cf", x"cc", x"cf", 
        x"d0", x"cf", x"cf", x"d0", x"d1", x"cf", x"cd", x"cd", x"ce", x"ce", x"d0", x"cf", x"ce", x"ce", x"ce", 
        x"cf", x"cf", x"cf", x"ce", x"ce", x"ce", x"ce", x"d9", x"cf", x"d1", x"cd", x"d4", x"ce", x"aa", x"95", 
        x"71", x"5f", x"61", x"60", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5b", x"61", 
        x"5f", x"5b", x"62", x"5e", x"5c", x"60", x"60", x"5d", x"5a", x"63", x"81", x"b4", x"e9", x"fa", x"f9", 
        x"fa", x"fa", x"fb", x"fb", x"f9", x"fb", x"fc", x"fa", x"fb", x"fb", x"f9", x"f9", x"fb", x"fc", x"fb", 
        x"f9", x"f9", x"fb", x"fc", x"fb", x"f9", x"f9", x"fb", x"f8", x"ee", x"e0", x"c9", x"a8", x"89", x"73", 
        x"61", x"5c", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"a3", x"e9", 
        x"ed", x"ed", x"ec", x"ed", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ed", x"ee", x"ed", x"ec", x"ec", x"ed", x"ed", x"ed", x"ee", x"ed", x"ec", x"ed", x"ee", x"ef", x"ef", 
        x"ee", x"ef", x"ed", x"e7", x"d6", x"c7", x"cd", x"dc", x"e3", x"d6", x"b2", x"83", x"6f", x"6e", x"74", 
        x"7b", x"7f", x"7d", x"7a", x"7c", x"7e", x"7d", x"7c", x"7b", x"7a", x"79", x"7a", x"7b", x"7b", x"7b", 
        x"7a", x"7a", x"7b", x"7c", x"7b", x"7a", x"7b", x"7c", x"7b", x"7b", x"7b", x"7c", x"79", x"79", x"79", 
        x"7a", x"7b", x"7b", x"79", x"77", x"7a", x"7b", x"7b", x"7b", x"7a", x"79", x"78", x"79", x"78", x"78", 
        x"7a", x"7a", x"78", x"78", x"78", x"78", x"79", x"7a", x"7a", x"7a", x"79", x"79", x"79", x"7a", x"7e", 
        x"7c", x"78", x"79", x"7b", x"78", x"76", x"76", x"79", x"7b", x"7b", x"79", x"7a", x"79", x"79", x"79", 
        x"7a", x"79", x"78", x"77", x"7a", x"7b", x"78", x"7b", x"78", x"76", x"76", x"75", x"76", x"77", x"78", 
        x"78", x"79", x"79", x"77", x"77", x"79", x"77", x"77", x"7a", x"77", x"77", x"79", x"79", x"77", x"76", 
        x"76", x"77", x"78", x"77", x"77", x"76", x"75", x"75", x"72", x"77", x"79", x"78", x"77", x"77", x"77", 
        x"78", x"77", x"78", x"78", x"78", x"77", x"77", x"77", x"78", x"78", x"75", x"74", x"76", x"77", x"77", 
        x"77", x"75", x"76", x"75", x"74", x"75", x"73", x"74", x"72", x"74", x"72", x"75", x"76", x"73", x"75", 
        x"76", x"78", x"75", x"75", x"79", x"77", x"75", x"76", x"75", x"74", x"75", x"76", x"77", x"74", x"76", 
        x"78", x"76", x"76", x"76", x"75", x"75", x"75", x"75", x"78", x"77", x"73", x"73", x"73", x"77", x"78", 
        x"78", x"77", x"74", x"75", x"77", x"75", x"73", x"72", x"72", x"74", x"75", x"76", x"75", x"76", x"76", 
        x"75", x"74", x"75", x"75", x"76", x"74", x"76", x"75", x"73", x"73", x"75", x"74", x"73", x"72", x"71", 
        x"72", x"72", x"75", x"76", x"77", x"76", x"74", x"72", x"74", x"76", x"76", x"75", x"74", x"73", x"72", 
        x"72", x"73", x"72", x"72", x"74", x"74", x"73", x"73", x"73", x"72", x"72", x"6f", x"6f", x"72", x"72", 
        x"70", x"6f", x"70", x"6f", x"6f", x"71", x"72", x"71", x"72", x"73", x"72", x"71", x"72", x"71", x"70", 
        x"71", x"70", x"6f", x"6f", x"70", x"71", x"71", x"72", x"70", x"6f", x"6d", x"70", x"70", x"71", x"71", 
        x"71", x"73", x"73", x"71", x"71", x"6e", x"6d", x"71", x"70", x"6c", x"6c", x"6d", x"6d", x"6d", x"6c", 
        x"6c", x"6f", x"6d", x"6b", x"6f", x"6e", x"6e", x"6f", x"6d", x"6f", x"6e", x"6d", x"6e", x"6d", x"71", 
        x"71", x"70", x"72", x"73", x"6d", x"6b", x"6b", x"6f", x"71", x"72", x"70", x"6e", x"6e", x"70", x"70", 
        x"6f", x"6e", x"6f", x"70", x"6e", x"6c", x"6f", x"6f", x"6e", x"6f", x"70", x"6f", x"6f", x"6f", x"6e", 
        x"6e", x"6d", x"6f", x"71", x"6f", x"74", x"72", x"70", x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"6d", 
        x"6c", x"6c", x"6c", x"6c", x"6d", x"6e", x"6e", x"71", x"6f", x"6d", x"6d", x"6c", x"6e", x"6f", x"6d", 
        x"72", x"71", x"71", x"6e", x"6f", x"6e", x"6d", x"6f", x"6e", x"6c", x"6b", x"6b", x"6b", x"6a", x"6b", 
        x"6d", x"6e", x"6f", x"6f", x"6e", x"6b", x"6b", x"6c", x"6c", x"6c", x"6a", x"6b", x"6c", x"6b", x"6a", 
        x"6a", x"6b", x"6c", x"6d", x"6d", x"6e", x"6c", x"6c", x"6e", x"6d", x"6b", x"6b", x"6d", x"71", x"6e", 
        x"6a", x"6b", x"6c", x"6e", x"6f", x"6d", x"6c", x"6e", x"6d", x"6b", x"6c", x"6f", x"6d", x"6e", x"70", 
        x"6f", x"6d", x"6f", x"70", x"6f", x"6b", x"6d", x"71", x"71", x"70", x"6b", x"6c", x"6e", x"6f", x"71", 
        x"6f", x"6b", x"6b", x"6f", x"6b", x"6c", x"70", x"70", x"6e", x"6d", x"6d", x"6f", x"6f", x"6f", x"70", 
        x"6e", x"6e", x"70", x"70", x"6f", x"6f", x"70", x"71", x"71", x"71", x"70", x"71", x"72", x"72", x"70", 
        x"6e", x"6f", x"71", x"72", x"74", x"71", x"71", x"71", x"70", x"72", x"70", x"70", x"72", x"71", x"6f", 
        x"71", x"73", x"74", x"74", x"73", x"71", x"71", x"72", x"75", x"72", x"72", x"75", x"73", x"72", x"72", 
        x"73", x"72", x"73", x"74", x"73", x"73", x"75", x"74", x"74", x"77", x"77", x"78", x"79", x"75", x"6b", 
        x"8e", x"d8", x"d2", x"cf", x"d1", x"d4", x"d9", x"d0", x"cd", x"ce", x"d0", x"d0", x"cf", x"cf", x"d0", 
        x"cf", x"ce", x"cd", x"cd", x"ce", x"cf", x"ce", x"ce", x"cf", x"cd", x"cc", x"cf", x"cd", x"cc", x"cf", 
        x"d1", x"cf", x"cf", x"d0", x"d1", x"cf", x"ce", x"cd", x"cd", x"cf", x"d0", x"d0", x"cf", x"cf", x"ce", 
        x"cd", x"ce", x"cf", x"cd", x"cf", x"cf", x"ce", x"d7", x"cc", x"d3", x"d7", x"bf", x"a1", x"a1", x"b8", 
        x"92", x"62", x"5e", x"5e", x"5c", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5c", x"5c", 
        x"5f", x"5d", x"5d", x"5e", x"5f", x"60", x"5c", x"60", x"5e", x"5b", x"70", x"ae", x"e8", x"f9", x"f5", 
        x"f7", x"f5", x"e9", x"e6", x"ea", x"ed", x"f4", x"f9", x"f9", x"f8", x"f8", x"f7", x"f1", x"ea", x"e3", 
        x"e2", x"ed", x"f0", x"f0", x"ef", x"ea", x"e4", x"da", x"c6", x"a9", x"8a", x"71", x"63", x"5c", x"5d", 
        x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"a1", x"e9", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ed", 
        x"ed", x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ed", x"ec", x"ed", x"ed", x"ec", x"ec", x"ec", 
        x"ee", x"ee", x"ee", x"ec", x"ee", x"ea", x"db", x"cb", x"cf", x"d7", x"df", x"da", x"b9", x"90", x"77", 
        x"70", x"72", x"78", x"7c", x"7d", x"7b", x"7d", x"7e", x"7d", x"7a", x"79", x"7a", x"79", x"7a", x"7d", 
        x"7d", x"7c", x"7d", x"7e", x"7d", x"7b", x"7a", x"7b", x"7b", x"7c", x"7d", x"7f", x"7b", x"79", x"79", 
        x"79", x"7a", x"7b", x"79", x"78", x"7a", x"7b", x"7b", x"7b", x"7a", x"7a", x"79", x"7a", x"7a", x"78", 
        x"78", x"78", x"77", x"76", x"79", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", x"79", x"78", x"79", x"7c", 
        x"7a", x"77", x"78", x"79", x"77", x"76", x"76", x"78", x"7a", x"7a", x"79", x"78", x"79", x"7c", x"7b", 
        x"7a", x"7a", x"77", x"76", x"77", x"78", x"77", x"7b", x"77", x"73", x"75", x"76", x"78", x"7a", x"7a", 
        x"79", x"77", x"78", x"76", x"75", x"77", x"76", x"78", x"7b", x"78", x"76", x"79", x"79", x"78", x"78", 
        x"79", x"78", x"78", x"77", x"77", x"76", x"76", x"78", x"75", x"74", x"76", x"78", x"78", x"77", x"77", 
        x"77", x"77", x"76", x"74", x"73", x"72", x"73", x"76", x"79", x"79", x"78", x"77", x"76", x"77", x"78", 
        x"78", x"75", x"74", x"76", x"77", x"76", x"73", x"73", x"74", x"74", x"73", x"76", x"76", x"73", x"75", 
        x"77", x"78", x"74", x"75", x"79", x"79", x"77", x"78", x"75", x"74", x"75", x"76", x"76", x"75", x"73", 
        x"74", x"74", x"73", x"73", x"74", x"74", x"75", x"77", x"79", x"77", x"75", x"75", x"74", x"78", x"77", 
        x"78", x"78", x"74", x"75", x"77", x"76", x"74", x"74", x"74", x"73", x"74", x"76", x"77", x"76", x"75", 
        x"74", x"75", x"75", x"76", x"77", x"75", x"75", x"75", x"74", x"75", x"77", x"76", x"76", x"75", x"74", 
        x"73", x"74", x"76", x"77", x"76", x"76", x"75", x"74", x"76", x"78", x"75", x"73", x"74", x"73", x"72", 
        x"72", x"73", x"73", x"72", x"72", x"72", x"73", x"73", x"73", x"72", x"71", x"70", x"72", x"73", x"71", 
        x"6f", x"6e", x"6e", x"6e", x"70", x"72", x"72", x"72", x"73", x"72", x"72", x"72", x"71", x"71", x"70", 
        x"6f", x"71", x"72", x"71", x"70", x"71", x"71", x"72", x"70", x"70", x"71", x"72", x"70", x"6e", x"6f", 
        x"6f", x"72", x"71", x"71", x"72", x"70", x"6e", x"72", x"72", x"6e", x"6f", x"6f", x"6f", x"6f", x"6f", 
        x"6e", x"70", x"6f", x"6e", x"72", x"72", x"72", x"71", x"6f", x"70", x"70", x"6e", x"70", x"70", x"72", 
        x"71", x"6d", x"70", x"71", x"6d", x"6e", x"6d", x"6f", x"70", x"70", x"6f", x"6e", x"6e", x"70", x"71", 
        x"71", x"71", x"70", x"70", x"6f", x"6d", x"6f", x"6e", x"6c", x"6e", x"71", x"72", x"71", x"71", x"70", 
        x"6e", x"70", x"70", x"6e", x"6a", x"6e", x"6e", x"72", x"71", x"6f", x"6e", x"6f", x"6e", x"6e", x"6e", 
        x"6d", x"6e", x"6c", x"6d", x"6f", x"71", x"6e", x"70", x"6e", x"6e", x"6f", x"70", x"72", x"70", x"6d", 
        x"6f", x"71", x"72", x"70", x"6b", x"6e", x"6d", x"6f", x"6f", x"6b", x"6a", x"6b", x"6c", x"6c", x"6d", 
        x"6d", x"6e", x"6e", x"6d", x"6b", x"68", x"68", x"6b", x"6c", x"6c", x"6d", x"6e", x"6e", x"6d", x"6a", 
        x"6c", x"6f", x"6f", x"6c", x"6a", x"6d", x"6c", x"6c", x"6d", x"6b", x"6a", x"6d", x"6e", x"70", x"71", 
        x"6e", x"6b", x"6d", x"70", x"6c", x"6a", x"6a", x"6e", x"6f", x"6b", x"6e", x"70", x"6d", x"6d", x"6f", 
        x"71", x"70", x"6f", x"6e", x"6e", x"6e", x"70", x"71", x"70", x"6e", x"6f", x"71", x"72", x"6f", x"6f", 
        x"70", x"6e", x"6e", x"70", x"6c", x"6b", x"6f", x"6f", x"6c", x"6e", x"6d", x"6f", x"70", x"71", x"71", 
        x"70", x"70", x"6e", x"6f", x"70", x"70", x"72", x"72", x"71", x"71", x"70", x"70", x"71", x"71", x"70", 
        x"70", x"71", x"72", x"72", x"72", x"72", x"73", x"73", x"72", x"72", x"75", x"73", x"72", x"72", x"70", 
        x"71", x"74", x"72", x"72", x"73", x"72", x"72", x"72", x"74", x"73", x"73", x"77", x"74", x"74", x"71", 
        x"74", x"74", x"74", x"75", x"75", x"74", x"74", x"73", x"73", x"74", x"75", x"74", x"77", x"77", x"6e", 
        x"8c", x"d6", x"d1", x"d1", x"d0", x"d3", x"dc", x"d1", x"cc", x"ce", x"cf", x"cf", x"cf", x"cf", x"d0", 
        x"d0", x"cf", x"ce", x"ce", x"cf", x"d0", x"cf", x"d0", x"d0", x"d0", x"cf", x"cd", x"cd", x"ce", x"d0", 
        x"d0", x"d1", x"d1", x"d1", x"d0", x"d0", x"cf", x"cf", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"ce", 
        x"cd", x"cd", x"cf", x"cc", x"d1", x"d0", x"cf", x"db", x"d1", x"d1", x"af", x"90", x"a7", x"d1", x"cd", 
        x"94", x"64", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"5e", x"5f", x"5e", x"75", x"bd", x"ec", x"f8", x"f7", x"f6", 
        x"f3", x"d9", x"a0", x"96", x"9d", x"aa", x"bd", x"ce", x"d4", x"cd", x"c8", x"c8", x"b0", x"9e", x"8e", 
        x"8f", x"ad", x"ae", x"a5", x"a2", x"9c", x"8f", x"7d", x"68", x"59", x"5b", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5d", x"5e", x"a0", x"e9", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", x"ed", x"ed", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ee", x"ed", x"ee", x"f0", x"ec", x"e3", x"cf", x"c6", x"d6", x"e5", x"e6", x"c6", 
        x"9c", x"7b", x"6f", x"72", x"77", x"7b", x"7c", x"7c", x"7b", x"79", x"7b", x"7e", x"7b", x"79", x"7c", 
        x"7c", x"7a", x"7c", x"7b", x"7a", x"7c", x"7c", x"7b", x"7b", x"7c", x"7d", x"7c", x"7b", x"7a", x"7a", 
        x"79", x"78", x"7a", x"7a", x"77", x"7a", x"79", x"7b", x"7b", x"79", x"7c", x"7c", x"7a", x"7b", x"7d", 
        x"7a", x"7a", x"7a", x"77", x"76", x"79", x"7a", x"7a", x"79", x"78", x"7a", x"7b", x"79", x"79", x"7c", 
        x"79", x"79", x"7a", x"77", x"7a", x"7a", x"7a", x"79", x"79", x"7a", x"7b", x"78", x"78", x"7c", x"78", 
        x"76", x"7b", x"7a", x"79", x"78", x"77", x"78", x"7a", x"78", x"76", x"77", x"76", x"78", x"7d", x"7b", 
        x"79", x"79", x"7a", x"7a", x"77", x"79", x"7c", x"7a", x"7b", x"7a", x"77", x"79", x"79", x"78", x"77", 
        x"78", x"78", x"78", x"78", x"78", x"79", x"79", x"78", x"76", x"77", x"78", x"78", x"77", x"76", x"77", 
        x"78", x"77", x"75", x"75", x"77", x"76", x"74", x"75", x"79", x"79", x"77", x"76", x"77", x"78", x"77", 
        x"77", x"73", x"71", x"74", x"79", x"77", x"78", x"76", x"77", x"74", x"75", x"78", x"77", x"75", x"75", 
        x"75", x"74", x"72", x"74", x"74", x"75", x"74", x"74", x"74", x"74", x"79", x"79", x"77", x"79", x"73", 
        x"74", x"77", x"73", x"74", x"77", x"77", x"75", x"77", x"77", x"75", x"78", x"76", x"74", x"77", x"75", 
        x"77", x"78", x"76", x"77", x"76", x"79", x"76", x"77", x"76", x"74", x"75", x"78", x"78", x"75", x"73", 
        x"75", x"78", x"77", x"75", x"76", x"75", x"74", x"76", x"76", x"77", x"77", x"77", x"76", x"76", x"76", 
        x"75", x"75", x"75", x"75", x"75", x"77", x"78", x"75", x"75", x"78", x"77", x"74", x"75", x"75", x"74", 
        x"73", x"73", x"73", x"73", x"72", x"73", x"75", x"76", x"76", x"75", x"74", x"71", x"74", x"72", x"6f", 
        x"70", x"71", x"70", x"71", x"72", x"73", x"74", x"75", x"75", x"70", x"6f", x"71", x"71", x"72", x"70", 
        x"6e", x"72", x"75", x"73", x"71", x"70", x"6f", x"71", x"73", x"73", x"72", x"71", x"70", x"6f", x"6f", 
        x"70", x"73", x"70", x"70", x"72", x"72", x"71", x"71", x"71", x"70", x"72", x"6f", x"71", x"71", x"72", 
        x"71", x"6f", x"6e", x"6c", x"70", x"74", x"73", x"71", x"70", x"70", x"72", x"6f", x"70", x"71", x"6f", 
        x"71", x"70", x"71", x"71", x"6e", x"71", x"6f", x"6e", x"6f", x"6d", x"6e", x"70", x"6f", x"6d", x"70", 
        x"72", x"73", x"6f", x"6e", x"71", x"6f", x"6f", x"6f", x"6e", x"6f", x"70", x"70", x"6f", x"71", x"71", 
        x"70", x"72", x"72", x"6f", x"6e", x"71", x"74", x"71", x"70", x"6f", x"6e", x"6e", x"6e", x"6e", x"6d", 
        x"6d", x"70", x"6c", x"6e", x"70", x"74", x"72", x"6f", x"6c", x"71", x"72", x"72", x"6e", x"6e", x"6b", 
        x"70", x"72", x"71", x"71", x"6e", x"6e", x"6e", x"6e", x"6e", x"6d", x"6c", x"6c", x"6c", x"6d", x"6e", 
        x"6e", x"6c", x"6d", x"70", x"70", x"6d", x"6d", x"6f", x"6e", x"6d", x"6d", x"6d", x"6c", x"6d", x"6e", 
        x"6c", x"6e", x"70", x"6e", x"6b", x"6b", x"6e", x"6f", x"70", x"6f", x"6e", x"6f", x"6f", x"6f", x"73", 
        x"74", x"70", x"6f", x"71", x"71", x"70", x"6e", x"70", x"70", x"6d", x"6f", x"70", x"6f", x"70", x"71", 
        x"71", x"70", x"6f", x"6f", x"71", x"70", x"6d", x"6e", x"70", x"6f", x"6f", x"70", x"70", x"6f", x"71", 
        x"72", x"70", x"6e", x"6f", x"70", x"6d", x"6d", x"6d", x"6b", x"6f", x"70", x"6f", x"70", x"71", x"71", 
        x"71", x"70", x"6f", x"70", x"71", x"71", x"71", x"71", x"71", x"71", x"71", x"71", x"71", x"71", x"70", 
        x"70", x"71", x"71", x"70", x"71", x"72", x"72", x"73", x"72", x"72", x"73", x"74", x"74", x"74", x"72", 
        x"72", x"73", x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"72", x"72", x"74", x"73", x"74", x"72", 
        x"75", x"74", x"73", x"74", x"74", x"74", x"74", x"74", x"74", x"74", x"74", x"74", x"77", x"78", x"70", 
        x"8e", x"d7", x"d1", x"d0", x"d0", x"d4", x"de", x"d4", x"cd", x"cd", x"ce", x"ce", x"ce", x"cf", x"d0", 
        x"d1", x"d0", x"ce", x"cd", x"cd", x"cf", x"d0", x"d0", x"d0", x"d1", x"d0", x"ce", x"cc", x"cc", x"ce", 
        x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", x"cf", x"d0", x"d0", x"d0", x"cf", x"cf", x"ce", x"ce", x"ce", 
        x"d2", x"cd", x"cd", x"cf", x"d2", x"cc", x"d1", x"dd", x"be", x"94", x"89", x"b8", x"d4", x"d1", x"c6", 
        x"94", x"64", x"5d", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"60", x"5c", x"77", x"bd", x"f0", x"f7", x"f8", x"f7", x"f7", 
        x"e6", x"9b", x"5f", x"5e", x"61", x"60", x"69", x"75", x"7a", x"74", x"6f", x"73", x"64", x"5e", x"5c", 
        x"5e", x"68", x"61", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5c", x"5d", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5d", x"5f", x"9d", x"e8", 
        x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"ec", x"ef", x"eb", x"e4", x"d9", x"d5", x"d4", x"d9", 
        x"e0", x"d4", x"b2", x"8e", x"74", x"6e", x"77", x"7b", x"80", x"81", x"7b", x"79", x"7c", x"7d", x"7e", 
        x"7c", x"7b", x"7e", x"7d", x"7d", x"7e", x"7b", x"7c", x"7d", x"7d", x"7d", x"7c", x"7b", x"7d", x"7d", 
        x"7c", x"7d", x"7d", x"7b", x"79", x"79", x"78", x"7b", x"7b", x"7a", x"7b", x"7a", x"79", x"7a", x"7a", 
        x"79", x"7a", x"7b", x"79", x"76", x"77", x"79", x"79", x"79", x"79", x"7b", x"7c", x"7a", x"7a", x"7c", 
        x"7a", x"7b", x"7d", x"7a", x"79", x"79", x"79", x"79", x"79", x"7a", x"7b", x"79", x"7a", x"7c", x"79", 
        x"78", x"7b", x"7a", x"78", x"78", x"77", x"79", x"7a", x"7a", x"78", x"7b", x"79", x"79", x"7c", x"79", 
        x"79", x"79", x"7a", x"7a", x"78", x"79", x"7a", x"7a", x"7a", x"7a", x"77", x"78", x"79", x"78", x"78", 
        x"7a", x"7b", x"7a", x"77", x"77", x"78", x"78", x"78", x"78", x"78", x"78", x"78", x"78", x"78", x"78", 
        x"78", x"79", x"78", x"77", x"79", x"78", x"76", x"77", x"79", x"77", x"77", x"78", x"77", x"78", x"77", 
        x"77", x"75", x"76", x"75", x"77", x"77", x"77", x"74", x"76", x"74", x"75", x"78", x"77", x"77", x"77", 
        x"75", x"76", x"77", x"79", x"77", x"77", x"76", x"76", x"76", x"75", x"78", x"77", x"76", x"79", x"75", 
        x"76", x"7a", x"79", x"77", x"7a", x"7a", x"77", x"79", x"7a", x"78", x"79", x"77", x"76", x"78", x"77", 
        x"76", x"75", x"74", x"75", x"74", x"76", x"78", x"76", x"76", x"77", x"76", x"75", x"76", x"76", x"76", 
        x"77", x"77", x"75", x"73", x"74", x"73", x"73", x"76", x"76", x"74", x"74", x"76", x"76", x"76", x"75", 
        x"74", x"75", x"76", x"76", x"77", x"78", x"78", x"74", x"73", x"75", x"76", x"75", x"75", x"76", x"76", 
        x"75", x"74", x"73", x"73", x"75", x"74", x"73", x"73", x"74", x"73", x"72", x"71", x"73", x"72", x"70", 
        x"72", x"72", x"72", x"74", x"74", x"73", x"71", x"72", x"74", x"73", x"70", x"70", x"73", x"74", x"72", 
        x"71", x"71", x"71", x"6f", x"6e", x"70", x"71", x"72", x"74", x"74", x"71", x"71", x"72", x"71", x"70", 
        x"70", x"72", x"73", x"72", x"71", x"70", x"70", x"71", x"72", x"71", x"72", x"71", x"73", x"72", x"71", 
        x"72", x"72", x"70", x"6d", x"6f", x"71", x"70", x"70", x"70", x"70", x"70", x"6f", x"70", x"70", x"6e", 
        x"70", x"6f", x"6f", x"70", x"6f", x"6f", x"6d", x"6e", x"72", x"70", x"6e", x"6e", x"70", x"71", x"70", 
        x"6f", x"6f", x"6c", x"6c", x"6f", x"6d", x"6d", x"6e", x"6e", x"6f", x"70", x"70", x"71", x"71", x"72", 
        x"72", x"70", x"6f", x"6f", x"6f", x"6f", x"70", x"72", x"71", x"6f", x"6f", x"6f", x"70", x"70", x"6f", 
        x"6e", x"71", x"6d", x"6f", x"6e", x"70", x"70", x"6f", x"6c", x"6f", x"70", x"71", x"70", x"6e", x"6e", 
        x"71", x"72", x"6f", x"72", x"70", x"6e", x"6f", x"6d", x"6d", x"6e", x"6e", x"6d", x"6d", x"6e", x"6e", 
        x"6c", x"6a", x"6c", x"6f", x"71", x"70", x"6e", x"6f", x"6f", x"6e", x"6e", x"6e", x"6d", x"6d", x"6d", 
        x"6d", x"6f", x"70", x"6d", x"6c", x"6e", x"6d", x"6f", x"6e", x"6f", x"70", x"6d", x"6f", x"6f", x"71", 
        x"72", x"71", x"70", x"71", x"71", x"6e", x"70", x"73", x"71", x"6c", x"6c", x"6f", x"6e", x"6d", x"6f", 
        x"70", x"70", x"70", x"70", x"71", x"70", x"6c", x"6d", x"70", x"70", x"6f", x"70", x"70", x"6f", x"71", 
        x"71", x"6f", x"6e", x"6f", x"71", x"6f", x"6d", x"6e", x"6e", x"70", x"6f", x"71", x"71", x"6f", x"6e", 
        x"6f", x"70", x"72", x"72", x"72", x"72", x"71", x"71", x"71", x"71", x"72", x"72", x"71", x"71", x"71", 
        x"71", x"71", x"70", x"70", x"71", x"72", x"73", x"73", x"73", x"72", x"70", x"73", x"75", x"75", x"75", 
        x"75", x"74", x"74", x"73", x"72", x"73", x"74", x"74", x"73", x"74", x"75", x"75", x"73", x"75", x"76", 
        x"77", x"74", x"73", x"73", x"73", x"73", x"74", x"74", x"74", x"73", x"75", x"76", x"7a", x"79", x"70", 
        x"8d", x"d8", x"d3", x"d1", x"d1", x"d4", x"dd", x"d2", x"cd", x"ce", x"ce", x"cd", x"cd", x"ce", x"d0", 
        x"d1", x"d1", x"cf", x"cd", x"cd", x"ce", x"d0", x"d0", x"cf", x"d0", x"d0", x"ce", x"cc", x"cb", x"ce", 
        x"d1", x"d0", x"d0", x"d2", x"d1", x"cf", x"ce", x"d0", x"d0", x"d0", x"cf", x"cf", x"cf", x"ce", x"cd", 
        x"d0", x"ce", x"cc", x"ce", x"d0", x"d3", x"d7", x"bf", x"88", x"93", x"c5", x"d5", x"d1", x"cc", x"c6", 
        x"98", x"64", x"5c", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"6a", x"b1", x"ea", x"f7", x"f8", x"f8", x"f8", x"f0", 
        x"bd", x"6d", x"5b", x"5d", x"5e", x"5d", x"5b", x"5a", x"5b", x"5c", x"5b", x"5a", x"5b", x"5d", x"5b", 
        x"59", x"5b", x"5b", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", 
        x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5d", x"5e", x"98", x"e5", 
        x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"e8", x"dd", x"d1", 
        x"d1", x"d9", x"e1", x"d6", x"b7", x"90", x"78", x"72", x"78", x"7b", x"78", x"79", x"7a", x"7b", x"7e", 
        x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7a", x"7d", x"7e", x"7d", x"7c", x"7c", x"7c", x"7f", x"7b", 
        x"7a", x"7a", x"7a", x"7a", x"7c", x"7b", x"7a", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7a", x"79", 
        x"78", x"7a", x"7b", x"7a", x"79", x"79", x"79", x"79", x"78", x"78", x"78", x"79", x"79", x"7a", x"7b", 
        x"7a", x"7b", x"7c", x"7a", x"79", x"7a", x"79", x"79", x"78", x"79", x"7a", x"7a", x"7a", x"7b", x"79", 
        x"79", x"7c", x"7a", x"78", x"78", x"79", x"7a", x"7a", x"7a", x"79", x"7c", x"7b", x"7a", x"7a", x"78", 
        x"79", x"7a", x"7a", x"79", x"78", x"79", x"7a", x"7a", x"7a", x"7a", x"79", x"7a", x"7a", x"79", x"78", 
        x"79", x"7a", x"7a", x"78", x"77", x"78", x"79", x"79", x"78", x"77", x"76", x"76", x"77", x"78", x"78", 
        x"78", x"77", x"76", x"76", x"77", x"76", x"75", x"75", x"77", x"76", x"78", x"79", x"79", x"78", x"77", 
        x"78", x"76", x"77", x"75", x"75", x"75", x"76", x"74", x"76", x"75", x"75", x"77", x"77", x"77", x"77", 
        x"77", x"78", x"77", x"77", x"76", x"78", x"79", x"78", x"77", x"77", x"7a", x"78", x"75", x"76", x"74", 
        x"76", x"7a", x"78", x"77", x"78", x"78", x"76", x"76", x"78", x"78", x"78", x"79", x"7a", x"7b", x"78", 
        x"76", x"75", x"75", x"77", x"77", x"78", x"77", x"74", x"75", x"77", x"75", x"73", x"75", x"75", x"76", 
        x"78", x"77", x"74", x"73", x"75", x"76", x"76", x"75", x"76", x"77", x"77", x"76", x"75", x"76", x"75", 
        x"75", x"75", x"76", x"78", x"78", x"77", x"77", x"74", x"72", x"74", x"74", x"75", x"75", x"74", x"73", 
        x"73", x"74", x"75", x"76", x"73", x"73", x"72", x"73", x"73", x"73", x"72", x"70", x"72", x"72", x"71", 
        x"74", x"73", x"73", x"73", x"72", x"71", x"6e", x"6f", x"73", x"74", x"72", x"71", x"74", x"73", x"71", 
        x"72", x"73", x"72", x"6f", x"70", x"71", x"71", x"72", x"72", x"72", x"70", x"72", x"73", x"73", x"71", 
        x"71", x"72", x"75", x"74", x"71", x"6f", x"71", x"72", x"73", x"71", x"70", x"71", x"73", x"72", x"6f", 
        x"71", x"72", x"70", x"6e", x"70", x"72", x"71", x"70", x"71", x"70", x"70", x"70", x"71", x"6f", x"6e", 
        x"71", x"6f", x"6e", x"70", x"70", x"6e", x"6d", x"70", x"72", x"72", x"70", x"6e", x"70", x"73", x"71", 
        x"6f", x"70", x"6e", x"6e", x"71", x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"70", x"72", x"71", x"6f", 
        x"6f", x"6f", x"70", x"70", x"70", x"6f", x"70", x"73", x"72", x"70", x"6f", x"6f", x"70", x"71", x"71", 
        x"6f", x"71", x"6f", x"70", x"6e", x"6e", x"70", x"70", x"6e", x"6f", x"6f", x"6f", x"6f", x"6f", x"70", 
        x"6f", x"6f", x"6d", x"71", x"70", x"6c", x"6f", x"6c", x"6c", x"6f", x"70", x"6f", x"6e", x"6f", x"6f", 
        x"6f", x"6f", x"6f", x"6e", x"6e", x"6f", x"6f", x"70", x"6f", x"6f", x"6e", x"6e", x"6d", x"6c", x"6b", 
        x"6e", x"71", x"70", x"6c", x"6e", x"71", x"6c", x"6e", x"6c", x"6e", x"6f", x"6b", x"6d", x"71", x"70", 
        x"6e", x"6e", x"6e", x"6e", x"6d", x"6d", x"6d", x"6d", x"6d", x"6e", x"6d", x"6d", x"6b", x"6b", x"6d", 
        x"6f", x"70", x"71", x"71", x"70", x"70", x"6f", x"72", x"72", x"70", x"6f", x"72", x"71", x"70", x"6f", 
        x"6f", x"6f", x"70", x"70", x"71", x"71", x"70", x"70", x"71", x"70", x"6e", x"71", x"72", x"71", x"71", 
        x"70", x"6f", x"6f", x"72", x"73", x"72", x"71", x"71", x"71", x"71", x"72", x"73", x"71", x"71", x"71", 
        x"72", x"71", x"70", x"70", x"70", x"71", x"72", x"73", x"73", x"72", x"70", x"74", x"75", x"73", x"73", 
        x"74", x"72", x"72", x"71", x"71", x"73", x"75", x"76", x"75", x"76", x"76", x"74", x"72", x"74", x"76", 
        x"74", x"73", x"76", x"74", x"75", x"75", x"76", x"77", x"77", x"74", x"76", x"76", x"79", x"79", x"6f", 
        x"8c", x"d7", x"d3", x"d2", x"d1", x"d3", x"da", x"cf", x"cd", x"ce", x"ce", x"cd", x"cd", x"ce", x"d0", 
        x"cf", x"d0", x"d0", x"ce", x"cd", x"ce", x"d0", x"cf", x"cd", x"ce", x"cf", x"cd", x"cc", x"cd", x"d0", 
        x"d1", x"d0", x"d0", x"d2", x"d3", x"d0", x"ce", x"d0", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", 
        x"d4", x"ca", x"ce", x"d6", x"d8", x"c9", x"98", x"97", x"b3", x"d1", x"d4", x"d1", x"d3", x"d0", x"c9", 
        x"9e", x"65", x"5c", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"61", x"5d", x"5a", x"77", x"d8", x"f7", x"f7", x"fa", x"f7", x"f6", x"d8", 
        x"82", x"5f", x"60", x"5c", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5c", x"5b", x"5c", x"5d", x"5e", 
        x"5f", x"5c", x"5e", x"5d", x"5d", x"5d", x"5d", x"5c", x"5c", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5d", x"5e", x"92", x"e2", 
        x"ed", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ed", x"ec", x"ef", x"ef", x"ee", x"ed", x"eb", 
        x"e1", x"d6", x"c4", x"c5", x"d8", x"e2", x"cf", x"a7", x"79", x"65", x"71", x"7e", x"7d", x"7c", x"7f", 
        x"7e", x"7d", x"7e", x"7e", x"7c", x"7a", x"7c", x"7e", x"7e", x"7c", x"7c", x"7c", x"7d", x"7a", x"78", 
        x"79", x"7b", x"7a", x"79", x"7b", x"7d", x"7c", x"7b", x"7b", x"7c", x"7d", x"7e", x"7e", x"7b", x"79", 
        x"79", x"7a", x"7a", x"7a", x"7a", x"7a", x"7a", x"7a", x"79", x"79", x"79", x"79", x"79", x"7a", x"7b", 
        x"7b", x"7a", x"79", x"79", x"7a", x"7b", x"7b", x"79", x"78", x"77", x"78", x"79", x"7b", x"7a", x"78", 
        x"79", x"7a", x"79", x"79", x"7a", x"7a", x"7b", x"7a", x"79", x"79", x"7b", x"7a", x"7a", x"7a", x"79", 
        x"7a", x"7c", x"7a", x"79", x"78", x"78", x"79", x"7a", x"7a", x"7a", x"7b", x"7c", x"7b", x"7a", x"78", 
        x"78", x"79", x"79", x"79", x"78", x"79", x"7a", x"79", x"78", x"77", x"76", x"75", x"77", x"78", x"78", 
        x"77", x"78", x"78", x"78", x"77", x"77", x"77", x"77", x"77", x"76", x"7a", x"7b", x"79", x"78", x"76", 
        x"78", x"77", x"76", x"77", x"76", x"75", x"75", x"76", x"78", x"78", x"77", x"76", x"76", x"77", x"77", 
        x"76", x"77", x"77", x"78", x"76", x"78", x"78", x"76", x"75", x"76", x"7b", x"7a", x"77", x"78", x"74", 
        x"75", x"77", x"75", x"74", x"75", x"77", x"78", x"79", x"78", x"77", x"75", x"76", x"78", x"79", x"77", 
        x"76", x"76", x"78", x"79", x"79", x"78", x"75", x"74", x"75", x"77", x"76", x"75", x"75", x"74", x"77", 
        x"78", x"76", x"75", x"75", x"77", x"78", x"75", x"73", x"75", x"78", x"78", x"74", x"74", x"76", x"76", 
        x"75", x"75", x"77", x"79", x"78", x"77", x"76", x"76", x"74", x"73", x"73", x"75", x"78", x"76", x"74", 
        x"73", x"74", x"76", x"77", x"71", x"73", x"75", x"75", x"73", x"73", x"74", x"71", x"72", x"72", x"71", 
        x"73", x"71", x"71", x"74", x"74", x"73", x"6e", x"6e", x"70", x"71", x"71", x"72", x"74", x"71", x"70", 
        x"73", x"74", x"73", x"72", x"72", x"73", x"72", x"71", x"6f", x"6f", x"70", x"72", x"72", x"71", x"71", 
        x"71", x"72", x"73", x"72", x"70", x"70", x"73", x"74", x"74", x"73", x"71", x"73", x"75", x"73", x"71", 
        x"73", x"75", x"73", x"71", x"72", x"72", x"70", x"6f", x"71", x"70", x"6f", x"71", x"72", x"6f", x"6f", 
        x"72", x"72", x"71", x"71", x"70", x"6d", x"6d", x"71", x"71", x"75", x"75", x"70", x"70", x"72", x"72", 
        x"71", x"73", x"71", x"72", x"73", x"71", x"72", x"71", x"6f", x"6f", x"6e", x"70", x"72", x"71", x"6d", 
        x"6d", x"6f", x"72", x"72", x"71", x"70", x"71", x"74", x"72", x"70", x"6e", x"6d", x"6e", x"70", x"72", 
        x"70", x"6f", x"6e", x"71", x"70", x"6f", x"6f", x"6f", x"6f", x"6f", x"6d", x"6c", x"6b", x"70", x"71", 
        x"70", x"71", x"70", x"73", x"71", x"70", x"71", x"6d", x"6c", x"6f", x"6f", x"6f", x"6f", x"6e", x"6b", 
        x"6b", x"6e", x"6e", x"6b", x"6b", x"6e", x"6f", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", x"6e", 
        x"6e", x"6f", x"6f", x"6d", x"6d", x"6e", x"6e", x"6f", x"6e", x"70", x"71", x"6e", x"6c", x"6c", x"6e", 
        x"6d", x"6b", x"6b", x"6d", x"70", x"6f", x"6f", x"6e", x"6f", x"72", x"71", x"70", x"72", x"72", x"70", 
        x"6f", x"70", x"71", x"72", x"70", x"6e", x"71", x"72", x"70", x"6e", x"6f", x"70", x"70", x"71", x"70", 
        x"6f", x"70", x"70", x"6f", x"72", x"73", x"70", x"70", x"70", x"6f", x"6e", x"70", x"71", x"71", x"71", 
        x"71", x"71", x"71", x"72", x"72", x"72", x"71", x"71", x"71", x"71", x"72", x"72", x"71", x"71", x"71", 
        x"73", x"72", x"72", x"71", x"71", x"72", x"73", x"74", x"73", x"72", x"71", x"73", x"74", x"72", x"72", 
        x"73", x"72", x"71", x"71", x"71", x"73", x"75", x"75", x"75", x"76", x"78", x"75", x"73", x"73", x"77", 
        x"73", x"73", x"75", x"74", x"74", x"74", x"74", x"75", x"76", x"77", x"76", x"74", x"76", x"77", x"6f", 
        x"8d", x"d7", x"d1", x"cf", x"cf", x"d2", x"db", x"d1", x"ce", x"ce", x"ce", x"ce", x"cd", x"cd", x"cf", 
        x"cf", x"d0", x"cf", x"cf", x"ce", x"ce", x"cf", x"ce", x"cd", x"ce", x"ce", x"cd", x"cd", x"cf", x"d1", 
        x"d1", x"cf", x"cf", x"d1", x"d2", x"cf", x"cd", x"cf", x"d0", x"d1", x"d1", x"d1", x"d2", x"d1", x"cc", 
        x"cd", x"d0", x"cf", x"ce", x"af", x"95", x"a4", x"cc", x"d7", x"d2", x"d1", x"cd", x"ce", x"cf", x"ca", 
        x"a0", x"64", x"5c", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"60", x"5f", x"5d", x"85", x"e0", x"f5", x"f9", x"f8", x"f9", x"ee", x"a7", 
        x"63", x"60", x"5f", x"5e", x"60", x"5d", x"5c", x"5e", x"5f", x"5e", x"5d", x"5e", x"61", x"60", x"5e", 
        x"5d", x"5d", x"5f", x"5d", x"5d", x"5d", x"5d", x"5d", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5e", x"5e", x"8c", x"df", 
        x"ec", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ec", x"ed", x"ec", x"ec", x"ed", x"ed", x"ec", x"ee", 
        x"f0", x"ec", x"e3", x"d7", x"cc", x"c8", x"d7", x"de", x"d3", x"b5", x"8d", x"71", x"71", x"7a", x"7d", 
        x"7d", x"7e", x"7c", x"7d", x"7e", x"7d", x"7d", x"7e", x"7d", x"7c", x"7c", x"7d", x"7e", x"7b", x"7a", 
        x"7b", x"7c", x"7b", x"7b", x"7d", x"7a", x"7b", x"7a", x"7b", x"7c", x"7b", x"7b", x"7c", x"7b", x"7b", 
        x"7b", x"7a", x"79", x"7a", x"7b", x"7b", x"7a", x"7a", x"7a", x"7a", x"79", x"79", x"7c", x"7d", x"7c", 
        x"7d", x"7c", x"79", x"7a", x"7b", x"7b", x"7c", x"7a", x"78", x"78", x"78", x"79", x"7b", x"78", x"78", 
        x"7a", x"7a", x"79", x"7a", x"7b", x"7a", x"7b", x"7a", x"79", x"78", x"79", x"79", x"7a", x"7a", x"79", 
        x"7b", x"7c", x"79", x"79", x"79", x"78", x"79", x"7b", x"7b", x"7a", x"79", x"7a", x"7b", x"7a", x"78", 
        x"79", x"7a", x"79", x"79", x"79", x"7a", x"7a", x"79", x"77", x"79", x"79", x"79", x"79", x"7a", x"7a", 
        x"79", x"78", x"78", x"78", x"77", x"77", x"77", x"77", x"78", x"78", x"79", x"7a", x"7a", x"78", x"77", 
        x"79", x"77", x"75", x"77", x"77", x"77", x"76", x"79", x"79", x"7a", x"78", x"76", x"76", x"77", x"77", 
        x"77", x"78", x"77", x"78", x"77", x"78", x"78", x"77", x"77", x"76", x"79", x"78", x"77", x"7a", x"78", 
        x"77", x"77", x"75", x"74", x"75", x"78", x"7a", x"79", x"77", x"77", x"74", x"75", x"77", x"77", x"78", 
        x"78", x"77", x"77", x"76", x"76", x"74", x"76", x"75", x"76", x"77", x"77", x"77", x"77", x"76", x"78", 
        x"79", x"76", x"74", x"76", x"76", x"76", x"77", x"77", x"77", x"77", x"76", x"75", x"76", x"77", x"76", 
        x"76", x"76", x"78", x"78", x"78", x"75", x"74", x"76", x"75", x"74", x"74", x"75", x"74", x"74", x"74", 
        x"74", x"74", x"74", x"74", x"72", x"74", x"75", x"73", x"70", x"71", x"74", x"72", x"73", x"72", x"73", 
        x"74", x"70", x"70", x"75", x"76", x"75", x"71", x"71", x"73", x"72", x"71", x"71", x"73", x"73", x"73", 
        x"73", x"73", x"73", x"73", x"73", x"74", x"73", x"72", x"71", x"70", x"72", x"72", x"72", x"72", x"71", 
        x"71", x"73", x"72", x"72", x"71", x"72", x"72", x"73", x"73", x"71", x"6f", x"72", x"72", x"72", x"71", 
        x"71", x"74", x"75", x"71", x"70", x"70", x"6f", x"71", x"73", x"72", x"71", x"73", x"72", x"71", x"72", 
        x"72", x"71", x"70", x"70", x"70", x"6f", x"72", x"73", x"70", x"74", x"75", x"71", x"6f", x"70", x"71", 
        x"70", x"74", x"73", x"72", x"73", x"71", x"71", x"71", x"70", x"6f", x"6e", x"6f", x"71", x"70", x"71", 
        x"72", x"6f", x"6f", x"71", x"72", x"70", x"70", x"73", x"73", x"71", x"6f", x"6e", x"6e", x"6f", x"73", 
        x"71", x"6e", x"6f", x"71", x"72", x"72", x"71", x"70", x"73", x"72", x"71", x"6f", x"6d", x"71", x"70", 
        x"6d", x"6f", x"70", x"70", x"6e", x"6f", x"70", x"6e", x"6d", x"6e", x"6e", x"6f", x"6f", x"6e", x"6e", 
        x"70", x"70", x"6f", x"6d", x"6c", x"6e", x"6e", x"6b", x"6c", x"6d", x"6d", x"6e", x"6f", x"70", x"6f", 
        x"6e", x"6e", x"6e", x"6d", x"6c", x"6e", x"70", x"6f", x"70", x"71", x"72", x"71", x"6d", x"6a", x"6d", 
        x"6e", x"6c", x"6e", x"72", x"72", x"6c", x"6e", x"6f", x"6e", x"6f", x"6d", x"6f", x"75", x"74", x"71", 
        x"6f", x"70", x"71", x"72", x"72", x"71", x"73", x"71", x"70", x"72", x"72", x"70", x"70", x"71", x"6f", 
        x"6e", x"70", x"70", x"6f", x"71", x"74", x"70", x"70", x"70", x"6d", x"6f", x"73", x"73", x"72", x"70", 
        x"70", x"70", x"70", x"70", x"71", x"72", x"72", x"72", x"72", x"72", x"71", x"71", x"71", x"71", x"72", 
        x"73", x"74", x"74", x"72", x"72", x"73", x"73", x"74", x"73", x"72", x"71", x"72", x"73", x"74", x"72", 
        x"72", x"74", x"72", x"72", x"72", x"73", x"73", x"73", x"73", x"75", x"78", x"76", x"75", x"75", x"79", 
        x"75", x"75", x"77", x"77", x"77", x"77", x"77", x"76", x"76", x"75", x"75", x"73", x"76", x"77", x"6f", 
        x"8e", x"d8", x"d2", x"d0", x"cf", x"d2", x"db", x"d2", x"ce", x"cf", x"cf", x"cf", x"ce", x"cd", x"cf", 
        x"d0", x"cf", x"ce", x"ce", x"cf", x"cf", x"d0", x"ce", x"ce", x"cf", x"cf", x"ce", x"ce", x"cf", x"d0", 
        x"d0", x"cf", x"cf", x"d0", x"d0", x"ce", x"ce", x"cf", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", x"cf", 
        x"cb", x"d3", x"c4", x"93", x"91", x"bf", x"d0", x"dc", x"d5", x"d2", x"d0", x"cd", x"d0", x"cf", x"c8", 
        x"a0", x"64", x"5d", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5c", x"60", x"64", x"ab", x"ed", x"fa", x"fa", x"f6", x"f7", x"e3", x"82", 
        x"61", x"5c", x"5f", x"5d", x"5c", x"5f", x"61", x"62", x"60", x"5f", x"5f", x"60", x"5f", x"5e", x"5f", 
        x"5e", x"5d", x"5d", x"5c", x"5e", x"60", x"5f", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5e", x"5e", x"89", x"dd", 
        x"ec", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ee", x"ed", x"ee", x"ef", x"ef", x"ee", x"eb", x"ef", x"ed", x"ea", x"ee", x"ef", x"eb", x"ec", 
        x"ee", x"eb", x"ed", x"ef", x"e7", x"de", x"cf", x"ca", x"d4", x"e1", x"dc", x"c0", x"8d", x"71", x"6a", 
        x"75", x"80", x"7f", x"7b", x"7e", x"80", x"7d", x"7d", x"7d", x"7d", x"7e", x"7d", x"7d", x"7f", x"7f", 
        x"7c", x"7a", x"7a", x"7d", x"7f", x"7a", x"7c", x"7b", x"7c", x"7d", x"7b", x"7b", x"7b", x"7a", x"7c", 
        x"7d", x"7b", x"79", x"7b", x"7d", x"7b", x"7a", x"7a", x"7b", x"7a", x"79", x"7a", x"7e", x"7d", x"7a", 
        x"7c", x"7b", x"7a", x"7c", x"7a", x"7b", x"7c", x"7c", x"7a", x"7a", x"7a", x"7a", x"7c", x"79", x"79", 
        x"7c", x"7a", x"79", x"7a", x"7a", x"79", x"7a", x"7b", x"7a", x"78", x"79", x"79", x"7a", x"79", x"78", 
        x"7b", x"7b", x"78", x"7a", x"7a", x"78", x"79", x"7c", x"7c", x"79", x"79", x"7a", x"7a", x"79", x"78", 
        x"78", x"79", x"79", x"78", x"78", x"78", x"79", x"78", x"77", x"79", x"7a", x"7a", x"7a", x"79", x"79", 
        x"79", x"77", x"78", x"78", x"76", x"76", x"77", x"76", x"78", x"78", x"79", x"7a", x"7a", x"79", x"77", 
        x"7a", x"79", x"77", x"76", x"76", x"79", x"76", x"78", x"78", x"7a", x"78", x"75", x"77", x"79", x"79", 
        x"7a", x"79", x"77", x"77", x"77", x"79", x"7a", x"7a", x"7a", x"77", x"79", x"78", x"75", x"78", x"79", 
        x"78", x"76", x"76", x"76", x"77", x"78", x"79", x"77", x"76", x"78", x"77", x"79", x"79", x"77", x"7a", 
        x"79", x"78", x"77", x"75", x"77", x"76", x"78", x"75", x"75", x"77", x"76", x"75", x"79", x"78", x"79", 
        x"79", x"76", x"76", x"78", x"78", x"77", x"79", x"7a", x"7a", x"77", x"76", x"77", x"78", x"78", x"78", 
        x"77", x"77", x"77", x"77", x"77", x"75", x"73", x"75", x"76", x"77", x"76", x"77", x"73", x"73", x"75", 
        x"76", x"76", x"76", x"76", x"74", x"74", x"75", x"75", x"75", x"76", x"76", x"73", x"73", x"73", x"75", 
        x"76", x"72", x"71", x"73", x"74", x"72", x"71", x"72", x"75", x"73", x"72", x"72", x"72", x"73", x"74", 
        x"73", x"73", x"73", x"73", x"73", x"74", x"74", x"73", x"73", x"72", x"71", x"72", x"73", x"72", x"71", 
        x"71", x"72", x"72", x"73", x"72", x"72", x"71", x"70", x"70", x"72", x"71", x"74", x"73", x"74", x"75", 
        x"72", x"73", x"70", x"6f", x"70", x"70", x"70", x"71", x"73", x"70", x"70", x"72", x"6f", x"70", x"72", 
        x"70", x"71", x"72", x"70", x"71", x"70", x"72", x"70", x"72", x"72", x"71", x"71", x"70", x"6f", x"70", 
        x"70", x"74", x"73", x"72", x"73", x"6f", x"70", x"72", x"71", x"70", x"6f", x"6e", x"6e", x"70", x"73", 
        x"74", x"70", x"6f", x"70", x"72", x"71", x"70", x"71", x"71", x"72", x"72", x"71", x"6f", x"6f", x"73", 
        x"72", x"70", x"70", x"71", x"72", x"72", x"70", x"6e", x"70", x"70", x"70", x"70", x"6e", x"71", x"6e", 
        x"70", x"72", x"73", x"71", x"6f", x"71", x"70", x"6f", x"6e", x"6d", x"6e", x"6e", x"6e", x"6e", x"6f", 
        x"6f", x"6e", x"6d", x"6e", x"6e", x"70", x"70", x"6e", x"6d", x"6d", x"6d", x"6d", x"6c", x"6c", x"6d", 
        x"6e", x"6f", x"6e", x"6c", x"6d", x"71", x"6f", x"6e", x"6f", x"70", x"70", x"71", x"6d", x"70", x"71", 
        x"6f", x"6e", x"72", x"73", x"6e", x"6c", x"6f", x"6c", x"6c", x"6f", x"6f", x"6e", x"71", x"71", x"70", 
        x"6f", x"70", x"72", x"72", x"70", x"70", x"71", x"6e", x"6e", x"73", x"72", x"6e", x"72", x"71", x"6d", 
        x"6c", x"6f", x"72", x"71", x"71", x"74", x"71", x"71", x"70", x"6d", x"6e", x"6f", x"70", x"71", x"72", 
        x"72", x"72", x"71", x"70", x"71", x"72", x"73", x"73", x"73", x"73", x"71", x"71", x"72", x"72", x"72", 
        x"72", x"75", x"75", x"73", x"74", x"74", x"74", x"73", x"73", x"73", x"73", x"74", x"76", x"76", x"72", 
        x"71", x"72", x"73", x"73", x"73", x"72", x"71", x"71", x"72", x"72", x"75", x"75", x"74", x"74", x"78", 
        x"75", x"75", x"76", x"76", x"76", x"76", x"76", x"74", x"73", x"72", x"74", x"75", x"78", x"77", x"6e", 
        x"8b", x"d8", x"d5", x"d3", x"d2", x"d4", x"db", x"d0", x"ce", x"cf", x"d1", x"cf", x"ce", x"ce", x"cf", 
        x"d0", x"cf", x"cd", x"cd", x"ce", x"d0", x"d0", x"cf", x"ce", x"d0", x"d0", x"d0", x"ce", x"cf", x"ce", 
        x"cf", x"ce", x"ce", x"cf", x"ce", x"ce", x"ce", x"d0", x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"d3", 
        x"d1", x"af", x"90", x"a4", x"ca", x"d0", x"ca", x"d9", x"d3", x"d0", x"d0", x"d2", x"d1", x"cf", x"c8", 
        x"a0", x"64", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"6f", x"d7", x"f6", x"fa", x"fa", x"f9", x"f7", x"cd", x"6c", 
        x"5f", x"61", x"60", x"5f", x"5e", x"5d", x"5d", x"5d", x"5d", x"5c", x"5d", x"5e", x"5e", x"5d", x"5e", 
        x"5d", x"5e", x"5c", x"5c", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5e", x"5e", x"87", x"dc", 
        x"ec", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ee", x"ed", x"ee", x"ef", x"ef", x"ee", x"eb", x"ea", x"ea", x"ec", x"ed", x"ec", x"ee", x"ed", 
        x"eb", x"eb", x"eb", x"ed", x"f0", x"ed", x"ec", x"e3", x"d2", x"c4", x"ca", x"dc", x"dc", x"c3", x"9d", 
        x"7b", x"71", x"74", x"79", x"7c", x"7c", x"7d", x"7e", x"7e", x"7e", x"7f", x"7b", x"7b", x"7e", x"7f", 
        x"7e", x"7b", x"7a", x"7b", x"7b", x"7c", x"7e", x"7b", x"7b", x"7d", x"7c", x"7d", x"7a", x"78", x"7c", 
        x"7d", x"7c", x"7a", x"7d", x"7d", x"7a", x"79", x"7a", x"7d", x"7e", x"7d", x"7c", x"7c", x"7b", x"78", 
        x"7a", x"7a", x"7a", x"7c", x"79", x"7a", x"7b", x"7c", x"7c", x"7c", x"7c", x"7a", x"7c", x"7a", x"7a", 
        x"7d", x"7b", x"7a", x"7a", x"78", x"78", x"79", x"7b", x"7b", x"79", x"7a", x"7b", x"7b", x"79", x"77", 
        x"79", x"7a", x"79", x"7b", x"7b", x"78", x"79", x"7c", x"7b", x"79", x"7a", x"7b", x"7a", x"79", x"78", 
        x"78", x"78", x"78", x"77", x"77", x"77", x"78", x"78", x"78", x"77", x"78", x"79", x"78", x"77", x"76", 
        x"76", x"78", x"7a", x"7a", x"78", x"78", x"7a", x"79", x"79", x"78", x"78", x"79", x"79", x"7a", x"78", 
        x"7a", x"79", x"78", x"76", x"75", x"7a", x"77", x"76", x"78", x"7a", x"78", x"76", x"77", x"7a", x"7a", 
        x"79", x"79", x"78", x"79", x"7a", x"79", x"77", x"77", x"78", x"78", x"7b", x"79", x"76", x"77", x"78", 
        x"76", x"75", x"75", x"76", x"76", x"76", x"79", x"79", x"79", x"7b", x"79", x"79", x"77", x"74", x"7a", 
        x"7a", x"79", x"78", x"77", x"7b", x"7b", x"7a", x"76", x"76", x"78", x"75", x"74", x"79", x"76", x"77", 
        x"77", x"75", x"76", x"7a", x"79", x"77", x"77", x"77", x"76", x"76", x"75", x"75", x"77", x"79", x"78", 
        x"78", x"78", x"78", x"77", x"76", x"75", x"72", x"73", x"76", x"77", x"78", x"78", x"75", x"75", x"74", 
        x"74", x"74", x"74", x"74", x"71", x"71", x"73", x"76", x"79", x"77", x"75", x"73", x"73", x"74", x"77", 
        x"77", x"73", x"73", x"73", x"72", x"71", x"6f", x"71", x"73", x"72", x"72", x"73", x"70", x"71", x"73", 
        x"73", x"74", x"74", x"74", x"75", x"74", x"73", x"73", x"73", x"72", x"71", x"73", x"74", x"74", x"72", 
        x"72", x"72", x"74", x"75", x"73", x"71", x"6f", x"6f", x"6f", x"72", x"73", x"74", x"72", x"74", x"76", 
        x"73", x"70", x"6f", x"70", x"73", x"72", x"6f", x"6e", x"6f", x"70", x"71", x"73", x"6f", x"70", x"73", 
        x"6f", x"6e", x"70", x"6f", x"72", x"71", x"73", x"70", x"75", x"71", x"6e", x"71", x"71", x"6e", x"6e", 
        x"70", x"74", x"74", x"72", x"72", x"6f", x"6f", x"71", x"70", x"70", x"6f", x"6e", x"6d", x"70", x"72", 
        x"71", x"72", x"72", x"71", x"71", x"72", x"72", x"6f", x"70", x"72", x"73", x"72", x"71", x"70", x"72", 
        x"72", x"71", x"71", x"71", x"71", x"71", x"70", x"6e", x"70", x"70", x"72", x"72", x"71", x"71", x"6d", 
        x"74", x"73", x"72", x"72", x"71", x"70", x"6e", x"6d", x"6d", x"6e", x"6f", x"6e", x"6c", x"70", x"71", 
        x"6f", x"70", x"70", x"6e", x"6b", x"6d", x"6f", x"6f", x"6e", x"6d", x"6e", x"6e", x"6d", x"6b", x"6c", 
        x"70", x"70", x"6f", x"71", x"71", x"6e", x"6f", x"6f", x"6f", x"6f", x"6e", x"6d", x"6d", x"6e", x"6e", 
        x"6e", x"6f", x"71", x"6f", x"6e", x"6e", x"71", x"6e", x"6c", x"6c", x"6f", x"73", x"72", x"72", x"73", 
        x"70", x"70", x"73", x"73", x"70", x"6c", x"6f", x"72", x"70", x"72", x"72", x"6e", x"70", x"6f", x"70", 
        x"70", x"72", x"73", x"73", x"74", x"72", x"70", x"70", x"72", x"70", x"6e", x"6f", x"70", x"70", x"72", 
        x"73", x"74", x"74", x"74", x"74", x"74", x"73", x"72", x"72", x"71", x"72", x"74", x"75", x"74", x"71", 
        x"71", x"75", x"75", x"71", x"73", x"73", x"72", x"71", x"72", x"73", x"72", x"75", x"77", x"74", x"71", 
        x"71", x"74", x"72", x"71", x"70", x"71", x"73", x"74", x"73", x"76", x"74", x"73", x"75", x"75", x"73", 
        x"74", x"76", x"77", x"74", x"75", x"77", x"77", x"76", x"75", x"75", x"74", x"74", x"76", x"73", x"6b", 
        x"86", x"d7", x"d4", x"d0", x"d1", x"d3", x"dc", x"d2", x"ce", x"cf", x"d0", x"ce", x"cd", x"cd", x"ce", 
        x"cf", x"cf", x"ce", x"ce", x"cf", x"d0", x"d0", x"cf", x"cf", x"cf", x"ce", x"d0", x"cf", x"cf", x"d1", 
        x"d0", x"cd", x"cc", x"ce", x"cf", x"ce", x"d0", x"d2", x"cf", x"d2", x"d1", x"cf", x"d4", x"d8", x"c8", 
        x"96", x"90", x"bb", x"d6", x"ce", x"cc", x"cb", x"d9", x"d5", x"d1", x"d0", x"d1", x"d1", x"d1", x"c8", 
        x"9d", x"62", x"5c", x"5d", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"8b", x"ed", x"fb", x"fa", x"fa", x"f9", x"f8", x"ba", x"65", 
        x"5d", x"61", x"5d", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", x"5e", 
        x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", 
        x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"60", x"86", x"dd", 
        x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ef", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ea", x"d5", x"c3", x"c8", x"da", x"e6", 
        x"d7", x"ab", x"81", x"6d", x"70", x"78", x"7e", x"82", x"80", x"7e", x"7f", x"7a", x"79", x"7c", x"7c", 
        x"7a", x"7d", x"7b", x"7c", x"7c", x"7e", x"7e", x"7d", x"7c", x"7c", x"7b", x"7b", x"7a", x"7a", x"7b", 
        x"7a", x"7c", x"7e", x"7e", x"7f", x"7f", x"7d", x"7c", x"7d", x"7e", x"7c", x"7a", x"7b", x"7c", x"7d", 
        x"7c", x"7b", x"7a", x"7a", x"7c", x"7a", x"79", x"79", x"7b", x"7c", x"7a", x"76", x"77", x"7a", x"7a", 
        x"7a", x"7a", x"7b", x"7c", x"7a", x"7c", x"79", x"79", x"79", x"7a", x"7b", x"7b", x"7d", x"7d", x"7c", 
        x"7b", x"7b", x"7c", x"7c", x"7c", x"7a", x"79", x"7b", x"79", x"77", x"79", x"79", x"79", x"79", x"79", 
        x"7a", x"79", x"78", x"79", x"7a", x"79", x"78", x"7a", x"7c", x"79", x"76", x"7c", x"7b", x"7c", x"79", 
        x"76", x"79", x"79", x"77", x"76", x"78", x"7a", x"7a", x"79", x"79", x"7a", x"79", x"78", x"78", x"79", 
        x"79", x"77", x"7a", x"7b", x"79", x"7a", x"7a", x"77", x"7b", x"7b", x"7b", x"79", x"7a", x"79", x"78", 
        x"79", x"7a", x"78", x"76", x"79", x"7b", x"7b", x"78", x"78", x"77", x"75", x"76", x"79", x"79", x"77", 
        x"75", x"75", x"76", x"76", x"75", x"7a", x"7a", x"78", x"78", x"78", x"78", x"78", x"79", x"78", x"77", 
        x"77", x"7a", x"77", x"77", x"7a", x"79", x"77", x"78", x"78", x"76", x"77", x"79", x"79", x"77", x"79", 
        x"79", x"76", x"76", x"79", x"78", x"77", x"78", x"79", x"77", x"75", x"76", x"79", x"7a", x"7a", x"79", 
        x"77", x"78", x"79", x"78", x"75", x"75", x"76", x"76", x"76", x"76", x"76", x"75", x"75", x"77", x"79", 
        x"76", x"74", x"73", x"73", x"74", x"76", x"77", x"76", x"74", x"73", x"73", x"71", x"72", x"74", x"75", 
        x"73", x"73", x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"72", x"71", x"72", x"75", 
        x"75", x"72", x"71", x"72", x"74", x"73", x"71", x"71", x"71", x"71", x"72", x"74", x"71", x"70", x"73", 
        x"74", x"75", x"75", x"74", x"72", x"70", x"71", x"73", x"74", x"73", x"76", x"73", x"73", x"75", x"73", 
        x"75", x"73", x"73", x"72", x"75", x"73", x"74", x"72", x"72", x"6f", x"70", x"71", x"6e", x"6e", x"71", 
        x"70", x"70", x"73", x"73", x"70", x"71", x"71", x"71", x"75", x"73", x"72", x"74", x"74", x"70", x"6d", 
        x"6d", x"72", x"70", x"6f", x"71", x"6d", x"6c", x"6c", x"6d", x"6f", x"71", x"71", x"70", x"71", x"71", 
        x"71", x"70", x"6e", x"6d", x"6e", x"70", x"72", x"6f", x"6f", x"70", x"72", x"72", x"72", x"72", x"70", 
        x"70", x"70", x"71", x"72", x"74", x"75", x"73", x"72", x"71", x"71", x"71", x"71", x"71", x"6f", x"6e", 
        x"71", x"70", x"6f", x"6f", x"70", x"70", x"70", x"6e", x"6e", x"6f", x"70", x"6e", x"6d", x"6f", x"70", 
        x"6e", x"6f", x"70", x"6e", x"6c", x"6e", x"6e", x"6d", x"6c", x"6d", x"6e", x"6f", x"6d", x"6c", x"6c", 
        x"6f", x"6f", x"6f", x"6f", x"6e", x"6c", x"6f", x"6f", x"6d", x"6c", x"6c", x"6d", x"6e", x"70", x"6e", 
        x"6c", x"6d", x"6f", x"72", x"72", x"70", x"71", x"70", x"6f", x"6e", x"6e", x"71", x"71", x"72", x"71", 
        x"6f", x"6e", x"70", x"71", x"71", x"72", x"72", x"74", x"71", x"71", x"73", x"70", x"6f", x"71", x"72", 
        x"71", x"6f", x"71", x"74", x"72", x"73", x"73", x"74", x"75", x"73", x"71", x"74", x"73", x"72", x"72", 
        x"72", x"73", x"73", x"72", x"72", x"72", x"71", x"72", x"72", x"71", x"71", x"71", x"73", x"73", x"72", 
        x"72", x"73", x"73", x"72", x"74", x"73", x"72", x"71", x"73", x"74", x"72", x"74", x"75", x"74", x"72", 
        x"73", x"75", x"72", x"73", x"74", x"76", x"76", x"76", x"75", x"76", x"75", x"73", x"75", x"75", x"73", 
        x"74", x"75", x"77", x"77", x"76", x"75", x"73", x"75", x"76", x"76", x"75", x"75", x"77", x"75", x"6d", 
        x"88", x"d7", x"d4", x"d0", x"d1", x"d3", x"dc", x"d2", x"ce", x"cf", x"cf", x"ce", x"ce", x"ce", x"cf", 
        x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"cf", x"ce", x"d0", x"cf", x"cf", x"cf", 
        x"ce", x"cf", x"d0", x"d2", x"cf", x"cf", x"d2", x"d0", x"d1", x"d0", x"d2", x"d6", x"ce", x"b7", x"9d", 
        x"a8", x"c7", x"cf", x"ca", x"cb", x"cf", x"cb", x"d8", x"d3", x"d0", x"cf", x"d0", x"cf", x"d1", x"c9", 
        x"9e", x"63", x"5d", x"5e", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5c", x"63", x"a6", x"f6", x"fb", x"fa", x"fb", x"fa", x"f9", x"b4", x"66", 
        x"5d", x"5f", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"60", x"83", x"db", 
        x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"f0", x"f1", x"eb", x"d9", x"cb", x"c8", 
        x"d4", x"da", x"d3", x"b9", x"95", x"7b", x"71", x"74", x"7e", x"80", x"7d", x"7e", x"7c", x"7d", x"7e", 
        x"7c", x"7d", x"7d", x"7e", x"7d", x"7d", x"7d", x"7e", x"7d", x"7c", x"7b", x"7a", x"7c", x"7d", x"7d", 
        x"7b", x"7b", x"7b", x"7b", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7c", x"7b", x"7c", x"7c", x"7c", 
        x"7c", x"7b", x"7a", x"7a", x"7d", x"7c", x"7a", x"7b", x"7c", x"7c", x"7c", x"7d", x"7b", x"77", x"77", 
        x"78", x"7a", x"7b", x"7a", x"7a", x"7d", x"7c", x"7b", x"7a", x"79", x"7b", x"7b", x"7a", x"7b", x"7c", 
        x"7b", x"7a", x"78", x"78", x"79", x"79", x"7a", x"7c", x"79", x"77", x"7a", x"7b", x"7b", x"7b", x"7a", 
        x"7b", x"7b", x"78", x"79", x"7c", x"7c", x"7a", x"7a", x"7b", x"78", x"76", x"79", x"79", x"7c", x"7b", 
        x"7a", x"79", x"78", x"77", x"78", x"7a", x"7b", x"7b", x"79", x"79", x"79", x"79", x"79", x"7a", x"7b", 
        x"79", x"78", x"7a", x"7a", x"79", x"7a", x"7a", x"78", x"79", x"78", x"77", x"77", x"79", x"79", x"7a", 
        x"79", x"7a", x"79", x"77", x"79", x"7a", x"7a", x"79", x"79", x"78", x"76", x"77", x"7a", x"7a", x"77", 
        x"74", x"76", x"78", x"77", x"77", x"7a", x"7b", x"7a", x"7a", x"7a", x"79", x"79", x"78", x"78", x"76", 
        x"76", x"78", x"77", x"78", x"7a", x"79", x"77", x"79", x"78", x"77", x"78", x"79", x"77", x"77", x"79", 
        x"79", x"76", x"76", x"78", x"78", x"75", x"76", x"78", x"77", x"74", x"74", x"76", x"79", x"78", x"75", 
        x"77", x"79", x"77", x"76", x"78", x"77", x"77", x"76", x"77", x"76", x"77", x"77", x"78", x"78", x"78", 
        x"76", x"75", x"75", x"75", x"74", x"75", x"76", x"75", x"74", x"74", x"74", x"73", x"74", x"75", x"75", 
        x"74", x"74", x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"74", x"76", x"75", x"73", 
        x"71", x"6f", x"71", x"74", x"75", x"74", x"72", x"72", x"71", x"70", x"73", x"74", x"70", x"6e", x"73", 
        x"74", x"76", x"72", x"71", x"73", x"73", x"73", x"72", x"70", x"73", x"75", x"72", x"73", x"73", x"73", 
        x"74", x"72", x"71", x"71", x"73", x"71", x"72", x"70", x"72", x"72", x"72", x"72", x"71", x"71", x"73", 
        x"72", x"70", x"72", x"72", x"70", x"72", x"73", x"73", x"72", x"71", x"71", x"72", x"73", x"72", x"71", 
        x"71", x"74", x"73", x"72", x"73", x"71", x"70", x"6f", x"6f", x"70", x"70", x"70", x"70", x"71", x"71", 
        x"70", x"70", x"71", x"70", x"70", x"70", x"71", x"71", x"71", x"71", x"71", x"73", x"74", x"75", x"72", 
        x"72", x"72", x"72", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"73", x"70", x"6f", 
        x"71", x"71", x"72", x"72", x"72", x"70", x"6e", x"6f", x"6f", x"6f", x"70", x"6e", x"6d", x"6e", x"6f", 
        x"6e", x"6f", x"6f", x"6f", x"6e", x"6f", x"6f", x"6d", x"6d", x"6e", x"6f", x"6e", x"6d", x"6b", x"6d", 
        x"6e", x"6d", x"6d", x"6e", x"6f", x"6e", x"6f", x"6f", x"70", x"70", x"6f", x"6e", x"6d", x"70", x"70", 
        x"6e", x"6e", x"70", x"72", x"72", x"70", x"70", x"71", x"73", x"71", x"6f", x"6f", x"71", x"72", x"71", 
        x"6f", x"6f", x"70", x"71", x"73", x"74", x"72", x"72", x"70", x"6f", x"70", x"71", x"71", x"70", x"70", 
        x"72", x"74", x"71", x"6f", x"6f", x"71", x"74", x"75", x"74", x"72", x"71", x"73", x"72", x"71", x"71", 
        x"72", x"73", x"72", x"71", x"71", x"71", x"72", x"73", x"73", x"73", x"72", x"70", x"72", x"73", x"73", 
        x"73", x"73", x"73", x"73", x"74", x"74", x"73", x"72", x"74", x"74", x"72", x"73", x"74", x"75", x"74", 
        x"74", x"75", x"72", x"72", x"74", x"74", x"74", x"74", x"75", x"76", x"75", x"74", x"75", x"75", x"74", 
        x"74", x"73", x"76", x"77", x"77", x"74", x"73", x"77", x"78", x"77", x"77", x"76", x"78", x"77", x"70", 
        x"8a", x"d8", x"d5", x"d0", x"d1", x"d2", x"db", x"d2", x"ce", x"cf", x"cf", x"ce", x"ce", x"ce", x"cf", 
        x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"cf", x"ce", x"d0", x"cf", x"cf", x"cf", 
        x"cf", x"d0", x"cd", x"cf", x"d0", x"cd", x"cf", x"d0", x"cf", x"d1", x"d8", x"c7", x"a2", x"a1", x"bc", 
        x"d4", x"d0", x"ca", x"ca", x"ca", x"cc", x"cb", x"d8", x"d4", x"cf", x"d0", x"d1", x"cf", x"d0", x"c8", 
        x"9e", x"64", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"65", x"b9", x"fa", x"fb", x"fb", x"fa", x"fb", x"f9", x"ae", x"66", 
        x"5d", x"5e", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"80", x"d8", 
        x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ec", x"ee", x"f2", x"f2", x"ed", x"de", 
        x"cb", x"c5", x"cd", x"de", x"dd", x"bf", x"95", x"7c", x"71", x"71", x"79", x"7d", x"7d", x"7f", x"7f", 
        x"7d", x"7c", x"79", x"7c", x"7e", x"7d", x"7d", x"7e", x"7e", x"7d", x"7b", x"7a", x"7b", x"7b", x"7c", 
        x"7b", x"7c", x"7d", x"7d", x"7e", x"7e", x"7e", x"7c", x"7b", x"7b", x"7a", x"7b", x"7b", x"7b", x"7b", 
        x"7b", x"7a", x"7a", x"7a", x"7b", x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", x"7d", x"7c", x"7a", x"7a", 
        x"7b", x"7a", x"78", x"7a", x"7a", x"7d", x"7c", x"7b", x"7b", x"7b", x"7c", x"7a", x"79", x"7a", x"7b", 
        x"7b", x"79", x"78", x"79", x"78", x"78", x"7a", x"7c", x"7c", x"7a", x"7a", x"7b", x"7c", x"7a", x"79", 
        x"7a", x"7b", x"78", x"7a", x"7c", x"7d", x"7b", x"7a", x"79", x"7c", x"7a", x"7a", x"78", x"79", x"7a", 
        x"7a", x"79", x"79", x"79", x"7a", x"7b", x"7b", x"7a", x"7a", x"79", x"78", x"79", x"7a", x"7c", x"7c", 
        x"7a", x"7a", x"7c", x"79", x"79", x"7a", x"78", x"78", x"79", x"78", x"78", x"78", x"78", x"77", x"78", 
        x"79", x"7a", x"79", x"78", x"79", x"79", x"78", x"79", x"7a", x"79", x"78", x"79", x"7a", x"7b", x"7a", 
        x"78", x"77", x"77", x"77", x"76", x"79", x"7c", x"7c", x"7b", x"7b", x"7a", x"78", x"78", x"78", x"78", 
        x"78", x"78", x"78", x"79", x"79", x"77", x"78", x"79", x"79", x"78", x"79", x"78", x"76", x"78", x"79", 
        x"78", x"76", x"75", x"78", x"79", x"77", x"77", x"79", x"78", x"76", x"75", x"75", x"77", x"76", x"76", 
        x"77", x"78", x"78", x"77", x"78", x"78", x"77", x"75", x"74", x"74", x"76", x"76", x"78", x"77", x"77", 
        x"77", x"77", x"77", x"75", x"72", x"73", x"75", x"76", x"76", x"77", x"78", x"76", x"76", x"76", x"75", 
        x"74", x"74", x"75", x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"72", x"73", x"74", x"75", x"73", 
        x"72", x"72", x"73", x"74", x"74", x"73", x"73", x"75", x"74", x"72", x"73", x"75", x"72", x"71", x"73", 
        x"73", x"73", x"70", x"70", x"72", x"73", x"72", x"71", x"6f", x"71", x"72", x"72", x"74", x"72", x"72", 
        x"73", x"71", x"72", x"72", x"73", x"72", x"73", x"71", x"73", x"74", x"73", x"70", x"73", x"73", x"72", 
        x"73", x"73", x"73", x"72", x"70", x"70", x"71", x"71", x"71", x"71", x"71", x"71", x"72", x"73", x"73", 
        x"73", x"74", x"74", x"74", x"75", x"74", x"73", x"72", x"72", x"71", x"70", x"6f", x"70", x"73", x"73", 
        x"72", x"71", x"72", x"72", x"72", x"71", x"71", x"72", x"73", x"74", x"74", x"73", x"72", x"72", x"74", 
        x"74", x"73", x"73", x"72", x"72", x"72", x"72", x"73", x"73", x"72", x"72", x"71", x"71", x"72", x"72", 
        x"6f", x"71", x"74", x"76", x"75", x"74", x"71", x"71", x"6f", x"6f", x"70", x"6f", x"6d", x"6e", x"6f", 
        x"6f", x"6f", x"6f", x"6f", x"6f", x"6f", x"6e", x"6d", x"6f", x"70", x"70", x"70", x"70", x"6f", x"6f", 
        x"70", x"70", x"70", x"6e", x"6c", x"6c", x"70", x"70", x"6f", x"6f", x"6f", x"6f", x"6f", x"70", x"71", 
        x"72", x"71", x"71", x"70", x"6f", x"71", x"70", x"71", x"73", x"72", x"6f", x"6e", x"70", x"70", x"70", 
        x"71", x"71", x"72", x"72", x"73", x"72", x"6f", x"70", x"70", x"6e", x"6e", x"71", x"73", x"72", x"70", 
        x"6f", x"6f", x"70", x"70", x"6f", x"71", x"74", x"73", x"71", x"6f", x"70", x"71", x"71", x"71", x"72", 
        x"74", x"73", x"72", x"72", x"73", x"74", x"75", x"75", x"76", x"77", x"75", x"72", x"72", x"73", x"73", 
        x"74", x"74", x"73", x"73", x"75", x"76", x"75", x"74", x"74", x"74", x"74", x"74", x"74", x"75", x"75", 
        x"74", x"74", x"73", x"74", x"75", x"74", x"73", x"74", x"76", x"76", x"76", x"75", x"74", x"74", x"75", 
        x"75", x"75", x"76", x"76", x"76", x"74", x"73", x"75", x"76", x"77", x"78", x"76", x"78", x"77", x"70", 
        x"89", x"d7", x"d5", x"d1", x"d1", x"d2", x"db", x"d2", x"ce", x"ce", x"cf", x"ce", x"ce", x"ce", x"d0", 
        x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"cf", x"ce", x"d0", x"cf", x"cf", x"cc", 
        x"cd", x"d2", x"ce", x"ce", x"d0", x"ce", x"cb", x"cc", x"d4", x"cd", x"a7", x"98", x"b4", x"ca", x"d1", 
        x"ca", x"cd", x"cd", x"d0", x"d2", x"cd", x"cb", x"da", x"d6", x"d0", x"d1", x"d2", x"d0", x"d0", x"c8", 
        x"9f", x"65", x"5f", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"62", x"be", x"f9", x"fb", x"fc", x"fb", x"fb", x"f7", x"aa", x"65", 
        x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5f", x"79", x"d1", 
        x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", x"f1", 
        x"f2", x"e5", x"d3", x"cb", x"cf", x"d9", x"e2", x"d0", x"aa", x"84", x"6f", x"6c", x"78", x"7d", x"81", 
        x"7f", x"7d", x"7d", x"80", x"7f", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7d", x"7d", 
        x"7c", x"7c", x"7d", x"7d", x"7e", x"7f", x"7e", x"7d", x"7b", x"7a", x"79", x"7a", x"7c", x"7b", x"7b", 
        x"7b", x"7b", x"7c", x"7b", x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7a", x"7c", x"7c", x"7b", x"7b", 
        x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7a", x"79", x"7b", x"7e", x"7d", x"7c", x"7c", x"7b", x"7a", 
        x"7a", x"7a", x"7a", x"7a", x"7a", x"7b", x"7d", x"7d", x"7c", x"7a", x"7a", x"7b", x"7b", x"7a", x"78", 
        x"79", x"7a", x"79", x"7a", x"7b", x"7b", x"7a", x"79", x"79", x"7d", x"7c", x"7a", x"7a", x"79", x"7a", 
        x"7a", x"79", x"79", x"79", x"7a", x"7a", x"7c", x"7d", x"7c", x"7a", x"78", x"79", x"7a", x"7c", x"7c", 
        x"79", x"7b", x"7c", x"78", x"79", x"7b", x"79", x"7a", x"79", x"79", x"7b", x"7c", x"79", x"77", x"78", 
        x"79", x"7a", x"7a", x"7a", x"79", x"78", x"78", x"7a", x"7b", x"7a", x"7a", x"7a", x"7a", x"7b", x"79", 
        x"76", x"77", x"7a", x"7b", x"79", x"7a", x"7b", x"79", x"79", x"79", x"79", x"78", x"78", x"79", x"7a", 
        x"79", x"79", x"7a", x"7b", x"79", x"77", x"78", x"7a", x"79", x"79", x"79", x"78", x"76", x"78", x"79", 
        x"78", x"77", x"77", x"78", x"7a", x"7a", x"7a", x"7b", x"7b", x"78", x"77", x"77", x"75", x"77", x"79", 
        x"77", x"78", x"7b", x"7a", x"79", x"79", x"79", x"78", x"77", x"76", x"76", x"76", x"76", x"76", x"76", 
        x"77", x"78", x"77", x"74", x"74", x"74", x"75", x"75", x"75", x"74", x"74", x"76", x"77", x"76", x"75", 
        x"74", x"74", x"75", x"76", x"75", x"75", x"75", x"75", x"75", x"75", x"74", x"73", x"73", x"73", x"74", 
        x"74", x"74", x"74", x"75", x"75", x"74", x"73", x"75", x"74", x"72", x"71", x"73", x"70", x"70", x"74", 
        x"74", x"76", x"72", x"71", x"71", x"70", x"70", x"71", x"71", x"72", x"71", x"71", x"74", x"71", x"72", 
        x"73", x"72", x"74", x"74", x"74", x"74", x"74", x"74", x"74", x"73", x"72", x"6f", x"72", x"72", x"6f", 
        x"72", x"72", x"72", x"71", x"71", x"71", x"73", x"73", x"70", x"72", x"72", x"71", x"72", x"72", x"70", 
        x"71", x"73", x"74", x"74", x"74", x"74", x"73", x"73", x"73", x"72", x"72", x"72", x"74", x"75", x"75", 
        x"73", x"73", x"72", x"72", x"73", x"73", x"73", x"75", x"74", x"73", x"72", x"71", x"71", x"71", x"75", 
        x"74", x"73", x"72", x"72", x"72", x"73", x"73", x"74", x"74", x"74", x"73", x"72", x"71", x"70", x"70", 
        x"6e", x"70", x"71", x"72", x"72", x"72", x"73", x"71", x"6f", x"6e", x"70", x"70", x"6e", x"6f", x"70", 
        x"70", x"6f", x"6f", x"6f", x"70", x"6f", x"6e", x"6f", x"70", x"71", x"70", x"71", x"71", x"70", x"6d", 
        x"6f", x"72", x"73", x"71", x"6e", x"6d", x"6f", x"6e", x"6d", x"6d", x"6d", x"6e", x"6f", x"6f", x"70", 
        x"71", x"71", x"71", x"71", x"72", x"73", x"71", x"71", x"71", x"72", x"70", x"6f", x"70", x"6d", x"6e", 
        x"71", x"72", x"71", x"71", x"71", x"71", x"71", x"72", x"73", x"72", x"70", x"73", x"72", x"73", x"72", 
        x"70", x"6f", x"70", x"72", x"73", x"75", x"75", x"73", x"70", x"70", x"71", x"70", x"71", x"72", x"73", 
        x"74", x"73", x"72", x"71", x"71", x"72", x"73", x"74", x"74", x"75", x"74", x"72", x"72", x"72", x"72", 
        x"72", x"73", x"73", x"73", x"75", x"76", x"76", x"75", x"74", x"74", x"75", x"75", x"75", x"75", x"75", 
        x"74", x"73", x"73", x"74", x"75", x"76", x"75", x"74", x"75", x"76", x"77", x"76", x"74", x"74", x"75", 
        x"76", x"77", x"78", x"75", x"75", x"76", x"75", x"75", x"74", x"76", x"78", x"76", x"77", x"77", x"70", 
        x"88", x"d6", x"d5", x"d2", x"d2", x"d3", x"dc", x"d4", x"cd", x"cd", x"cf", x"ce", x"ce", x"ce", x"d0", 
        x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"cf", x"ce", x"d0", x"cf", x"cf", x"cc", 
        x"ca", x"ce", x"ce", x"cf", x"d0", x"d0", x"cf", x"cc", x"b7", x"9e", x"a5", x"c0", x"cd", x"c8", x"cc", 
        x"ca", x"ca", x"cf", x"ce", x"ce", x"d0", x"cb", x"d9", x"d7", x"ce", x"cf", x"d1", x"cf", x"d0", x"c8", 
        x"9f", x"65", x"5f", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"63", x"be", x"f8", x"fa", x"fc", x"fb", x"fa", x"f7", x"b2", x"66", 
        x"5c", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"74", x"cb", 
        x"ed", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", 
        x"ef", x"ed", x"ef", x"e7", x"db", x"d5", x"d0", x"d3", x"d7", x"cd", x"b1", x"90", x"7b", x"71", x"76", 
        x"7c", x"7f", x"7e", x"7e", x"7f", x"7e", x"7e", x"7d", x"7d", x"7d", x"7e", x"7e", x"7d", x"7c", x"7d", 
        x"7c", x"7c", x"7d", x"7d", x"7d", x"7d", x"7c", x"7b", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7b", 
        x"7b", x"7c", x"7d", x"7c", x"7b", x"7c", x"7c", x"7c", x"7b", x"7c", x"7c", x"7b", x"7c", x"7b", x"7a", 
        x"79", x"7c", x"7e", x"7b", x"7b", x"7b", x"7b", x"7a", x"7b", x"7e", x"7d", x"7e", x"7e", x"7d", x"7a", 
        x"7a", x"7c", x"7c", x"7a", x"7a", x"7c", x"7d", x"7c", x"79", x"79", x"7c", x"7c", x"7b", x"7b", x"7a", 
        x"7a", x"7a", x"7b", x"7a", x"79", x"79", x"7a", x"79", x"7a", x"79", x"7b", x"7a", x"7b", x"7b", x"7d", 
        x"7d", x"7a", x"7a", x"79", x"79", x"79", x"7b", x"7d", x"7d", x"7b", x"7a", x"79", x"7a", x"7a", x"7a", 
        x"79", x"7b", x"7c", x"78", x"79", x"7b", x"7b", x"7c", x"7d", x"7a", x"7b", x"7c", x"79", x"78", x"7b", 
        x"7a", x"79", x"79", x"7a", x"79", x"78", x"79", x"7b", x"7b", x"7b", x"7b", x"7b", x"7a", x"7b", x"7a", 
        x"79", x"7a", x"7c", x"7d", x"7a", x"78", x"78", x"77", x"78", x"78", x"79", x"79", x"79", x"78", x"77", 
        x"78", x"79", x"7b", x"7c", x"7a", x"79", x"78", x"7a", x"7a", x"78", x"78", x"79", x"78", x"78", x"78", 
        x"79", x"79", x"78", x"78", x"79", x"7a", x"79", x"7a", x"7a", x"79", x"78", x"77", x"77", x"77", x"78", 
        x"79", x"7a", x"7a", x"7b", x"7b", x"7a", x"7a", x"7a", x"79", x"78", x"76", x"75", x"77", x"75", x"75", 
        x"75", x"76", x"76", x"75", x"75", x"74", x"75", x"75", x"76", x"75", x"75", x"75", x"76", x"76", x"75", 
        x"74", x"74", x"75", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"75", x"75", x"75", x"75", x"73", 
        x"72", x"72", x"74", x"75", x"76", x"74", x"73", x"75", x"74", x"72", x"73", x"75", x"71", x"70", x"73", 
        x"73", x"74", x"73", x"72", x"72", x"71", x"71", x"72", x"72", x"72", x"72", x"72", x"74", x"72", x"72", 
        x"73", x"72", x"73", x"73", x"72", x"73", x"72", x"73", x"74", x"76", x"74", x"72", x"73", x"73", x"72", 
        x"73", x"72", x"71", x"71", x"73", x"73", x"73", x"73", x"6f", x"72", x"73", x"72", x"73", x"74", x"71", 
        x"72", x"71", x"73", x"74", x"73", x"73", x"72", x"72", x"72", x"73", x"74", x"75", x"75", x"75", x"73", 
        x"72", x"73", x"74", x"72", x"72", x"72", x"73", x"73", x"72", x"71", x"70", x"71", x"72", x"73", x"74", 
        x"74", x"73", x"72", x"73", x"74", x"74", x"74", x"74", x"75", x"75", x"74", x"73", x"72", x"71", x"71", 
        x"71", x"72", x"71", x"70", x"6f", x"6f", x"72", x"71", x"6e", x"6e", x"71", x"71", x"70", x"70", x"70", 
        x"70", x"6f", x"6e", x"70", x"71", x"70", x"70", x"73", x"72", x"71", x"6f", x"6f", x"71", x"72", x"71", 
        x"70", x"71", x"71", x"6f", x"6e", x"6f", x"6d", x"6e", x"6f", x"70", x"6f", x"6f", x"6e", x"70", x"70", 
        x"71", x"70", x"70", x"72", x"75", x"74", x"71", x"72", x"71", x"72", x"73", x"71", x"72", x"70", x"6f", 
        x"71", x"71", x"70", x"70", x"72", x"72", x"73", x"72", x"75", x"75", x"72", x"74", x"72", x"71", x"72", 
        x"75", x"75", x"71", x"6e", x"74", x"76", x"75", x"73", x"72", x"72", x"73", x"6f", x"70", x"72", x"73", 
        x"72", x"74", x"74", x"72", x"71", x"72", x"72", x"73", x"74", x"74", x"73", x"72", x"74", x"73", x"71", 
        x"70", x"71", x"73", x"74", x"74", x"75", x"74", x"74", x"74", x"74", x"75", x"75", x"76", x"76", x"75", 
        x"74", x"74", x"72", x"73", x"75", x"76", x"75", x"74", x"72", x"74", x"77", x"78", x"74", x"74", x"75", 
        x"76", x"76", x"77", x"74", x"75", x"77", x"76", x"76", x"76", x"77", x"79", x"76", x"77", x"77", x"70", 
        x"87", x"d5", x"d5", x"d2", x"d2", x"d3", x"dd", x"d5", x"cd", x"cd", x"cf", x"ce", x"ce", x"cf", x"d0", 
        x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"cf", x"ce", x"d0", x"cf", x"cf", x"ce", 
        x"cb", x"cf", x"cf", x"cb", x"d1", x"d3", x"c2", x"a0", x"9a", x"bb", x"ce", x"ce", x"cc", x"c8", x"ca", 
        x"cb", x"ce", x"ce", x"ce", x"cb", x"cb", x"c7", x"d8", x"d8", x"cd", x"ce", x"d0", x"cf", x"d0", x"c8", 
        x"9f", x"65", x"5f", x"5f", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"65", x"b9", x"f7", x"f9", x"fc", x"fb", x"f9", x"f7", x"c0", x"6a", 
        x"5b", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"6f", x"c6", 
        x"ed", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"f1", x"ec", x"eb", x"ee", x"f0", x"ee", x"ef", 
        x"ef", x"ec", x"ee", x"f1", x"f0", x"ec", x"e0", x"d0", x"c7", x"c7", x"d9", x"db", x"c4", x"94", x"75", 
        x"68", x"79", x"81", x"7f", x"79", x"7d", x"7e", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", x"7e", x"7d", 
        x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7d", x"7f", x"7e", x"7d", x"7d", x"7c", x"7c", 
        x"7c", x"7d", x"7e", x"7e", x"7d", x"7e", x"7d", x"7c", x"7c", x"7d", x"7e", x"7b", x"7c", x"7e", x"7e", 
        x"7d", x"7d", x"7d", x"78", x"7a", x"7b", x"7d", x"7c", x"7c", x"7d", x"7c", x"7c", x"7c", x"7c", x"7b", 
        x"7b", x"7d", x"7e", x"7c", x"79", x"79", x"7a", x"79", x"79", x"7b", x"7e", x"7d", x"7b", x"7c", x"7c", 
        x"7b", x"7a", x"7d", x"7c", x"7a", x"79", x"7a", x"7b", x"7b", x"79", x"7b", x"79", x"7c", x"7c", x"7e", 
        x"7e", x"7c", x"7c", x"7b", x"79", x"78", x"78", x"7a", x"7b", x"7b", x"7a", x"7a", x"79", x"79", x"79", 
        x"79", x"7b", x"7b", x"79", x"78", x"7b", x"7c", x"7c", x"80", x"7b", x"7a", x"7b", x"77", x"78", x"7c", 
        x"7a", x"78", x"77", x"79", x"78", x"78", x"7a", x"7c", x"7b", x"7b", x"7c", x"7b", x"79", x"7a", x"7c", 
        x"7a", x"78", x"79", x"7a", x"7a", x"7c", x"7a", x"77", x"77", x"78", x"79", x"79", x"7a", x"78", x"76", 
        x"79", x"79", x"7c", x"7c", x"7a", x"7b", x"78", x"7b", x"7b", x"77", x"77", x"79", x"7a", x"78", x"78", 
        x"7a", x"7b", x"7a", x"77", x"79", x"79", x"79", x"79", x"79", x"79", x"78", x"79", x"79", x"77", x"78", 
        x"7a", x"7a", x"78", x"7a", x"7c", x"79", x"79", x"78", x"77", x"76", x"75", x"75", x"78", x"77", x"75", 
        x"73", x"73", x"76", x"77", x"78", x"77", x"77", x"77", x"77", x"76", x"74", x"73", x"73", x"75", x"75", 
        x"74", x"74", x"74", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"75", x"76", x"76", x"75", x"73", 
        x"72", x"74", x"74", x"73", x"75", x"74", x"74", x"75", x"76", x"74", x"70", x"73", x"72", x"73", x"76", 
        x"74", x"73", x"73", x"72", x"73", x"73", x"73", x"73", x"72", x"73", x"74", x"73", x"73", x"73", x"73", 
        x"74", x"73", x"72", x"73", x"71", x"72", x"71", x"73", x"74", x"76", x"75", x"74", x"73", x"72", x"73", 
        x"74", x"75", x"72", x"72", x"74", x"73", x"71", x"71", x"70", x"72", x"72", x"71", x"75", x"77", x"73", 
        x"73", x"71", x"74", x"74", x"72", x"73", x"72", x"71", x"71", x"71", x"72", x"73", x"73", x"72", x"70", 
        x"71", x"73", x"74", x"71", x"70", x"71", x"73", x"71", x"71", x"73", x"74", x"74", x"73", x"73", x"73", 
        x"74", x"74", x"74", x"74", x"73", x"73", x"72", x"73", x"74", x"74", x"73", x"72", x"70", x"72", x"74", 
        x"71", x"73", x"73", x"72", x"72", x"72", x"74", x"71", x"6e", x"6d", x"70", x"71", x"70", x"71", x"70", 
        x"6f", x"6f", x"6e", x"70", x"73", x"71", x"70", x"72", x"71", x"70", x"6e", x"6e", x"71", x"72", x"6f", 
        x"6e", x"70", x"72", x"70", x"6f", x"71", x"72", x"72", x"72", x"71", x"72", x"72", x"72", x"71", x"72", 
        x"72", x"71", x"70", x"71", x"73", x"72", x"70", x"73", x"71", x"73", x"74", x"71", x"76", x"77", x"74", 
        x"74", x"73", x"71", x"73", x"73", x"72", x"74", x"70", x"72", x"73", x"70", x"71", x"73", x"74", x"73", 
        x"72", x"72", x"72", x"73", x"73", x"73", x"73", x"72", x"71", x"72", x"73", x"72", x"73", x"73", x"71", 
        x"70", x"71", x"74", x"74", x"73", x"74", x"74", x"74", x"75", x"75", x"74", x"74", x"77", x"77", x"75", 
        x"72", x"72", x"73", x"75", x"74", x"73", x"72", x"73", x"75", x"75", x"74", x"75", x"76", x"76", x"75", 
        x"75", x"76", x"76", x"76", x"76", x"77", x"77", x"77", x"75", x"75", x"77", x"78", x"75", x"74", x"75", 
        x"76", x"77", x"78", x"77", x"76", x"77", x"75", x"77", x"77", x"79", x"7a", x"77", x"77", x"78", x"71", 
        x"87", x"d4", x"d5", x"d2", x"d2", x"d4", x"de", x"d6", x"cd", x"cd", x"cf", x"cf", x"cf", x"cf", x"d0", 
        x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"cf", x"d0", x"cf", x"ce", x"d0", x"cf", x"cf", x"cf", 
        x"cd", x"cd", x"ce", x"d2", x"d1", x"b4", x"92", x"ad", x"ca", x"d3", x"ce", x"cc", x"cb", x"cb", x"cc", 
        x"ce", x"ce", x"cd", x"cc", x"cd", x"cc", x"c8", x"da", x"db", x"cf", x"ce", x"d1", x"d1", x"d1", x"c9", 
        x"a0", x"66", x"5f", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"63", x"ae", x"f4", x"f8", x"fc", x"fa", x"f8", x"f8", x"d0", x"70", 
        x"5a", x"5c", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5c", x"5d", x"6d", x"c4", 
        x"ed", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ee", x"ed", x"ed", x"ef", x"f0", x"ef", x"ee", 
        x"ef", x"f1", x"ee", x"ee", x"f0", x"ee", x"ee", x"ee", x"e4", x"d5", x"c8", x"ca", x"d7", x"df", x"ce", 
        x"ac", x"84", x"71", x"74", x"7b", x"7c", x"7f", x"80", x"80", x"80", x"80", x"7f", x"7c", x"7b", x"7c", 
        x"7d", x"7d", x"7e", x"7f", x"7f", x"7d", x"7c", x"7c", x"7e", x"80", x"7e", x"7c", x"7d", x"7d", x"7d", 
        x"7d", x"7e", x"7e", x"7e", x"7d", x"7e", x"7d", x"7b", x"7b", x"7d", x"7e", x"7d", x"7c", x"7d", x"7f", 
        x"7f", x"7d", x"7b", x"77", x"7a", x"7a", x"7e", x"7c", x"7c", x"7c", x"7b", x"7b", x"79", x"79", x"7b", 
        x"7c", x"7c", x"7d", x"7b", x"7a", x"7c", x"7e", x"7b", x"7a", x"7c", x"7d", x"7b", x"79", x"7b", x"7c", 
        x"7a", x"79", x"7e", x"7d", x"7c", x"7b", x"7c", x"7d", x"7c", x"7a", x"7c", x"79", x"7c", x"7b", x"7d", 
        x"7f", x"7a", x"7b", x"7b", x"7b", x"79", x"79", x"7a", x"7a", x"7b", x"7b", x"79", x"78", x"78", x"78", 
        x"79", x"7a", x"7b", x"7b", x"78", x"7b", x"7d", x"7a", x"7c", x"78", x"78", x"7b", x"78", x"79", x"7d", 
        x"7b", x"78", x"77", x"79", x"78", x"79", x"7c", x"7c", x"7a", x"7a", x"7c", x"7b", x"79", x"79", x"7d", 
        x"7c", x"79", x"79", x"7a", x"7a", x"7b", x"7b", x"79", x"79", x"79", x"7a", x"7b", x"7b", x"7a", x"79", 
        x"7d", x"7b", x"7c", x"7a", x"77", x"79", x"77", x"7b", x"7a", x"77", x"76", x"79", x"7c", x"79", x"78", 
        x"7a", x"7c", x"7a", x"77", x"78", x"7b", x"7b", x"7b", x"7a", x"7b", x"7c", x"7c", x"79", x"78", x"79", 
        x"78", x"77", x"78", x"7a", x"7b", x"7c", x"7a", x"79", x"77", x"77", x"77", x"77", x"78", x"79", x"78", 
        x"76", x"75", x"75", x"76", x"76", x"75", x"76", x"77", x"77", x"77", x"75", x"72", x"72", x"74", x"75", 
        x"74", x"74", x"74", x"75", x"75", x"75", x"76", x"76", x"76", x"76", x"76", x"76", x"74", x"73", x"74", 
        x"75", x"75", x"73", x"74", x"76", x"75", x"73", x"74", x"75", x"74", x"72", x"75", x"72", x"72", x"75", 
        x"74", x"74", x"75", x"74", x"73", x"73", x"73", x"74", x"74", x"73", x"76", x"73", x"72", x"74", x"73", 
        x"74", x"75", x"74", x"75", x"72", x"74", x"73", x"75", x"75", x"74", x"74", x"75", x"70", x"6f", x"71", 
        x"72", x"73", x"71", x"72", x"75", x"74", x"72", x"73", x"74", x"74", x"72", x"71", x"75", x"77", x"73", 
        x"74", x"73", x"75", x"76", x"73", x"73", x"72", x"72", x"71", x"70", x"70", x"71", x"70", x"6f", x"6f", 
        x"72", x"73", x"72", x"6f", x"6e", x"72", x"76", x"75", x"74", x"74", x"74", x"73", x"73", x"73", x"72", 
        x"74", x"75", x"76", x"75", x"72", x"70", x"72", x"74", x"75", x"76", x"75", x"73", x"72", x"71", x"71", 
        x"73", x"73", x"70", x"70", x"73", x"71", x"72", x"72", x"70", x"6f", x"70", x"71", x"71", x"70", x"72", 
        x"74", x"73", x"71", x"70", x"72", x"70", x"6f", x"71", x"71", x"71", x"71", x"71", x"71", x"72", x"73", 
        x"71", x"71", x"71", x"72", x"72", x"72", x"70", x"72", x"73", x"70", x"70", x"70", x"6f", x"6f", x"70", 
        x"70", x"71", x"72", x"72", x"71", x"70", x"71", x"74", x"73", x"71", x"72", x"73", x"75", x"74", x"71", 
        x"72", x"71", x"70", x"71", x"73", x"73", x"72", x"70", x"70", x"70", x"6f", x"6e", x"70", x"75", x"73", 
        x"73", x"76", x"70", x"74", x"72", x"73", x"75", x"72", x"6f", x"73", x"72", x"72", x"74", x"74", x"73", 
        x"73", x"74", x"75", x"75", x"75", x"74", x"74", x"73", x"73", x"74", x"73", x"73", x"74", x"75", x"74", 
        x"74", x"74", x"74", x"73", x"74", x"73", x"73", x"75", x"76", x"75", x"78", x"76", x"76", x"75", x"73", 
        x"75", x"72", x"72", x"75", x"76", x"74", x"75", x"76", x"75", x"77", x"77", x"76", x"76", x"74", x"74", 
        x"79", x"79", x"78", x"75", x"74", x"77", x"77", x"76", x"78", x"77", x"79", x"76", x"78", x"7b", x"71", 
        x"87", x"d4", x"d6", x"d3", x"d3", x"d3", x"dc", x"d6", x"cb", x"cc", x"cd", x"cd", x"cf", x"d1", x"d0", 
        x"cf", x"cf", x"ce", x"ce", x"ce", x"cf", x"cf", x"d0", x"d0", x"cd", x"ce", x"d2", x"ce", x"ce", x"d1", 
        x"d1", x"d2", x"d5", x"c2", x"98", x"99", x"c6", x"cf", x"d2", x"d0", x"cd", x"cd", x"cd", x"cc", x"cd", 
        x"ce", x"ce", x"cd", x"cd", x"ce", x"ce", x"cb", x"d9", x"da", x"d0", x"cf", x"d2", x"d3", x"d2", x"cc", 
        x"a3", x"68", x"61", x"5e", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"61", x"a4", x"e3", x"ed", x"fa", x"fb", x"fa", x"f9", x"e0", x"81", 
        x"5f", x"61", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5c", x"5c", x"6c", x"c6", 
        x"eb", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ef", x"ef", x"ee", x"f0", x"f0", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ec", x"ec", x"ed", x"ee", x"ee", x"ef", x"ef", x"ee", 
        x"ef", x"ef", x"f1", x"f0", x"ee", x"ec", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ed", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"ee", x"ed", x"e8", x"dc", x"ce", x"cb", x"d5", 
        x"de", x"d7", x"b7", x"90", x"74", x"72", x"7a", x"7e", x"7e", x"7f", x"7f", x"81", x"7d", x"7d", x"7f", 
        x"7e", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", x"80", x"83", x"82", x"7e", x"7b", x"7c", x"7d", 
        x"7e", x"7d", x"7c", x"7c", x"7d", x"7d", x"7f", x"81", x"7f", x"7e", x"7e", x"7c", x"7a", x"7b", x"7d", 
        x"7d", x"7c", x"7c", x"7a", x"7b", x"7d", x"7e", x"7d", x"7d", x"7d", x"7d", x"7c", x"7b", x"7b", x"7a", 
        x"7a", x"7a", x"7c", x"7e", x"7c", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7c", 
        x"7c", x"7c", x"7d", x"7b", x"7b", x"7c", x"7c", x"7b", x"7a", x"7b", x"7c", x"7a", x"7a", x"7a", x"7b", 
        x"7b", x"7a", x"7a", x"7b", x"7b", x"7c", x"7b", x"7c", x"7a", x"7b", x"7b", x"7a", x"7b", x"7a", x"7a", 
        x"7c", x"7a", x"7c", x"7b", x"7a", x"7c", x"7c", x"7a", x"79", x"7a", x"79", x"78", x"79", x"7a", x"7a", 
        x"7b", x"7a", x"79", x"79", x"7a", x"7b", x"7c", x"79", x"79", x"79", x"78", x"7a", x"7c", x"7c", x"7b", 
        x"7a", x"79", x"78", x"79", x"7b", x"7b", x"7a", x"79", x"7a", x"7a", x"7b", x"7a", x"7a", x"7a", x"7c", 
        x"7b", x"7a", x"79", x"78", x"79", x"7a", x"7b", x"7a", x"78", x"77", x"78", x"7a", x"7b", x"7a", x"79", 
        x"7a", x"7a", x"78", x"77", x"7a", x"78", x"78", x"7a", x"7b", x"7c", x"7b", x"7a", x"79", x"79", x"79", 
        x"79", x"79", x"79", x"79", x"79", x"7a", x"79", x"78", x"79", x"79", x"77", x"77", x"78", x"77", x"77", 
        x"77", x"77", x"77", x"76", x"76", x"72", x"75", x"76", x"74", x"76", x"77", x"76", x"75", x"74", x"75", 
        x"75", x"74", x"73", x"73", x"73", x"72", x"75", x"76", x"76", x"76", x"75", x"76", x"76", x"76", x"77", 
        x"77", x"77", x"77", x"77", x"74", x"74", x"72", x"74", x"76", x"74", x"75", x"76", x"74", x"72", x"75", 
        x"74", x"72", x"75", x"73", x"71", x"72", x"74", x"75", x"73", x"70", x"74", x"74", x"71", x"73", x"73", 
        x"74", x"72", x"74", x"77", x"73", x"72", x"76", x"75", x"73", x"75", x"74", x"76", x"74", x"71", x"71", 
        x"73", x"76", x"75", x"73", x"75", x"75", x"72", x"73", x"74", x"72", x"71", x"74", x"76", x"76", x"73", 
        x"73", x"70", x"72", x"73", x"73", x"73", x"71", x"73", x"72", x"70", x"72", x"74", x"73", x"72", x"72", 
        x"73", x"71", x"75", x"76", x"71", x"74", x"77", x"75", x"74", x"75", x"75", x"73", x"72", x"72", x"70", 
        x"70", x"71", x"74", x"75", x"74", x"73", x"74", x"72", x"72", x"75", x"76", x"74", x"73", x"75", x"73", 
        x"72", x"73", x"71", x"72", x"74", x"72", x"73", x"72", x"72", x"72", x"72", x"70", x"6f", x"6e", x"71", 
        x"73", x"73", x"71", x"70", x"72", x"72", x"70", x"71", x"71", x"71", x"70", x"6f", x"6e", x"6f", x"71", 
        x"70", x"70", x"70", x"73", x"74", x"74", x"70", x"72", x"73", x"70", x"70", x"70", x"6f", x"71", x"71", 
        x"71", x"71", x"72", x"71", x"6f", x"70", x"73", x"74", x"73", x"71", x"72", x"75", x"74", x"70", x"6f", 
        x"71", x"72", x"71", x"72", x"74", x"72", x"71", x"6f", x"70", x"71", x"72", x"71", x"72", x"74", x"70", 
        x"71", x"75", x"71", x"76", x"72", x"71", x"73", x"72", x"71", x"74", x"73", x"74", x"75", x"74", x"74", 
        x"75", x"76", x"77", x"73", x"72", x"73", x"74", x"74", x"75", x"77", x"75", x"73", x"75", x"75", x"73", 
        x"72", x"73", x"73", x"71", x"73", x"72", x"71", x"73", x"74", x"73", x"74", x"73", x"76", x"76", x"74", 
        x"74", x"71", x"72", x"74", x"74", x"72", x"73", x"75", x"75", x"77", x"75", x"74", x"75", x"75", x"75", 
        x"78", x"78", x"77", x"76", x"75", x"77", x"77", x"76", x"78", x"76", x"78", x"76", x"78", x"7b", x"72", 
        x"88", x"d3", x"d5", x"d3", x"d3", x"d2", x"db", x"d5", x"cb", x"cc", x"cd", x"cd", x"cf", x"d1", x"d0", 
        x"cf", x"cf", x"ce", x"ce", x"ce", x"ce", x"cf", x"cf", x"ce", x"ce", x"cd", x"ce", x"d0", x"d1", x"ce", 
        x"d0", x"cf", x"b1", x"96", x"ae", x"ce", x"d1", x"cc", x"cc", x"cf", x"cb", x"ca", x"cc", x"cb", x"cd", 
        x"ce", x"ce", x"cd", x"cd", x"ce", x"ce", x"cc", x"d9", x"da", x"d0", x"d0", x"d1", x"d2", x"d2", x"cc", 
        x"a4", x"68", x"61", x"5e", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"9d", x"d8", x"e1", x"f8", x"fb", x"fb", x"fa", x"ef", x"a8", 
        x"61", x"62", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"6c", x"c3", 
        x"ea", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ed", x"ef", x"ee", x"ee", x"ef", x"f0", 
        x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", 
        x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ec", x"ec", x"ed", x"ee", x"ee", x"ef", x"ef", x"ee", 
        x"ef", x"ef", x"f0", x"ef", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"ef", x"f2", x"ef", x"eb", x"e4", x"d0", 
        x"c6", x"d1", x"de", x"da", x"c3", x"97", x"7a", x"72", x"7c", x"7d", x"7d", x"80", x"80", x"81", x"7f", 
        x"7c", x"7c", x"7f", x"7d", x"7d", x"7f", x"7f", x"7e", x"7c", x"7e", x"7e", x"7e", x"7c", x"7d", x"7e", 
        x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7f", x"82", x"7f", x"7f", x"7e", x"7c", x"7b", x"7b", x"7c", 
        x"7c", x"7c", x"7d", x"7c", x"7d", x"7e", x"7e", x"7d", x"7c", x"7b", x"7c", x"7d", x"7c", x"7c", x"7c", 
        x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7c", x"7d", x"7d", x"7d", x"7e", x"7d", x"7c", x"7b", x"7a", 
        x"7a", x"7b", x"7b", x"7c", x"7c", x"7c", x"7c", x"7b", x"7a", x"7b", x"7c", x"7b", x"7b", x"7b", x"7a", 
        x"7a", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"78", x"7a", x"7c", x"7a", x"7b", x"79", x"7a", 
        x"7c", x"7c", x"7d", x"7b", x"7a", x"7c", x"7c", x"7b", x"7c", x"7d", x"7b", x"7a", x"7b", x"7b", x"77", 
        x"78", x"77", x"77", x"77", x"78", x"79", x"79", x"79", x"7c", x"7c", x"78", x"78", x"7a", x"7c", x"7a", 
        x"7a", x"7a", x"79", x"7a", x"7b", x"7b", x"7a", x"7a", x"7a", x"7b", x"7b", x"7a", x"7a", x"79", x"79", 
        x"7a", x"7b", x"7b", x"7a", x"78", x"78", x"7b", x"7a", x"79", x"7a", x"7b", x"7b", x"7a", x"7c", x"7b", 
        x"7a", x"7a", x"79", x"78", x"7a", x"78", x"78", x"7a", x"7b", x"7b", x"7b", x"7a", x"78", x"77", x"78", 
        x"7a", x"7b", x"7a", x"79", x"7a", x"7b", x"7b", x"7a", x"7a", x"7a", x"79", x"78", x"77", x"77", x"77", 
        x"77", x"78", x"78", x"77", x"78", x"74", x"77", x"77", x"73", x"75", x"77", x"77", x"76", x"75", x"77", 
        x"78", x"77", x"76", x"76", x"76", x"75", x"76", x"76", x"76", x"74", x"75", x"76", x"76", x"77", x"77", 
        x"77", x"77", x"78", x"76", x"73", x"74", x"73", x"75", x"77", x"74", x"73", x"75", x"74", x"73", x"75", 
        x"75", x"73", x"74", x"73", x"73", x"74", x"75", x"75", x"73", x"72", x"76", x"74", x"71", x"73", x"74", 
        x"73", x"72", x"73", x"76", x"73", x"72", x"76", x"75", x"73", x"74", x"74", x"76", x"77", x"75", x"75", 
        x"77", x"76", x"75", x"72", x"75", x"75", x"72", x"73", x"75", x"73", x"71", x"72", x"74", x"74", x"74", 
        x"73", x"72", x"73", x"72", x"73", x"73", x"72", x"74", x"74", x"73", x"74", x"76", x"76", x"73", x"72", 
        x"70", x"6f", x"73", x"74", x"71", x"74", x"75", x"74", x"75", x"75", x"74", x"73", x"73", x"73", x"72", 
        x"72", x"72", x"73", x"75", x"75", x"74", x"75", x"72", x"72", x"75", x"76", x"74", x"74", x"75", x"72", 
        x"76", x"77", x"76", x"74", x"73", x"71", x"70", x"6e", x"6e", x"71", x"72", x"70", x"70", x"71", x"72", 
        x"72", x"71", x"70", x"70", x"73", x"73", x"72", x"71", x"73", x"73", x"71", x"71", x"72", x"74", x"74", 
        x"73", x"72", x"70", x"71", x"71", x"72", x"70", x"72", x"73", x"71", x"71", x"72", x"70", x"70", x"71", 
        x"72", x"72", x"71", x"71", x"72", x"73", x"74", x"74", x"72", x"71", x"72", x"75", x"74", x"70", x"6f", 
        x"71", x"71", x"6f", x"6f", x"71", x"72", x"70", x"6f", x"70", x"72", x"73", x"74", x"74", x"75", x"70", 
        x"71", x"75", x"71", x"75", x"75", x"74", x"74", x"72", x"72", x"73", x"71", x"73", x"74", x"74", x"74", 
        x"75", x"75", x"76", x"74", x"74", x"76", x"76", x"74", x"74", x"75", x"72", x"70", x"74", x"76", x"75", 
        x"76", x"79", x"79", x"72", x"74", x"73", x"72", x"74", x"75", x"73", x"76", x"76", x"77", x"76", x"75", 
        x"77", x"77", x"77", x"77", x"75", x"74", x"76", x"78", x"77", x"78", x"77", x"75", x"75", x"75", x"73", 
        x"73", x"73", x"74", x"76", x"76", x"78", x"78", x"78", x"79", x"76", x"79", x"78", x"78", x"79", x"73", 
        x"88", x"d2", x"d4", x"d2", x"d2", x"d2", x"da", x"d5", x"cc", x"cd", x"cd", x"cd", x"cf", x"d1", x"d0", 
        x"cf", x"cf", x"ce", x"ce", x"ce", x"ce", x"cf", x"cd", x"cf", x"d0", x"cf", x"d1", x"d2", x"d2", x"d1", 
        x"c0", x"9d", x"97", x"c1", x"cf", x"cc", x"d0", x"cc", x"cd", x"cf", x"ce", x"cd", x"ce", x"ce", x"ce", 
        x"ce", x"ce", x"cd", x"cd", x"cd", x"cd", x"cb", x"d9", x"da", x"d0", x"d1", x"d1", x"d1", x"d2", x"cc", 
        x"a6", x"68", x"61", x"5e", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"60", x"8f", x"d3", x"d2", x"f7", x"fb", x"fb", x"fa", x"f9", x"d3", 
        x"79", x"5f", x"5d", x"5c", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"6b", x"be", 
        x"eb", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"ec", x"ee", x"f2", x"f1", x"ef", 
        x"e6", x"d2", x"c8", x"d0", x"e0", x"e2", x"cc", x"a2", x"7e", x"73", x"76", x"77", x"7d", x"81", x"80", 
        x"7e", x"7d", x"7e", x"80", x"7f", x"7e", x"7d", x"7d", x"7b", x"7b", x"7e", x"80", x"7e", x"7f", x"7f", 
        x"7f", x"7f", x"7e", x"7e", x"7d", x"7d", x"7e", x"80", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7c", 
        x"7c", x"7d", x"7c", x"7c", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7d", x"7e", x"7e", 
        x"7e", x"7e", x"7b", x"79", x"7b", x"7b", x"7c", x"7c", x"7d", x"7d", x"7c", x"7b", x"7b", x"7b", x"7b", 
        x"7c", x"7c", x"7c", x"7d", x"7d", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", x"7c", x"7c", x"7c", x"7b", 
        x"7a", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"78", x"78", x"7a", x"79", x"79", x"77", x"76", 
        x"7a", x"7d", x"7d", x"7b", x"7a", x"7c", x"7d", x"7c", x"7c", x"7b", x"7a", x"7a", x"7a", x"78", x"74", 
        x"78", x"79", x"7a", x"7a", x"7a", x"7a", x"7a", x"79", x"7c", x"7d", x"7b", x"7a", x"7b", x"7d", x"7c", 
        x"7a", x"7a", x"7b", x"7b", x"79", x"7a", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7a", x"7b", 
        x"7b", x"7a", x"7a", x"7a", x"79", x"79", x"79", x"7a", x"7b", x"7c", x"7c", x"7a", x"79", x"7c", x"7a", 
        x"79", x"7a", x"7a", x"79", x"79", x"7a", x"7a", x"7a", x"7a", x"7a", x"7a", x"7b", x"7a", x"79", x"7b", 
        x"7c", x"7b", x"79", x"77", x"78", x"7b", x"7c", x"7b", x"7a", x"79", x"79", x"79", x"7a", x"78", x"77", 
        x"77", x"77", x"76", x"76", x"78", x"77", x"79", x"78", x"74", x"75", x"78", x"75", x"72", x"72", x"75", 
        x"76", x"75", x"76", x"78", x"77", x"77", x"78", x"78", x"76", x"75", x"75", x"77", x"76", x"75", x"75", 
        x"75", x"76", x"76", x"74", x"73", x"75", x"75", x"76", x"77", x"75", x"73", x"75", x"75", x"73", x"73", 
        x"73", x"73", x"73", x"74", x"75", x"75", x"74", x"74", x"74", x"75", x"76", x"74", x"72", x"73", x"74", 
        x"74", x"75", x"76", x"76", x"75", x"74", x"73", x"71", x"71", x"73", x"71", x"72", x"74", x"73", x"74", 
        x"76", x"76", x"72", x"71", x"76", x"76", x"73", x"74", x"75", x"74", x"73", x"72", x"72", x"72", x"72", 
        x"76", x"74", x"74", x"72", x"73", x"73", x"72", x"74", x"75", x"75", x"76", x"77", x"78", x"75", x"73", 
        x"74", x"73", x"73", x"73", x"72", x"75", x"74", x"72", x"75", x"75", x"74", x"75", x"76", x"74", x"74", 
        x"73", x"72", x"72", x"73", x"74", x"74", x"75", x"73", x"73", x"75", x"75", x"74", x"74", x"75", x"73", 
        x"71", x"73", x"75", x"75", x"74", x"73", x"74", x"70", x"6f", x"70", x"71", x"70", x"70", x"6f", x"71", 
        x"72", x"71", x"71", x"71", x"71", x"71", x"70", x"71", x"73", x"72", x"70", x"6f", x"71", x"73", x"72", 
        x"74", x"74", x"72", x"71", x"70", x"71", x"70", x"72", x"71", x"70", x"70", x"72", x"71", x"72", x"72", 
        x"73", x"73", x"71", x"70", x"72", x"72", x"73", x"73", x"72", x"71", x"71", x"74", x"73", x"71", x"72", 
        x"75", x"75", x"73", x"72", x"74", x"74", x"71", x"70", x"71", x"72", x"73", x"72", x"73", x"73", x"72", 
        x"74", x"77", x"73", x"73", x"73", x"75", x"76", x"75", x"74", x"74", x"76", x"72", x"72", x"72", x"73", 
        x"73", x"74", x"73", x"74", x"76", x"77", x"76", x"75", x"73", x"74", x"74", x"75", x"77", x"77", x"77", 
        x"76", x"78", x"78", x"75", x"77", x"75", x"74", x"76", x"76", x"75", x"75", x"75", x"76", x"74", x"73", 
        x"74", x"75", x"77", x"76", x"75", x"75", x"76", x"76", x"75", x"76", x"75", x"74", x"75", x"77", x"77", 
        x"76", x"76", x"77", x"79", x"79", x"78", x"76", x"76", x"77", x"77", x"7a", x"79", x"78", x"78", x"73", 
        x"87", x"d3", x"d5", x"d3", x"d3", x"d3", x"dc", x"d7", x"cd", x"ce", x"ce", x"ce", x"cf", x"d1", x"d0", 
        x"d0", x"cf", x"ce", x"ce", x"ce", x"ce", x"ce", x"cf", x"d1", x"d3", x"cf", x"d1", x"d5", x"c7", x"ac", 
        x"98", x"ac", x"d0", x"cf", x"ce", x"d2", x"cd", x"d1", x"cf", x"ce", x"cf", x"d0", x"ce", x"cd", x"ce", 
        x"cf", x"cf", x"ce", x"ce", x"ce", x"ce", x"cb", x"d9", x"d9", x"d0", x"d2", x"d0", x"d0", x"d2", x"cc", 
        x"a9", x"67", x"61", x"5e", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5c", x"62", x"7a", x"cf", x"ca", x"ee", x"fb", x"fc", x"fc", x"fa", x"eb", 
        x"a9", x"61", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"6a", x"b7", 
        x"ea", x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"f0", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"ed", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"eb", x"ee", x"f1", x"ef", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"eb", x"de", x"cf", x"d4", x"d8", x"df", x"d5", x"b1", x"8a", x"74", x"74", x"79", x"7d", 
        x"80", x"80", x"80", x"7e", x"7f", x"7f", x"7d", x"7e", x"7d", x"7b", x"7c", x"7f", x"7f", x"7e", x"7e", 
        x"7e", x"7e", x"7f", x"7f", x"7e", x"7c", x"7d", x"7f", x"7c", x"7d", x"7e", x"7e", x"7f", x"7e", x"7c", 
        x"7c", x"7e", x"7c", x"7c", x"7c", x"7b", x"7c", x"7e", x"7e", x"7e", x"7d", x"7d", x"7e", x"7e", x"7d", 
        x"7e", x"7e", x"7c", x"7c", x"7d", x"7e", x"7c", x"7b", x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", x"7d", 
        x"7d", x"7e", x"7c", x"7d", x"7d", x"7c", x"7b", x"7b", x"7b", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", 
        x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7c", x"7d", x"7d", x"7d", x"7b", x"7a", 
        x"7b", x"7d", x"7e", x"7d", x"7c", x"7d", x"7e", x"7d", x"7d", x"7b", x"7a", x"7b", x"7b", x"7a", x"77", 
        x"79", x"7a", x"7a", x"7a", x"79", x"7a", x"7c", x"7c", x"7d", x"7e", x"7d", x"7c", x"7b", x"7a", x"7c", 
        x"7b", x"7c", x"7d", x"7c", x"79", x"7a", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", 
        x"7b", x"7a", x"7a", x"7a", x"7a", x"7a", x"78", x"78", x"7a", x"7a", x"7a", x"79", x"78", x"7c", x"7a", 
        x"79", x"7b", x"7b", x"79", x"7a", x"7b", x"7c", x"7a", x"7a", x"79", x"7a", x"7a", x"7a", x"79", x"7a", 
        x"7b", x"7b", x"7a", x"7a", x"79", x"79", x"7a", x"7a", x"78", x"77", x"78", x"79", x"78", x"77", x"77", 
        x"78", x"79", x"78", x"77", x"77", x"77", x"78", x"77", x"75", x"76", x"78", x"78", x"75", x"74", x"77", 
        x"78", x"76", x"76", x"78", x"78", x"77", x"78", x"79", x"78", x"77", x"77", x"78", x"76", x"75", x"74", 
        x"75", x"76", x"75", x"72", x"73", x"74", x"75", x"76", x"76", x"76", x"73", x"74", x"75", x"74", x"73", 
        x"73", x"74", x"73", x"74", x"75", x"75", x"74", x"73", x"74", x"76", x"75", x"72", x"72", x"74", x"75", 
        x"76", x"75", x"73", x"72", x"74", x"76", x"75", x"74", x"75", x"75", x"71", x"72", x"74", x"73", x"72", 
        x"75", x"77", x"72", x"73", x"78", x"77", x"75", x"75", x"73", x"74", x"76", x"75", x"73", x"72", x"73", 
        x"75", x"73", x"73", x"72", x"73", x"74", x"73", x"73", x"75", x"76", x"75", x"76", x"77", x"74", x"72", 
        x"76", x"75", x"73", x"71", x"72", x"74", x"72", x"72", x"74", x"75", x"75", x"76", x"76", x"75", x"73", 
        x"73", x"72", x"73", x"73", x"73", x"74", x"74", x"74", x"74", x"75", x"75", x"75", x"75", x"75", x"75", 
        x"71", x"72", x"74", x"74", x"72", x"72", x"72", x"72", x"70", x"6f", x"70", x"71", x"71", x"6f", x"6e", 
        x"6d", x"6f", x"72", x"74", x"73", x"73", x"72", x"71", x"72", x"70", x"6d", x"6d", x"6f", x"71", x"72", 
        x"74", x"76", x"74", x"72", x"70", x"6f", x"71", x"71", x"70", x"6f", x"71", x"72", x"71", x"71", x"70", 
        x"71", x"73", x"72", x"72", x"75", x"73", x"71", x"72", x"72", x"72", x"71", x"72", x"74", x"74", x"74", 
        x"75", x"74", x"71", x"70", x"72", x"73", x"71", x"71", x"72", x"73", x"73", x"73", x"71", x"72", x"72", 
        x"76", x"76", x"75", x"75", x"74", x"77", x"79", x"77", x"73", x"72", x"77", x"75", x"74", x"73", x"73", 
        x"74", x"75", x"76", x"75", x"74", x"75", x"75", x"75", x"75", x"77", x"77", x"76", x"75", x"75", x"76", 
        x"76", x"75", x"75", x"75", x"77", x"75", x"74", x"75", x"75", x"74", x"73", x"76", x"77", x"77", x"76", 
        x"75", x"76", x"77", x"76", x"77", x"78", x"79", x"77", x"76", x"77", x"79", x"77", x"77", x"78", x"7a", 
        x"79", x"78", x"78", x"7a", x"7a", x"78", x"77", x"77", x"77", x"77", x"79", x"79", x"78", x"79", x"76", 
        x"88", x"d4", x"d6", x"d4", x"d4", x"d4", x"dd", x"d8", x"ce", x"ce", x"ce", x"ce", x"d0", x"d1", x"d0", 
        x"d0", x"d0", x"ce", x"ce", x"ce", x"ce", x"ce", x"d0", x"cc", x"ce", x"d5", x"cf", x"b9", x"a2", x"9d", 
        x"bd", x"d0", x"ce", x"cc", x"cd", x"cd", x"cc", x"ce", x"ce", x"cd", x"cd", x"cd", x"cb", x"cc", x"cf", 
        x"d0", x"cf", x"ce", x"ce", x"ce", x"cd", x"cb", x"da", x"d8", x"ce", x"d3", x"d0", x"cf", x"d2", x"cd", 
        x"ac", x"67", x"61", x"5e", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"6a", x"c1", x"d0", x"e1", x"fb", x"fc", x"fb", x"f9", x"f5", 
        x"d4", x"7f", x"5b", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5f", x"67", x"b0", 
        x"ea", x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"ef", x"ef", x"ef", x"ee", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"ef", x"ee", x"f2", 
        x"f0", x"ed", x"f0", x"f2", x"ef", x"e3", x"d6", x"d4", x"da", x"df", x"d9", x"b5", x"90", x"7e", x"74", 
        x"75", x"7b", x"80", x"7f", x"80", x"80", x"7d", x"7d", x"7e", x"7e", x"7f", x"80", x"7f", x"7e", x"7e", 
        x"7e", x"7e", x"7f", x"7f", x"7f", x"7d", x"7d", x"7e", x"7c", x"7d", x"7f", x"7e", x"80", x"7f", x"7d", 
        x"7d", x"7e", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", x"7d", x"7d", x"7e", x"7d", x"7d", x"7d", 
        x"7c", x"7c", x"7c", x"7d", x"7e", x"7e", x"7d", x"7b", x"7b", x"7c", x"7e", x"7d", x"7d", x"7c", x"7c", 
        x"7c", x"7d", x"7d", x"7e", x"7d", x"7c", x"7b", x"7b", x"7c", x"7c", x"7c", x"7b", x"7b", x"7c", x"7d", 
        x"7d", x"7d", x"7b", x"7b", x"7b", x"7c", x"7d", x"7e", x"7d", x"7b", x"79", x"7a", x"7a", x"7b", x"7a", 
        x"79", x"7c", x"7e", x"7d", x"7d", x"7e", x"7d", x"7c", x"7c", x"78", x"77", x"79", x"7a", x"79", x"79", 
        x"7b", x"7b", x"7b", x"79", x"79", x"7b", x"7e", x"7d", x"7b", x"7a", x"7b", x"7d", x"7d", x"7c", x"7c", 
        x"7b", x"7b", x"7c", x"7c", x"79", x"7a", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7a", x"7a", 
        x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7a", x"7b", x"7b", x"7b", x"7a", 
        x"7a", x"7c", x"7c", x"7a", x"7a", x"7c", x"7c", x"7b", x"7a", x"79", x"79", x"7a", x"7b", x"7c", x"7b", 
        x"7a", x"79", x"79", x"79", x"7a", x"7a", x"7b", x"7b", x"79", x"78", x"79", x"79", x"7a", x"79", x"78", 
        x"78", x"78", x"78", x"77", x"76", x"77", x"76", x"76", x"77", x"77", x"78", x"78", x"76", x"76", x"76", 
        x"77", x"76", x"75", x"78", x"79", x"78", x"78", x"78", x"78", x"76", x"77", x"77", x"76", x"75", x"75", 
        x"75", x"76", x"75", x"72", x"74", x"74", x"75", x"75", x"74", x"75", x"73", x"73", x"74", x"75", x"74", 
        x"75", x"77", x"75", x"76", x"77", x"76", x"74", x"75", x"76", x"76", x"74", x"72", x"73", x"74", x"76", 
        x"77", x"77", x"73", x"72", x"75", x"77", x"74", x"74", x"76", x"75", x"73", x"74", x"75", x"75", x"74", 
        x"77", x"77", x"74", x"75", x"77", x"77", x"77", x"75", x"74", x"74", x"76", x"75", x"73", x"73", x"75", 
        x"75", x"71", x"72", x"71", x"73", x"74", x"73", x"74", x"75", x"74", x"74", x"74", x"75", x"74", x"71", 
        x"74", x"73", x"71", x"71", x"72", x"75", x"72", x"72", x"72", x"75", x"77", x"76", x"75", x"76", x"73", 
        x"74", x"75", x"76", x"76", x"76", x"76", x"74", x"75", x"75", x"74", x"75", x"76", x"75", x"74", x"75", 
        x"75", x"73", x"74", x"72", x"70", x"70", x"70", x"74", x"74", x"72", x"71", x"71", x"70", x"6e", x"70", 
        x"70", x"71", x"74", x"73", x"70", x"6e", x"70", x"73", x"72", x"72", x"70", x"71", x"73", x"74", x"72", 
        x"73", x"74", x"74", x"74", x"72", x"71", x"72", x"72", x"70", x"70", x"72", x"74", x"73", x"74", x"71", 
        x"71", x"74", x"74", x"72", x"75", x"73", x"72", x"72", x"73", x"73", x"73", x"73", x"75", x"76", x"75", 
        x"76", x"75", x"72", x"71", x"73", x"72", x"71", x"72", x"74", x"75", x"75", x"74", x"76", x"75", x"73", 
        x"74", x"72", x"75", x"74", x"73", x"76", x"76", x"76", x"74", x"72", x"76", x"77", x"75", x"75", x"74", 
        x"75", x"76", x"77", x"76", x"74", x"72", x"72", x"74", x"75", x"76", x"76", x"74", x"74", x"74", x"74", 
        x"74", x"73", x"74", x"75", x"76", x"74", x"73", x"74", x"74", x"73", x"73", x"74", x"72", x"74", x"76", 
        x"76", x"78", x"76", x"75", x"76", x"78", x"77", x"76", x"76", x"78", x"79", x"78", x"76", x"77", x"7a", 
        x"7a", x"7b", x"7a", x"7a", x"7b", x"78", x"78", x"78", x"77", x"77", x"78", x"79", x"79", x"79", x"78", 
        x"87", x"d4", x"d7", x"d4", x"d4", x"d4", x"dd", x"d8", x"ce", x"ce", x"cf", x"cd", x"cf", x"d0", x"d0", 
        x"d0", x"d0", x"ce", x"ce", x"ce", x"cd", x"ce", x"ce", x"ce", x"d3", x"cb", x"a6", x"95", x"ae", x"cc", 
        x"d0", x"cd", x"cb", x"cb", x"cf", x"cf", x"ca", x"cb", x"cf", x"ce", x"ce", x"cd", x"cc", x"cf", x"d0", 
        x"d0", x"d0", x"cf", x"ce", x"ce", x"cd", x"ca", x"da", x"d6", x"cd", x"d4", x"d0", x"cf", x"d3", x"cd", 
        x"ae", x"67", x"61", x"5e", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5a", x"60", x"a2", x"d7", x"df", x"f9", x"fb", x"fa", x"f8", x"fa", 
        x"f1", x"b6", x"6b", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"65", x"a9", 
        x"e9", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ee", x"ef", x"f0", x"ee", x"ed", 
        x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"f1", x"f1", x"f1", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"f1", x"ef", x"ef", x"f1", x"f2", x"f0", x"e8", x"d9", x"d5", x"dc", x"e3", x"df", x"c8", x"a0", 
        x"80", x"70", x"6f", x"7a", x"80", x"80", x"7f", x"7e", x"7d", x"7d", x"7f", x"80", x"7f", x"7f", x"7e", 
        x"7e", x"7e", x"7f", x"80", x"80", x"7e", x"7e", x"7f", x"7d", x"7d", x"7f", x"7f", x"7f", x"7e", x"7f", 
        x"7e", x"7e", x"7e", x"7f", x"7e", x"7d", x"7c", x"7c", x"7c", x"7c", x"7d", x"7d", x"7d", x"7d", x"7d", 
        x"7d", x"7d", x"7d", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"7e", x"7e", x"7d", x"7d", x"7d", 
        x"7d", x"7e", x"7e", x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", x"7d", x"7d", x"7c", x"7c", x"7d", x"7d", 
        x"7e", x"7d", x"7d", x"7c", x"7b", x"7c", x"7d", x"7e", x"7e", x"7c", x"7a", x"7a", x"79", x"7b", x"7d", 
        x"7b", x"7b", x"7d", x"7c", x"7c", x"7d", x"7c", x"7b", x"7c", x"78", x"78", x"7b", x"7b", x"7b", x"7c", 
        x"7a", x"7a", x"7a", x"78", x"78", x"79", x"7d", x"7f", x"7c", x"79", x"7b", x"7c", x"7c", x"7c", x"7b", 
        x"7b", x"7b", x"7a", x"7a", x"7b", x"7b", x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7a", x"7b", x"7c", 
        x"7b", x"79", x"79", x"7b", x"7c", x"7d", x"7a", x"79", x"79", x"78", x"77", x"78", x"7a", x"7b", x"7a", 
        x"7b", x"7d", x"7c", x"7a", x"7a", x"7c", x"7c", x"7b", x"7a", x"7a", x"7a", x"7a", x"7c", x"7c", x"7b", 
        x"7a", x"79", x"79", x"7a", x"7b", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7a", x"79", x"78", x"78", 
        x"78", x"7a", x"79", x"78", x"77", x"79", x"76", x"76", x"7a", x"79", x"78", x"79", x"79", x"78", x"76", 
        x"77", x"78", x"76", x"78", x"7a", x"77", x"77", x"76", x"77", x"76", x"76", x"77", x"76", x"76", x"76", 
        x"76", x"77", x"76", x"75", x"77", x"76", x"76", x"75", x"73", x"75", x"75", x"74", x"74", x"76", x"75", 
        x"74", x"76", x"77", x"77", x"77", x"75", x"75", x"76", x"78", x"78", x"73", x"74", x"77", x"75", x"76", 
        x"78", x"76", x"73", x"73", x"76", x"77", x"74", x"75", x"76", x"72", x"71", x"73", x"74", x"74", x"74", 
        x"76", x"76", x"77", x"77", x"74", x"75", x"77", x"74", x"75", x"75", x"75", x"73", x"72", x"73", x"75", 
        x"75", x"73", x"74", x"73", x"75", x"76", x"74", x"76", x"75", x"74", x"73", x"74", x"74", x"74", x"73", 
        x"73", x"74", x"74", x"75", x"76", x"79", x"76", x"73", x"73", x"75", x"77", x"76", x"75", x"76", x"75", 
        x"76", x"78", x"78", x"77", x"77", x"77", x"74", x"75", x"76", x"75", x"74", x"76", x"76", x"73", x"75", 
        x"74", x"71", x"72", x"72", x"71", x"74", x"72", x"70", x"70", x"72", x"73", x"72", x"72", x"72", x"72", 
        x"70", x"70", x"72", x"72", x"70", x"70", x"73", x"74", x"73", x"71", x"71", x"72", x"73", x"74", x"75", 
        x"74", x"73", x"73", x"73", x"72", x"72", x"73", x"73", x"71", x"71", x"74", x"76", x"75", x"76", x"72", 
        x"71", x"74", x"73", x"72", x"74", x"75", x"74", x"73", x"73", x"73", x"74", x"75", x"75", x"73", x"72", 
        x"72", x"73", x"71", x"71", x"74", x"73", x"73", x"74", x"75", x"74", x"72", x"72", x"76", x"77", x"76", 
        x"74", x"71", x"73", x"72", x"73", x"72", x"71", x"73", x"75", x"71", x"73", x"73", x"73", x"75", x"77", 
        x"77", x"75", x"74", x"76", x"75", x"71", x"70", x"73", x"75", x"75", x"75", x"77", x"78", x"78", x"75", 
        x"74", x"75", x"77", x"77", x"78", x"76", x"74", x"76", x"76", x"74", x"75", x"76", x"73", x"75", x"77", 
        x"75", x"75", x"77", x"75", x"76", x"78", x"77", x"76", x"79", x"79", x"7a", x"79", x"75", x"75", x"78", 
        x"7a", x"7b", x"7a", x"79", x"7a", x"78", x"7a", x"7b", x"7a", x"7b", x"7a", x"7b", x"79", x"78", x"75", 
        x"83", x"d3", x"d5", x"d3", x"d3", x"d3", x"dc", x"d7", x"ce", x"ce", x"ce", x"cd", x"ce", x"cf", x"cf", 
        x"d0", x"d0", x"cf", x"cd", x"cd", x"cd", x"ce", x"d1", x"d3", x"b5", x"96", x"a6", x"c3", x"d0", x"d3", 
        x"cd", x"cc", x"ce", x"cd", x"ce", x"cf", x"ca", x"ce", x"ce", x"cb", x"cd", x"cf", x"cd", x"d0", x"d0", 
        x"d1", x"d0", x"cf", x"ce", x"ce", x"cd", x"ca", x"da", x"d5", x"cc", x"d4", x"d0", x"cf", x"d3", x"cd", 
        x"af", x"67", x"61", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"62", x"5e", x"7b", x"d0", x"eb", x"f5", x"f9", x"fb", x"fb", x"fa", 
        x"f7", x"e4", x"a8", x"6f", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", x"5e", x"5d", 
        x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"64", x"a5", 
        x"e8", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"f1", x"ef", x"ed", 
        x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"f0", x"f1", x"ee", x"ef", x"f1", x"ef", x"ef", 
        x"f0", x"f1", x"ef", x"f0", x"f1", x"f1", x"ee", x"f2", x"f0", x"e7", x"e4", x"de", x"dc", x"e0", x"e1", 
        x"d3", x"b3", x"8e", x"77", x"72", x"7a", x"80", x"82", x"7f", x"7f", x"7f", x"80", x"80", x"80", x"7f", 
        x"7f", x"80", x"80", x"81", x"80", x"7f", x"7f", x"80", x"7d", x"7e", x"7f", x"7f", x"7d", x"7e", x"7f", 
        x"7f", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7e", x"7d", x"7d", x"7d", x"7d", x"7e", 
        x"7e", x"7e", x"7f", x"7f", x"7e", x"7d", x"7e", x"7f", x"7f", x"7f", x"7e", x"7e", x"7d", x"7d", x"7d", 
        x"7e", x"7f", x"7f", x"7d", x"7c", x"7c", x"7d", x"7d", x"7c", x"7c", x"7c", x"7d", x"7e", x"7e", x"7e", 
        x"7e", x"7f", x"7e", x"7c", x"7b", x"7b", x"7c", x"7d", x"7e", x"7c", x"7d", x"7d", x"78", x"7a", x"80", 
        x"7f", x"7c", x"7d", x"7b", x"7a", x"7c", x"7c", x"7c", x"7b", x"7a", x"7c", x"7d", x"7c", x"7b", x"7d", 
        x"7a", x"7c", x"7d", x"7b", x"7a", x"7b", x"7d", x"7e", x"7c", x"7c", x"7e", x"7d", x"79", x"79", x"79", 
        x"7a", x"7a", x"79", x"79", x"7c", x"7b", x"7a", x"7a", x"7a", x"7b", x"7b", x"7a", x"7a", x"7a", x"7a", 
        x"7a", x"7b", x"7c", x"7c", x"7c", x"7b", x"7a", x"7a", x"7b", x"79", x"78", x"79", x"7a", x"7b", x"7b", 
        x"7c", x"7d", x"7b", x"79", x"7a", x"7b", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", x"7c", x"7b", x"7b", 
        x"7b", x"7a", x"79", x"79", x"7a", x"7c", x"7b", x"7a", x"7a", x"7a", x"79", x"79", x"7a", x"79", x"79", 
        x"79", x"79", x"79", x"78", x"7a", x"7c", x"77", x"76", x"7c", x"7a", x"78", x"77", x"79", x"78", x"75", 
        x"78", x"7b", x"78", x"77", x"77", x"76", x"75", x"76", x"77", x"78", x"77", x"77", x"76", x"77", x"77", 
        x"77", x"77", x"77", x"78", x"7a", x"78", x"77", x"75", x"72", x"75", x"75", x"73", x"74", x"77", x"76", 
        x"75", x"76", x"76", x"75", x"73", x"72", x"72", x"74", x"76", x"77", x"74", x"77", x"7a", x"75", x"74", 
        x"77", x"76", x"74", x"75", x"77", x"76", x"73", x"74", x"76", x"75", x"74", x"76", x"75", x"73", x"72", 
        x"74", x"74", x"77", x"77", x"71", x"72", x"76", x"72", x"75", x"75", x"75", x"74", x"72", x"71", x"72", 
        x"76", x"76", x"78", x"77", x"78", x"77", x"76", x"77", x"77", x"75", x"75", x"75", x"75", x"77", x"76", 
        x"74", x"74", x"76", x"76", x"75", x"78", x"74", x"74", x"75", x"75", x"75", x"76", x"76", x"75", x"75", 
        x"75", x"75", x"73", x"72", x"73", x"74", x"73", x"76", x"77", x"75", x"74", x"76", x"76", x"75", x"77", 
        x"76", x"73", x"72", x"72", x"73", x"74", x"73", x"71", x"70", x"71", x"71", x"70", x"71", x"72", x"71", 
        x"72", x"73", x"74", x"73", x"71", x"70", x"72", x"73", x"71", x"70", x"73", x"71", x"72", x"72", x"73", 
        x"73", x"72", x"73", x"73", x"74", x"72", x"71", x"74", x"73", x"74", x"75", x"75", x"76", x"74", x"74", 
        x"72", x"70", x"72", x"75", x"74", x"73", x"76", x"74", x"72", x"74", x"74", x"73", x"74", x"73", x"73", 
        x"73", x"74", x"73", x"71", x"72", x"72", x"72", x"74", x"75", x"73", x"72", x"73", x"77", x"77", x"74", 
        x"74", x"75", x"74", x"75", x"76", x"73", x"72", x"73", x"73", x"73", x"73", x"74", x"73", x"75", x"77", 
        x"76", x"77", x"75", x"75", x"75", x"75", x"75", x"76", x"76", x"76", x"75", x"77", x"78", x"76", x"76", 
        x"75", x"74", x"77", x"78", x"76", x"74", x"74", x"76", x"76", x"74", x"74", x"77", x"76", x"76", x"77", 
        x"76", x"75", x"78", x"75", x"75", x"78", x"78", x"77", x"78", x"79", x"7b", x"7a", x"76", x"76", x"79", 
        x"7a", x"7a", x"77", x"76", x"79", x"7a", x"7a", x"7b", x"7a", x"79", x"79", x"7a", x"7a", x"79", x"75", 
        x"85", x"d4", x"d6", x"d2", x"d2", x"d3", x"dc", x"d6", x"cc", x"d0", x"cf", x"cf", x"ce", x"cd", x"cf", 
        x"d0", x"d1", x"cd", x"cc", x"cf", x"ce", x"d3", x"cb", x"a5", x"9a", x"b2", x"cc", x"d0", x"cd", x"ce", 
        x"cd", x"cd", x"ce", x"cd", x"cd", x"cd", x"cf", x"cf", x"ce", x"cb", x"cc", x"ce", x"ce", x"d0", x"cf", 
        x"cf", x"d0", x"cf", x"cf", x"ce", x"ce", x"cb", x"d9", x"d7", x"cc", x"d3", x"d1", x"ce", x"d1", x"cc", 
        x"ac", x"67", x"60", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5f", x"63", x"60", x"63", x"af", x"eb", x"f5", x"f9", x"f9", x"fa", x"f9", 
        x"f6", x"f7", x"e4", x"a9", x"70", x"5e", x"60", x"5c", x"5b", x"5c", x"5c", x"5d", x"5e", x"5d", x"5c", 
        x"5d", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"66", x"a4", 
        x"e6", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ee", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ef", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f1", x"ef", x"ee", x"f1", x"ec", x"e7", x"e3", x"dd", 
        x"dc", x"e1", x"d9", x"bb", x"98", x"7a", x"73", x"7b", x"80", x"82", x"83", x"81", x"82", x"80", x"7c", 
        x"7f", x"81", x"80", x"81", x"81", x"81", x"7e", x"7d", x"7d", x"80", x"81", x"80", x"7d", x"7d", x"7e", 
        x"7d", x"7d", x"7f", x"7e", x"7e", x"7f", x"7f", x"7f", x"7e", x"7e", x"7e", x"7e", x"7d", x"7e", x"7e", 
        x"7d", x"7b", x"7d", x"7f", x"7d", x"7f", x"81", x"80", x"7e", x"7d", x"7c", x"7d", x"7c", x"7c", x"7d", 
        x"7d", x"7b", x"7b", x"7e", x"7e", x"7e", x"7e", x"7c", x"7d", x"7e", x"7b", x"7c", x"7e", x"7d", x"7c", 
        x"7c", x"7f", x"7e", x"7d", x"7c", x"7c", x"7d", x"7e", x"7f", x"7f", x"7e", x"7d", x"7a", x"7c", x"7f", 
        x"7f", x"7d", x"7e", x"7e", x"7c", x"7c", x"7d", x"7d", x"7a", x"7a", x"7b", x"7c", x"7c", x"7d", x"7d", 
        x"7d", x"7c", x"7c", x"7b", x"7c", x"7c", x"7d", x"7d", x"7a", x"7a", x"7e", x"7f", x"7b", x"7a", x"7b", 
        x"7b", x"7a", x"7b", x"7b", x"7a", x"7a", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7c", x"7d", 
        x"7b", x"7c", x"7e", x"7d", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", 
        x"7e", x"7d", x"7a", x"7b", x"7b", x"79", x"7b", x"7c", x"7b", x"79", x"7b", x"7d", x"7e", x"7b", x"7a", 
        x"7a", x"7a", x"7a", x"7a", x"78", x"79", x"7b", x"7b", x"79", x"78", x"79", x"7b", x"7c", x"7a", x"7a", 
        x"79", x"79", x"7a", x"79", x"7a", x"7a", x"78", x"78", x"7b", x"7b", x"7b", x"79", x"78", x"78", x"77", 
        x"79", x"7a", x"78", x"77", x"77", x"77", x"78", x"79", x"79", x"79", x"79", x"7a", x"77", x"75", x"77", 
        x"76", x"76", x"78", x"77", x"79", x"78", x"78", x"76", x"74", x"75", x"76", x"76", x"75", x"77", x"77", 
        x"75", x"76", x"75", x"77", x"75", x"74", x"76", x"76", x"75", x"75", x"77", x"77", x"75", x"75", x"76", 
        x"77", x"78", x"76", x"76", x"76", x"78", x"75", x"76", x"75", x"73", x"74", x"75", x"75", x"75", x"75", 
        x"76", x"75", x"76", x"76", x"72", x"72", x"75", x"74", x"73", x"75", x"75", x"75", x"74", x"74", x"76", 
        x"76", x"77", x"78", x"76", x"75", x"76", x"77", x"78", x"77", x"75", x"74", x"73", x"74", x"77", x"76", 
        x"75", x"75", x"76", x"75", x"75", x"78", x"77", x"75", x"75", x"75", x"75", x"76", x"77", x"76", x"75", 
        x"75", x"74", x"74", x"74", x"76", x"77", x"78", x"75", x"77", x"79", x"76", x"75", x"76", x"76", x"76", 
        x"74", x"73", x"72", x"72", x"73", x"74", x"75", x"73", x"71", x"72", x"73", x"72", x"74", x"75", x"72", 
        x"71", x"72", x"73", x"73", x"72", x"71", x"74", x"74", x"72", x"71", x"74", x"70", x"6f", x"6f", x"70", 
        x"71", x"71", x"73", x"72", x"74", x"74", x"72", x"75", x"73", x"74", x"75", x"72", x"74", x"73", x"75", 
        x"74", x"71", x"73", x"77", x"75", x"70", x"73", x"73", x"72", x"75", x"75", x"74", x"75", x"74", x"74", 
        x"72", x"72", x"74", x"73", x"75", x"73", x"71", x"73", x"73", x"73", x"74", x"76", x"74", x"74", x"71", 
        x"73", x"76", x"73", x"76", x"75", x"72", x"74", x"74", x"73", x"76", x"76", x"77", x"74", x"75", x"76", 
        x"74", x"76", x"75", x"74", x"75", x"76", x"76", x"77", x"76", x"75", x"74", x"75", x"75", x"72", x"74", 
        x"75", x"75", x"78", x"77", x"74", x"73", x"75", x"76", x"74", x"74", x"77", x"78", x"77", x"76", x"77", 
        x"76", x"74", x"79", x"77", x"76", x"79", x"7a", x"78", x"76", x"78", x"79", x"78", x"77", x"78", x"79", 
        x"7b", x"7a", x"78", x"76", x"79", x"7a", x"79", x"78", x"78", x"76", x"78", x"79", x"7a", x"7b", x"76", 
        x"88", x"d5", x"d5", x"d2", x"d2", x"d3", x"dd", x"d6", x"cd", x"ce", x"cf", x"cf", x"d0", x"d5", x"ce", 
        x"cb", x"ce", x"ce", x"ce", x"d2", x"d4", x"b4", x"96", x"a8", x"c8", x"d0", x"cc", x"ce", x"cc", x"cd", 
        x"ce", x"ce", x"ce", x"cc", x"cc", x"cd", x"cf", x"cf", x"ce", x"cd", x"cd", x"cd", x"cf", x"d0", x"ce", 
        x"ce", x"cf", x"cf", x"cf", x"ce", x"cd", x"cc", x"da", x"db", x"cf", x"d4", x"d4", x"d1", x"d2", x"cb", 
        x"ab", x"67", x"5f", x"5d", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5d", x"5a", x"85", x"d1", x"f2", x"f5", x"f9", x"fc", x"fb", 
        x"f9", x"f8", x"f8", x"e9", x"b4", x"73", x"5e", x"58", x"5c", x"5d", x"5c", x"60", x"5e", x"5d", x"60", 
        x"61", x"5f", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5e", x"5d", x"5b", x"5c", x"67", x"a4", 
        x"e6", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ed", x"ee", x"ec", 
        x"df", x"d5", x"d6", x"e1", x"e0", x"c8", x"a0", x"7e", x"72", x"74", x"7d", x"7f", x"81", x"85", x"7e", 
        x"7d", x"80", x"81", x"7e", x"7d", x"81", x"7f", x"7a", x"7c", x"81", x"81", x"80", x"7e", x"7d", x"7e", 
        x"7d", x"7d", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", x"7d", x"7c", x"7e", x"7f", x"7e", x"7e", x"7d", 
        x"7c", x"7a", x"7d", x"80", x"7f", x"81", x"82", x"80", x"7f", x"7f", x"7e", x"7e", x"7b", x"7b", x"7c", 
        x"7e", x"7d", x"7c", x"7f", x"7f", x"80", x"80", x"7e", x"7e", x"7f", x"7c", x"7b", x"7d", x"7d", x"7b", 
        x"7c", x"7c", x"7d", x"7e", x"7f", x"7e", x"7e", x"7d", x"7e", x"7f", x"7d", x"7c", x"7b", x"7c", x"7d", 
        x"7c", x"7c", x"7e", x"7e", x"7b", x"7a", x"7c", x"7e", x"7f", x"7f", x"7e", x"7d", x"7d", x"7c", x"7c", 
        x"7c", x"7a", x"7c", x"7c", x"7e", x"7d", x"7a", x"7d", x"7b", x"7b", x"7d", x"7d", x"7b", x"7b", x"7d", 
        x"7d", x"7c", x"7e", x"7e", x"7c", x"7e", x"7e", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7c", x"7e", 
        x"7b", x"7c", x"7d", x"7c", x"7a", x"7c", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", 
        x"7e", x"7d", x"7b", x"7d", x"7e", x"7a", x"7b", x"7b", x"79", x"7a", x"7c", x"7c", x"7b", x"7a", x"7a", 
        x"7c", x"79", x"7b", x"7c", x"79", x"7a", x"7b", x"7a", x"79", x"79", x"79", x"7b", x"7a", x"79", x"7c", 
        x"7a", x"79", x"7a", x"79", x"79", x"79", x"79", x"7a", x"7b", x"7b", x"7b", x"7c", x"7a", x"78", x"77", 
        x"79", x"79", x"79", x"78", x"78", x"78", x"7a", x"7a", x"79", x"79", x"7a", x"7b", x"77", x"75", x"78", 
        x"76", x"74", x"76", x"75", x"76", x"77", x"78", x"77", x"76", x"76", x"75", x"76", x"75", x"76", x"78", 
        x"76", x"77", x"76", x"78", x"75", x"73", x"76", x"77", x"77", x"75", x"78", x"77", x"74", x"77", x"78", 
        x"77", x"78", x"76", x"75", x"75", x"79", x"76", x"76", x"75", x"73", x"73", x"74", x"75", x"75", x"76", 
        x"76", x"75", x"74", x"74", x"76", x"76", x"75", x"74", x"75", x"74", x"73", x"74", x"74", x"74", x"74", 
        x"75", x"78", x"78", x"75", x"73", x"76", x"78", x"78", x"79", x"77", x"76", x"75", x"76", x"78", x"77", 
        x"72", x"74", x"75", x"75", x"77", x"79", x"7a", x"76", x"75", x"75", x"75", x"76", x"76", x"76", x"76", 
        x"76", x"75", x"75", x"76", x"77", x"77", x"77", x"73", x"76", x"78", x"75", x"75", x"76", x"77", x"76", 
        x"74", x"74", x"74", x"73", x"73", x"73", x"74", x"73", x"71", x"73", x"74", x"74", x"76", x"76", x"73", 
        x"71", x"71", x"72", x"72", x"71", x"72", x"73", x"72", x"72", x"71", x"74", x"72", x"72", x"71", x"71", 
        x"72", x"72", x"72", x"71", x"74", x"74", x"74", x"74", x"72", x"74", x"75", x"73", x"74", x"72", x"73", 
        x"74", x"75", x"75", x"76", x"75", x"73", x"72", x"74", x"74", x"73", x"74", x"73", x"72", x"74", x"76", 
        x"74", x"72", x"73", x"73", x"76", x"75", x"72", x"72", x"73", x"73", x"75", x"78", x"72", x"72", x"72", 
        x"73", x"75", x"73", x"76", x"77", x"75", x"77", x"77", x"74", x"74", x"73", x"76", x"74", x"74", x"74", 
        x"74", x"75", x"74", x"76", x"76", x"74", x"74", x"76", x"76", x"75", x"74", x"75", x"75", x"73", x"74", 
        x"74", x"73", x"75", x"76", x"75", x"75", x"76", x"77", x"75", x"74", x"78", x"78", x"76", x"75", x"77", 
        x"77", x"74", x"78", x"77", x"76", x"78", x"79", x"78", x"78", x"79", x"78", x"76", x"78", x"78", x"77", 
        x"79", x"7b", x"7a", x"78", x"79", x"7a", x"78", x"77", x"78", x"78", x"78", x"78", x"79", x"7b", x"76", 
        x"86", x"d5", x"d5", x"d2", x"d3", x"d4", x"dd", x"d5", x"cb", x"d1", x"ce", x"cd", x"ce", x"ce", x"d0", 
        x"d0", x"cf", x"cd", x"cf", x"c1", x"97", x"96", x"b9", x"cd", x"d1", x"ce", x"c9", x"ca", x"cb", x"ce", 
        x"ce", x"cf", x"ce", x"cd", x"cd", x"cd", x"cf", x"cf", x"ce", x"cd", x"cd", x"ce", x"cf", x"d0", x"cd", 
        x"ce", x"ce", x"cf", x"ce", x"ce", x"cd", x"ca", x"da", x"dc", x"cf", x"d1", x"d3", x"d3", x"d3", x"ca", 
        x"ab", x"67", x"5f", x"5d", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5f", x"61", x"5e", x"5e", x"64", x"9b", x"db", x"f0", x"fb", x"f8", x"f6", 
        x"fa", x"fb", x"f9", x"f6", x"eb", x"c0", x"86", x"60", x"5b", x"5a", x"5d", x"5d", x"5e", x"5f", x"5f", 
        x"5d", x"5c", x"5c", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"60", x"5f", x"5a", x"5a", x"65", x"a0", 
        x"e4", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f3", x"f0", x"ee", 
        x"ef", x"ed", x"e3", x"d8", x"d3", x"db", x"e0", x"d5", x"b1", x"86", x"75", x"75", x"7b", x"7f", x"7f", 
        x"80", x"82", x"80", x"81", x"84", x"84", x"81", x"7d", x"7e", x"80", x"7e", x"7f", x"80", x"7e", x"7d", 
        x"7d", x"7e", x"7e", x"7f", x"80", x"80", x"7f", x"7f", x"7f", x"7e", x"7f", x"7e", x"7e", x"7e", x"7f", 
        x"7e", x"7c", x"7d", x"7e", x"7e", x"7f", x"7e", x"7d", x"7e", x"80", x"7e", x"7d", x"7f", x"7f", x"7e", 
        x"7e", x"7e", x"7d", x"7e", x"7c", x"7f", x"82", x"7e", x"7c", x"7f", x"7d", x"7c", x"7d", x"7d", x"7c", 
        x"7c", x"7c", x"7d", x"7e", x"7f", x"7f", x"7e", x"7c", x"7d", x"7e", x"7d", x"7d", x"7d", x"7c", x"7d", 
        x"7c", x"7d", x"7e", x"7f", x"7d", x"7c", x"7d", x"7f", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", 
        x"7e", x"7c", x"7c", x"7b", x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", x"7e", x"7b", x"7a", x"7e", x"7e", 
        x"7b", x"7b", x"7c", x"7d", x"7c", x"7d", x"7c", x"79", x"7b", x"7c", x"7d", x"7c", x"7b", x"7c", x"7d", 
        x"7b", x"7c", x"7d", x"7c", x"7b", x"7c", x"7c", x"7c", x"7d", x"7d", x"7c", x"7c", x"7c", x"7e", x"7d", 
        x"7f", x"7d", x"7b", x"7d", x"7c", x"7b", x"7c", x"7c", x"7a", x"7b", x"7c", x"7b", x"79", x"7a", x"7b", 
        x"7d", x"7a", x"7b", x"7b", x"7a", x"7b", x"78", x"78", x"7b", x"7d", x"7a", x"77", x"79", x"78", x"7a", 
        x"7a", x"79", x"7a", x"79", x"7a", x"7a", x"78", x"77", x"78", x"7a", x"7b", x"7c", x"7a", x"78", x"77", 
        x"77", x"78", x"78", x"78", x"78", x"78", x"79", x"78", x"78", x"77", x"78", x"78", x"77", x"78", x"7a", 
        x"77", x"74", x"75", x"75", x"76", x"77", x"78", x"79", x"78", x"78", x"77", x"78", x"76", x"77", x"77", 
        x"75", x"76", x"74", x"76", x"75", x"74", x"78", x"77", x"76", x"76", x"78", x"78", x"77", x"79", x"78", 
        x"75", x"76", x"75", x"74", x"75", x"77", x"75", x"75", x"76", x"76", x"77", x"77", x"76", x"76", x"76", 
        x"75", x"73", x"73", x"74", x"77", x"78", x"76", x"74", x"77", x"74", x"71", x"73", x"75", x"74", x"71", 
        x"75", x"78", x"78", x"75", x"75", x"77", x"77", x"76", x"76", x"76", x"75", x"74", x"75", x"76", x"75", 
        x"72", x"73", x"73", x"75", x"77", x"78", x"79", x"77", x"77", x"76", x"76", x"76", x"75", x"75", x"77", 
        x"77", x"77", x"77", x"76", x"75", x"74", x"72", x"72", x"76", x"76", x"76", x"78", x"76", x"77", x"77", 
        x"73", x"75", x"75", x"74", x"73", x"74", x"75", x"72", x"70", x"73", x"74", x"72", x"74", x"73", x"74", 
        x"73", x"72", x"72", x"72", x"70", x"71", x"73", x"74", x"73", x"73", x"74", x"73", x"73", x"71", x"72", 
        x"73", x"74", x"74", x"71", x"73", x"73", x"73", x"72", x"71", x"73", x"75", x"76", x"76", x"73", x"71", 
        x"73", x"74", x"74", x"73", x"74", x"72", x"70", x"73", x"74", x"73", x"76", x"76", x"73", x"73", x"75", 
        x"75", x"74", x"74", x"73", x"76", x"75", x"74", x"75", x"76", x"74", x"74", x"75", x"73", x"74", x"76", 
        x"74", x"75", x"74", x"77", x"76", x"74", x"77", x"76", x"75", x"76", x"74", x"74", x"73", x"72", x"73", 
        x"74", x"75", x"75", x"77", x"75", x"73", x"74", x"77", x"77", x"75", x"75", x"78", x"78", x"78", x"79", 
        x"78", x"76", x"76", x"76", x"76", x"76", x"77", x"78", x"76", x"74", x"76", x"77", x"76", x"74", x"76", 
        x"78", x"78", x"77", x"76", x"76", x"77", x"79", x"7a", x"79", x"78", x"77", x"76", x"77", x"77", x"77", 
        x"79", x"7a", x"7a", x"79", x"79", x"79", x"79", x"77", x"79", x"7b", x"7a", x"79", x"79", x"7b", x"76", 
        x"83", x"d4", x"d5", x"d2", x"d4", x"d4", x"dd", x"d5", x"cd", x"cf", x"cf", x"cd", x"cf", x"d2", x"d1", 
        x"cd", x"d1", x"cf", x"b2", x"93", x"a7", x"c8", x"d0", x"cd", x"ce", x"cf", x"cd", x"d1", x"d0", x"ce", 
        x"ce", x"ce", x"ce", x"cd", x"ce", x"cf", x"cf", x"ce", x"ce", x"cd", x"cd", x"ce", x"d0", x"d0", x"ce", 
        x"ce", x"cf", x"cf", x"cf", x"ce", x"cd", x"ca", x"d9", x"dc", x"d0", x"d1", x"d2", x"d4", x"d4", x"ca", 
        x"aa", x"67", x"5f", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5c", x"5f", x"5d", x"61", x"5b", x"72", x"bd", x"e7", x"f7", x"fa", x"f8", 
        x"f9", x"fb", x"f9", x"f7", x"f8", x"f2", x"cf", x"98", x"6c", x"5d", x"5c", x"5d", x"5c", x"5d", x"5e", 
        x"5d", x"5c", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5e", x"5c", x"5c", x"64", x"9a", 
        x"e4", x"f0", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ed", x"ee", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"ed", x"ef", x"f1", x"ef", x"e9", x"db", x"d5", x"db", x"e1", x"db", x"bc", x"91", x"77", x"76", x"78", 
        x"7e", x"80", x"80", x"80", x"7f", x"81", x"83", x"82", x"7f", x"7f", x"7f", x"7f", x"81", x"80", x"7e", 
        x"7e", x"7f", x"7e", x"80", x"80", x"7f", x"7e", x"7f", x"7f", x"80", x"7f", x"7f", x"7f", x"7f", x"80", 
        x"7f", x"7f", x"7d", x"7d", x"7e", x"7e", x"7d", x"7c", x"7e", x"7f", x"7d", x"7c", x"7f", x"80", x"7e", 
        x"7d", x"7d", x"7c", x"7c", x"7a", x"7c", x"7e", x"7b", x"7b", x"7d", x"7c", x"7c", x"7e", x"7f", x"7e", 
        x"7d", x"7e", x"7e", x"7d", x"7d", x"7d", x"7e", x"7e", x"7d", x"7d", x"7e", x"7e", x"7e", x"7d", x"7d", 
        x"7c", x"7b", x"7c", x"7c", x"7b", x"7a", x"7b", x"7d", x"7d", x"7c", x"7c", x"7b", x"7b", x"7a", x"7b", 
        x"7e", x"7e", x"7c", x"7b", x"7c", x"7d", x"7e", x"7d", x"7d", x"7e", x"7d", x"7b", x"7b", x"7e", x"7f", 
        x"7d", x"7c", x"7c", x"7c", x"7a", x"7b", x"7b", x"7a", x"7a", x"7b", x"7c", x"7c", x"7c", x"7b", x"79", 
        x"79", x"7a", x"7a", x"7a", x"79", x"79", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7e", x"7d", 
        x"7f", x"7d", x"7a", x"7b", x"7a", x"79", x"7d", x"7f", x"7c", x"7a", x"7b", x"7b", x"7b", x"7a", x"7a", 
        x"7c", x"7b", x"7c", x"7b", x"7a", x"7b", x"79", x"7a", x"7c", x"7d", x"79", x"78", x"7c", x"7b", x"7a", 
        x"79", x"78", x"79", x"7a", x"7b", x"7a", x"78", x"77", x"78", x"79", x"7a", x"7a", x"7a", x"79", x"79", 
        x"79", x"78", x"77", x"78", x"78", x"78", x"78", x"78", x"77", x"77", x"78", x"78", x"77", x"79", x"7b", 
        x"77", x"74", x"76", x"76", x"77", x"78", x"78", x"79", x"79", x"79", x"79", x"7a", x"77", x"78", x"78", 
        x"76", x"76", x"73", x"76", x"76", x"75", x"78", x"77", x"76", x"78", x"7a", x"78", x"77", x"78", x"77", 
        x"74", x"74", x"75", x"74", x"75", x"76", x"74", x"75", x"76", x"76", x"76", x"76", x"76", x"76", x"77", 
        x"76", x"73", x"75", x"76", x"76", x"75", x"75", x"76", x"77", x"74", x"70", x"73", x"76", x"76", x"74", 
        x"75", x"78", x"78", x"76", x"76", x"78", x"76", x"75", x"77", x"78", x"77", x"76", x"76", x"76", x"76", 
        x"75", x"74", x"73", x"75", x"76", x"77", x"77", x"77", x"77", x"77", x"76", x"76", x"76", x"76", x"77", 
        x"77", x"78", x"77", x"76", x"75", x"74", x"72", x"72", x"75", x"76", x"75", x"78", x"76", x"75", x"75", 
        x"71", x"73", x"75", x"75", x"75", x"75", x"77", x"74", x"71", x"73", x"73", x"71", x"72", x"71", x"73", 
        x"74", x"73", x"74", x"73", x"71", x"72", x"73", x"73", x"73", x"73", x"73", x"75", x"74", x"74", x"72", 
        x"74", x"75", x"75", x"72", x"73", x"72", x"74", x"72", x"72", x"74", x"75", x"77", x"76", x"77", x"74", 
        x"73", x"75", x"74", x"71", x"73", x"73", x"70", x"73", x"75", x"74", x"75", x"75", x"75", x"75", x"74", 
        x"73", x"74", x"76", x"74", x"76", x"76", x"75", x"77", x"77", x"74", x"73", x"74", x"74", x"75", x"77", 
        x"74", x"74", x"74", x"76", x"76", x"73", x"75", x"75", x"73", x"76", x"74", x"74", x"74", x"72", x"72", 
        x"74", x"74", x"74", x"76", x"75", x"74", x"76", x"78", x"78", x"75", x"73", x"73", x"72", x"72", x"72", 
        x"73", x"75", x"76", x"77", x"77", x"77", x"77", x"77", x"76", x"75", x"75", x"79", x"78", x"74", x"74", 
        x"77", x"78", x"79", x"79", x"77", x"77", x"78", x"79", x"78", x"77", x"78", x"78", x"76", x"77", x"79", 
        x"79", x"79", x"7a", x"79", x"79", x"7a", x"7b", x"79", x"7a", x"7d", x"7c", x"7a", x"78", x"7b", x"76", 
        x"81", x"d3", x"d5", x"d2", x"d4", x"d5", x"dd", x"d5", x"ce", x"cf", x"ce", x"cf", x"d0", x"ce", x"d3", 
        x"d5", x"c4", x"99", x"91", x"b9", x"cf", x"ca", x"cc", x"ce", x"ce", x"ce", x"cb", x"cb", x"ce", x"cf", 
        x"ce", x"cd", x"cd", x"ce", x"ce", x"cf", x"cf", x"ce", x"ce", x"ce", x"ce", x"ce", x"cf", x"d0", x"d0", 
        x"d0", x"d0", x"d1", x"d1", x"d0", x"cf", x"cc", x"db", x"de", x"d3", x"d4", x"d4", x"d5", x"d4", x"cb", 
        x"aa", x"67", x"5f", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5f", x"5e", x"5d", x"5d", x"5e", x"5f", x"8e", x"d3", x"f6", x"f8", x"f8", 
        x"fb", x"fa", x"f9", x"f9", x"f8", x"fa", x"f7", x"e8", x"bc", x"8d", x"6d", x"5f", x"5c", x"5d", x"60", 
        x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5d", x"5e", x"5e", x"5f", x"63", x"93", 
        x"e2", x"f1", x"ee", x"ef", x"ef", x"ed", x"ec", x"ed", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"ed", x"eb", x"e3", x"d4", x"d3", x"df", x"e0", x"c6", x"9d", x"7b", 
        x"74", x"7d", x"81", x"80", x"80", x"81", x"81", x"81", x"81", x"82", x"81", x"80", x"81", x"80", x"7f", 
        x"80", x"80", x"7e", x"7e", x"7d", x"7c", x"7c", x"7c", x"7d", x"7e", x"7e", x"7f", x"7f", x"80", x"80", 
        x"80", x"7f", x"7f", x"7f", x"80", x"80", x"7f", x"7f", x"80", x"80", x"7f", x"7d", x"7d", x"7d", x"7d", 
        x"7d", x"7e", x"7d", x"80", x"7f", x"7e", x"7e", x"7c", x"7f", x"7c", x"7c", x"7d", x"7f", x"80", x"80", 
        x"7e", x"7e", x"7e", x"7d", x"7c", x"7c", x"7d", x"7f", x"7d", x"7d", x"7d", x"7e", x"7f", x"7e", x"7d", 
        x"7c", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7d", x"7b", x"7b", x"7c", x"7c", x"7c", x"7c", x"7c", 
        x"7d", x"7e", x"7e", x"7f", x"7e", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7d", x"7e", x"7f", 
        x"7f", x"7e", x"7f", x"7e", x"7c", x"7d", x"7d", x"7b", x"7b", x"7b", x"7b", x"7c", x"7d", x"7b", x"7a", 
        x"7b", x"7c", x"7c", x"7c", x"7b", x"7a", x"7a", x"7b", x"7b", x"7c", x"7b", x"7b", x"7a", x"7d", x"7b", 
        x"7c", x"7c", x"7b", x"7c", x"7b", x"7b", x"7d", x"7e", x"7c", x"7b", x"7c", x"7b", x"7d", x"7b", x"78", 
        x"7a", x"7b", x"7e", x"7d", x"79", x"7b", x"7c", x"7c", x"7b", x"7b", x"79", x"79", x"7c", x"7c", x"7a", 
        x"7b", x"7b", x"7b", x"7c", x"79", x"79", x"7b", x"7c", x"7b", x"79", x"77", x"79", x"7a", x"7a", x"7a", 
        x"79", x"79", x"79", x"79", x"79", x"78", x"78", x"77", x"77", x"77", x"78", x"78", x"78", x"7a", x"79", 
        x"77", x"77", x"78", x"79", x"79", x"78", x"78", x"78", x"79", x"78", x"78", x"79", x"78", x"78", x"79", 
        x"78", x"79", x"77", x"78", x"76", x"73", x"76", x"77", x"77", x"79", x"78", x"77", x"77", x"78", x"77", 
        x"77", x"76", x"75", x"74", x"76", x"75", x"74", x"75", x"76", x"75", x"76", x"76", x"76", x"77", x"78", 
        x"77", x"77", x"77", x"77", x"76", x"75", x"75", x"76", x"77", x"76", x"75", x"75", x"77", x"77", x"76", 
        x"75", x"77", x"78", x"76", x"77", x"78", x"76", x"74", x"75", x"77", x"77", x"76", x"75", x"76", x"76", 
        x"77", x"76", x"75", x"76", x"78", x"78", x"77", x"77", x"77", x"77", x"77", x"78", x"78", x"78", x"77", 
        x"77", x"77", x"78", x"77", x"76", x"76", x"76", x"73", x"76", x"77", x"75", x"76", x"77", x"76", x"74", 
        x"74", x"74", x"76", x"76", x"75", x"75", x"74", x"75", x"74", x"74", x"74", x"72", x"73", x"72", x"73", 
        x"73", x"72", x"75", x"75", x"73", x"75", x"75", x"72", x"73", x"74", x"72", x"75", x"75", x"74", x"75", 
        x"74", x"73", x"75", x"73", x"73", x"71", x"75", x"74", x"76", x"74", x"74", x"76", x"75", x"78", x"77", 
        x"75", x"76", x"75", x"73", x"74", x"75", x"72", x"74", x"76", x"75", x"73", x"73", x"75", x"73", x"74", 
        x"75", x"77", x"77", x"74", x"75", x"77", x"75", x"75", x"74", x"72", x"72", x"75", x"74", x"73", x"75", 
        x"72", x"73", x"74", x"74", x"76", x"73", x"75", x"74", x"73", x"76", x"76", x"76", x"76", x"73", x"71", 
        x"74", x"73", x"73", x"75", x"76", x"76", x"77", x"79", x"78", x"75", x"78", x"7a", x"78", x"76", x"74", 
        x"76", x"7a", x"79", x"77", x"77", x"77", x"77", x"77", x"76", x"75", x"77", x"7a", x"79", x"75", x"74", 
        x"75", x"75", x"7a", x"7b", x"79", x"76", x"76", x"77", x"76", x"77", x"79", x"7a", x"78", x"79", x"7b", 
        x"7a", x"79", x"7a", x"7b", x"79", x"7a", x"7d", x"7c", x"7b", x"7c", x"7c", x"7c", x"77", x"7b", x"78", 
        x"81", x"d2", x"d4", x"d2", x"d5", x"d6", x"dd", x"d5", x"cc", x"cc", x"cf", x"cc", x"d1", x"d4", x"ca", 
        x"ad", x"95", x"a6", x"cd", x"d4", x"cb", x"cc", x"cb", x"cd", x"cb", x"cc", x"cd", x"ce", x"ce", x"cb", 
        x"cd", x"cc", x"cc", x"ce", x"cf", x"d0", x"cf", x"ce", x"ce", x"ce", x"ce", x"cf", x"cf", x"cf", x"d0", 
        x"d0", x"d1", x"d1", x"d1", x"d0", x"cf", x"cc", x"d8", x"db", x"d3", x"d4", x"d2", x"d1", x"d3", x"cb", 
        x"ab", x"66", x"5f", x"5c", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5f", x"5a", x"5f", x"5c", x"62", x"5d", x"5f", x"a4", x"e4", x"f6", x"f5", 
        x"f8", x"fb", x"fb", x"fb", x"f9", x"fa", x"fc", x"fa", x"f9", x"e7", x"ba", x"80", x"68", x"59", x"5c", 
        x"60", x"60", x"60", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"5f", x"61", x"60", x"5f", x"60", x"8c", 
        x"dd", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ed", x"ed", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", 
        x"f0", x"ee", x"ef", x"f2", x"f3", x"f0", x"ee", x"f0", x"f0", x"e0", x"d5", x"d5", x"df", x"e6", x"db", 
        x"ab", x"84", x"79", x"79", x"79", x"80", x"83", x"80", x"7f", x"81", x"82", x"80", x"81", x"81", x"81", 
        x"80", x"80", x"7f", x"7f", x"7f", x"7e", x"7e", x"7e", x"7f", x"80", x"7f", x"7f", x"81", x"81", x"80", 
        x"80", x"80", x"7f", x"7e", x"7f", x"7e", x"7e", x"7f", x"7f", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", 
        x"7e", x"7e", x"7f", x"83", x"81", x"81", x"80", x"7f", x"82", x"7e", x"7d", x"7e", x"7f", x"81", x"81", 
        x"7e", x"7c", x"7c", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7d", x"7e", x"7f", x"7f", x"7e", 
        x"7e", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7e", x"7c", x"7d", x"7d", x"7e", x"7e", x"7f", x"80", 
        x"7e", x"7f", x"7c", x"7d", x"7b", x"7d", x"7f", x"7e", x"7e", x"7c", x"7c", x"7e", x"7f", x"7d", x"7c", 
        x"7c", x"7b", x"7d", x"7e", x"7d", x"7d", x"7e", x"7d", x"7d", x"7b", x"7b", x"7c", x"7d", x"7d", x"7d", 
        x"80", x"80", x"7e", x"7e", x"7e", x"7c", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7e", x"7c", 
        x"7c", x"7d", x"7b", x"7d", x"7c", x"7c", x"7c", x"7a", x"7a", x"7d", x"7f", x"7c", x"7d", x"7c", x"79", 
        x"7b", x"7c", x"7e", x"7e", x"79", x"7c", x"7d", x"7d", x"7b", x"79", x"79", x"7a", x"79", x"7b", x"7a", 
        x"7d", x"7e", x"7c", x"7d", x"79", x"79", x"7a", x"7b", x"7b", x"7a", x"7a", x"7b", x"7c", x"7b", x"79", 
        x"78", x"79", x"7c", x"7b", x"79", x"78", x"78", x"78", x"78", x"78", x"7a", x"78", x"78", x"7a", x"78", 
        x"77", x"79", x"7a", x"7a", x"78", x"78", x"77", x"78", x"78", x"79", x"7a", x"7b", x"79", x"79", x"79", 
        x"77", x"78", x"76", x"7a", x"78", x"76", x"78", x"77", x"75", x"77", x"75", x"75", x"78", x"78", x"79", 
        x"7b", x"78", x"76", x"75", x"78", x"75", x"75", x"75", x"77", x"76", x"76", x"76", x"77", x"77", x"77", 
        x"78", x"7a", x"77", x"76", x"77", x"78", x"77", x"76", x"79", x"79", x"78", x"77", x"77", x"77", x"76", 
        x"75", x"77", x"78", x"76", x"76", x"79", x"78", x"76", x"75", x"76", x"76", x"75", x"75", x"76", x"76", 
        x"76", x"76", x"76", x"78", x"79", x"79", x"79", x"77", x"77", x"77", x"78", x"78", x"79", x"78", x"76", 
        x"76", x"77", x"77", x"77", x"78", x"78", x"79", x"76", x"78", x"78", x"76", x"78", x"78", x"77", x"77", 
        x"76", x"75", x"76", x"76", x"76", x"74", x"73", x"74", x"73", x"74", x"74", x"72", x"74", x"74", x"75", 
        x"74", x"73", x"76", x"76", x"72", x"74", x"75", x"75", x"76", x"75", x"71", x"73", x"71", x"72", x"77", 
        x"74", x"71", x"73", x"73", x"73", x"71", x"73", x"73", x"77", x"75", x"74", x"78", x"76", x"75", x"75", 
        x"76", x"76", x"76", x"74", x"73", x"73", x"73", x"73", x"75", x"77", x"73", x"73", x"76", x"74", x"76", 
        x"75", x"75", x"76", x"75", x"76", x"75", x"73", x"74", x"74", x"73", x"74", x"77", x"75", x"72", x"74", 
        x"72", x"74", x"76", x"75", x"75", x"73", x"76", x"76", x"76", x"79", x"79", x"76", x"76", x"72", x"71", 
        x"75", x"74", x"74", x"77", x"77", x"77", x"78", x"77", x"77", x"77", x"78", x"78", x"77", x"77", x"75", 
        x"76", x"79", x"76", x"75", x"77", x"78", x"78", x"77", x"75", x"74", x"77", x"78", x"77", x"76", x"78", 
        x"77", x"74", x"77", x"7a", x"78", x"75", x"76", x"79", x"79", x"79", x"79", x"7a", x"7b", x"7c", x"7a", 
        x"7b", x"7b", x"7c", x"7c", x"7a", x"7b", x"7e", x"7c", x"7a", x"79", x"7c", x"7d", x"77", x"7c", x"7a", 
        x"83", x"d1", x"d3", x"d2", x"d5", x"d6", x"dd", x"d5", x"cb", x"cd", x"cf", x"d1", x"d3", x"b9", x"9b", 
        x"9c", x"bc", x"d1", x"cd", x"cb", x"c9", x"cb", x"cf", x"d0", x"cc", x"cd", x"ce", x"ca", x"cc", x"ce", 
        x"cc", x"cb", x"cb", x"cd", x"cf", x"d0", x"ce", x"ce", x"ce", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", 
        x"cf", x"d0", x"d0", x"d0", x"d0", x"cf", x"cc", x"d7", x"da", x"d3", x"d6", x"d2", x"cf", x"d2", x"ca", 
        x"ab", x"67", x"5f", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5c", x"5c", x"5f", x"5c", x"60", x"60", x"5d", x"70", x"a5", x"e1", x"f7", 
        x"f9", x"fa", x"fc", x"f9", x"fa", x"fa", x"f9", x"fb", x"fa", x"f9", x"ed", x"cc", x"a7", x"87", x"71", 
        x"64", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"5f", x"5a", x"5a", x"60", x"8c", 
        x"dd", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f1", x"ef", x"e7", x"da", x"d5", x"d7", 
        x"db", x"d5", x"bb", x"96", x"7e", x"73", x"75", x"80", x"82", x"80", x"80", x"80", x"80", x"81", x"82", 
        x"81", x"7f", x"7f", x"80", x"80", x"80", x"80", x"80", x"81", x"82", x"80", x"80", x"81", x"82", x"80", 
        x"7f", x"80", x"80", x"80", x"7f", x"7d", x"7d", x"80", x"80", x"7e", x"7f", x"81", x"81", x"80", x"81", 
        x"80", x"7e", x"7f", x"80", x"7d", x"7e", x"80", x"7e", x"7f", x"80", x"80", x"7e", x"7d", x"7f", x"80", 
        x"7e", x"7c", x"7c", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7d", x"7e", x"7f", x"7f", x"7f", 
        x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", 
        x"7d", x"7e", x"7c", x"7d", x"7b", x"7d", x"7f", x"7d", x"7e", x"7e", x"7d", x"7e", x"7f", x"7d", x"7d", 
        x"7d", x"7c", x"7e", x"7d", x"7c", x"7d", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7c", x"7b", x"7b", 
        x"7e", x"7e", x"7b", x"7b", x"7b", x"79", x"7c", x"7d", x"7d", x"7e", x"7d", x"7d", x"7d", x"7f", x"7d", 
        x"7e", x"7e", x"7d", x"7f", x"7e", x"7c", x"7d", x"7c", x"7a", x"7c", x"7f", x"7d", x"7c", x"7b", x"7c", 
        x"7e", x"7b", x"7c", x"7d", x"7c", x"7d", x"7d", x"7b", x"7b", x"7a", x"79", x"78", x"7a", x"7b", x"79", 
        x"7b", x"7c", x"7a", x"7c", x"7a", x"79", x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", 
        x"7a", x"7a", x"7c", x"7a", x"79", x"78", x"78", x"78", x"79", x"7a", x"7a", x"77", x"78", x"7b", x"79", 
        x"77", x"7a", x"79", x"78", x"78", x"78", x"78", x"79", x"7a", x"7a", x"7b", x"7b", x"79", x"79", x"7a", 
        x"78", x"78", x"78", x"7b", x"79", x"77", x"78", x"77", x"76", x"77", x"75", x"78", x"7a", x"77", x"77", 
        x"79", x"77", x"76", x"76", x"79", x"75", x"75", x"76", x"79", x"79", x"79", x"79", x"78", x"78", x"78", 
        x"77", x"78", x"78", x"79", x"79", x"79", x"79", x"78", x"78", x"77", x"76", x"77", x"78", x"79", x"78", 
        x"75", x"77", x"78", x"76", x"75", x"79", x"7b", x"79", x"78", x"78", x"78", x"77", x"77", x"79", x"79", 
        x"77", x"78", x"78", x"76", x"76", x"77", x"78", x"78", x"78", x"78", x"78", x"78", x"78", x"78", x"77", 
        x"77", x"77", x"77", x"77", x"77", x"77", x"76", x"77", x"7a", x"78", x"77", x"7a", x"77", x"77", x"77", 
        x"75", x"76", x"75", x"77", x"76", x"73", x"74", x"75", x"73", x"74", x"74", x"72", x"74", x"74", x"75", 
        x"75", x"75", x"76", x"74", x"72", x"74", x"74", x"74", x"75", x"74", x"73", x"74", x"73", x"75", x"77", 
        x"73", x"71", x"73", x"72", x"73", x"73", x"73", x"72", x"74", x"74", x"74", x"76", x"75", x"73", x"73", 
        x"74", x"75", x"75", x"74", x"75", x"74", x"75", x"74", x"76", x"79", x"74", x"74", x"78", x"77", x"77", 
        x"75", x"74", x"74", x"74", x"75", x"74", x"73", x"72", x"74", x"75", x"75", x"76", x"76", x"76", x"77", 
        x"75", x"75", x"76", x"75", x"75", x"74", x"75", x"75", x"76", x"78", x"78", x"73", x"75", x"74", x"74", 
        x"78", x"76", x"76", x"76", x"75", x"75", x"77", x"76", x"76", x"77", x"78", x"76", x"76", x"79", x"78", 
        x"78", x"78", x"77", x"76", x"78", x"78", x"78", x"77", x"76", x"76", x"78", x"78", x"76", x"75", x"78", 
        x"79", x"75", x"77", x"79", x"7a", x"77", x"78", x"7c", x"7c", x"7a", x"78", x"79", x"7b", x"7b", x"7a", 
        x"7c", x"7b", x"7a", x"79", x"79", x"7a", x"7b", x"7b", x"7b", x"7a", x"7b", x"7b", x"77", x"7b", x"79", 
        x"83", x"d1", x"d5", x"d3", x"d6", x"d4", x"dd", x"d6", x"c9", x"d4", x"d5", x"ce", x"ad", x"91", x"a4", 
        x"c8", x"d0", x"cd", x"cc", x"c9", x"cc", x"cf", x"cf", x"cf", x"cc", x"cb", x"cd", x"cf", x"cd", x"cb", 
        x"ce", x"cd", x"cb", x"cc", x"ce", x"d0", x"d0", x"ce", x"ce", x"ce", x"ce", x"ce", x"ce", x"ce", x"cf", 
        x"cf", x"d0", x"d0", x"d0", x"cf", x"ce", x"cc", x"d7", x"da", x"d3", x"d7", x"d2", x"ce", x"d2", x"ca", 
        x"ac", x"69", x"5d", x"5c", x"5e", x"5f", x"5d", x"5c", x"5e", x"5d", x"5e", x"5c", x"5b", x"5c", x"5f", 
        x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5c", x"5d", x"5f", x"60", x"5b", x"6a", x"a3", x"de", 
        x"f7", x"f8", x"f9", x"fa", x"fa", x"f9", x"f9", x"fa", x"fa", x"fb", x"f8", x"ed", x"dc", x"c9", x"b2", 
        x"96", x"7d", x"67", x"5d", x"5c", x"5d", x"5d", x"5d", x"5d", x"5e", x"5c", x"5c", x"5c", x"5c", x"5d", 
        x"5e", x"5e", x"5f", x"5e", x"5d", x"5b", x"5b", x"5c", x"5a", x"5c", x"5e", x"69", x"7a", x"8b", x"a8", 
        x"e3", x"f0", x"ee", x"ee", x"ef", x"ee", x"ed", x"ee", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"ef", 
        x"f1", x"f0", x"f0", x"f1", x"f0", x"ee", x"f0", x"f2", x"ed", x"ee", x"f0", x"f2", x"f0", x"e5", x"da", 
        x"d0", x"d4", x"df", x"df", x"c0", x"9e", x"7b", x"73", x"7a", x"80", x"7f", x"7f", x"81", x"82", x"80", 
        x"7f", x"7f", x"7f", x"80", x"7f", x"80", x"82", x"82", x"80", x"81", x"80", x"80", x"82", x"81", x"80", 
        x"80", x"81", x"80", x"80", x"80", x"7e", x"7e", x"80", x"80", x"7f", x"80", x"81", x"7f", x"80", x"81", 
        x"80", x"7f", x"7d", x"7e", x"7d", x"7e", x"80", x"7e", x"7e", x"82", x"81", x"7e", x"7d", x"7e", x"80", 
        x"7f", x"7d", x"7d", x"7e", x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", x"7e", x"7e", x"7d", x"7e", x"7d", 
        x"7e", x"7f", x"80", x"7f", x"7d", x"7d", x"7e", x"7f", x"7c", x"7c", x"7c", x"7c", x"7d", x"7e", x"7e", 
        x"7e", x"7d", x"7b", x"7d", x"7c", x"7c", x"7d", x"7e", x"7e", x"7e", x"7e", x"7d", x"7e", x"7d", x"7e", 
        x"7f", x"7e", x"7e", x"7e", x"7c", x"7d", x"7e", x"7e", x"7f", x"7f", x"7e", x"7d", x"7c", x"7b", x"7a", 
        x"7d", x"7d", x"7b", x"7c", x"7c", x"7a", x"7d", x"7e", x"7f", x"7d", x"7d", x"7d", x"7d", x"7c", x"7d", 
        x"7e", x"7f", x"80", x"7e", x"7d", x"7c", x"7e", x"7e", x"7b", x"7c", x"7e", x"7f", x"7d", x"79", x"7c", 
        x"7d", x"7b", x"7c", x"7b", x"7c", x"7c", x"7c", x"7b", x"7b", x"7c", x"76", x"76", x"7b", x"7b", x"79", 
        x"7a", x"7a", x"7a", x"7c", x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7a", x"7a", x"7a", x"7c", x"7b", 
        x"7a", x"79", x"79", x"78", x"78", x"78", x"78", x"79", x"79", x"79", x"79", x"78", x"79", x"7c", x"79", 
        x"78", x"7a", x"7a", x"78", x"79", x"79", x"78", x"79", x"7a", x"78", x"77", x"79", x"79", x"79", x"79", 
        x"79", x"7b", x"78", x"79", x"78", x"76", x"77", x"77", x"77", x"76", x"76", x"79", x"7a", x"78", x"77", 
        x"78", x"78", x"77", x"77", x"7b", x"78", x"78", x"79", x"79", x"79", x"7a", x"79", x"78", x"78", x"78", 
        x"77", x"76", x"76", x"77", x"79", x"78", x"78", x"78", x"76", x"76", x"76", x"77", x"78", x"78", x"77", 
        x"74", x"75", x"77", x"76", x"77", x"78", x"79", x"79", x"78", x"78", x"77", x"76", x"77", x"77", x"78", 
        x"78", x"78", x"78", x"76", x"76", x"76", x"77", x"79", x"77", x"76", x"77", x"77", x"78", x"78", x"78", 
        x"78", x"79", x"79", x"78", x"78", x"78", x"77", x"78", x"7a", x"76", x"77", x"7b", x"78", x"77", x"78", 
        x"73", x"75", x"76", x"77", x"76", x"71", x"74", x"74", x"73", x"73", x"72", x"72", x"72", x"71", x"72", 
        x"74", x"74", x"73", x"72", x"73", x"75", x"74", x"74", x"74", x"73", x"76", x"76", x"75", x"76", x"76", 
        x"74", x"74", x"74", x"74", x"75", x"76", x"75", x"73", x"72", x"73", x"74", x"74", x"73", x"72", x"72", 
        x"73", x"73", x"74", x"75", x"76", x"73", x"75", x"75", x"75", x"78", x"76", x"76", x"78", x"76", x"75", 
        x"75", x"76", x"75", x"74", x"74", x"75", x"74", x"73", x"74", x"77", x"76", x"73", x"75", x"79", x"79", 
        x"78", x"77", x"76", x"75", x"77", x"77", x"77", x"76", x"76", x"77", x"77", x"75", x"77", x"75", x"74", 
        x"78", x"77", x"77", x"78", x"76", x"75", x"77", x"78", x"77", x"77", x"77", x"77", x"78", x"7a", x"7b", 
        x"79", x"78", x"77", x"79", x"7a", x"79", x"78", x"79", x"7a", x"7b", x"76", x"77", x"75", x"74", x"77", 
        x"79", x"78", x"78", x"78", x"7b", x"78", x"78", x"7c", x"7b", x"79", x"7a", x"7a", x"7a", x"7a", x"7a", 
        x"7a", x"7a", x"78", x"78", x"7a", x"7b", x"7a", x"7a", x"7c", x"7d", x"7b", x"79", x"79", x"7a", x"77", 
        x"80", x"cc", x"d3", x"d2", x"d8", x"d8", x"de", x"d2", x"cc", x"d9", x"bf", x"93", x"99", x"bf", x"ce", 
        x"cb", x"cb", x"cb", x"cb", x"cc", x"cd", x"d0", x"cf", x"ce", x"ce", x"cd", x"cc", x"cc", x"ce", x"cf", 
        x"cf", x"cf", x"ce", x"cc", x"cd", x"ce", x"d0", x"cf", x"ce", x"cd", x"ce", x"cf", x"ce", x"ce", x"d0", 
        x"d0", x"d0", x"d0", x"d0", x"d0", x"ce", x"ca", x"d7", x"db", x"d2", x"d5", x"d2", x"ce", x"d1", x"c9", 
        x"af", x"6c", x"5d", x"5d", x"5e", x"60", x"5e", x"5d", x"5f", x"5e", x"5f", x"5e", x"5f", x"5d", x"5c", 
        x"5b", x"5d", x"60", x"60", x"5d", x"5d", x"5d", x"5c", x"5c", x"5e", x"5f", x"60", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5c", x"63", x"8b", 
        x"c9", x"f1", x"fa", x"fb", x"fa", x"f8", x"f9", x"fb", x"fb", x"fb", x"fb", x"fa", x"f4", x"ef", x"e7", 
        x"d7", x"bd", x"94", x"6f", x"63", x"59", x"57", x"5a", x"5c", x"5d", x"5b", x"5b", x"5a", x"59", x"59", 
        x"5a", x"5c", x"5c", x"62", x"77", x"84", x"89", x"8b", x"87", x"93", x"ac", x"b3", x"a2", x"9c", x"b4", 
        x"e4", x"f0", x"f0", x"ee", x"ee", x"ef", x"f0", x"ee", x"ed", x"ee", x"f0", x"f1", x"ef", x"ed", x"ec", 
        x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", 
        x"eb", x"de", x"d3", x"d1", x"d8", x"de", x"d6", x"ae", x"87", x"73", x"71", x"7d", x"81", x"81", x"81", 
        x"83", x"83", x"83", x"82", x"81", x"82", x"83", x"80", x"7d", x"81", x"81", x"81", x"82", x"81", x"80", 
        x"82", x"80", x"7d", x"7d", x"7e", x"7f", x"80", x"80", x"7f", x"7f", x"7f", x"80", x"7f", x"81", x"81", 
        x"7e", x"7f", x"7e", x"7f", x"80", x"7f", x"7f", x"80", x"81", x"81", x"80", x"7f", x"7f", x"7f", x"7f", 
        x"7f", x"7d", x"7d", x"7e", x"7e", x"7c", x"7c", x"7c", x"7e", x"7e", x"7f", x"7d", x"7d", x"7e", x"7d", 
        x"7e", x"80", x"81", x"7f", x"7c", x"7b", x"7e", x"7f", x"7b", x"7c", x"7c", x"7d", x"7e", x"7f", x"7f", 
        x"7f", x"7c", x"7b", x"7d", x"7c", x"7b", x"7d", x"80", x"7c", x"7d", x"7e", x"7d", x"7d", x"7e", x"7c", 
        x"7c", x"7c", x"7c", x"7b", x"7b", x"7c", x"7c", x"7e", x"7f", x"7f", x"7d", x"7d", x"7d", x"7c", x"7a", 
        x"7d", x"7d", x"7b", x"7c", x"7d", x"7c", x"7c", x"7e", x"7f", x"7e", x"7c", x"7c", x"7c", x"79", x"7c", 
        x"7d", x"7e", x"7e", x"7a", x"7b", x"7c", x"7d", x"7e", x"7c", x"7c", x"7d", x"7e", x"7e", x"7b", x"7c", 
        x"7c", x"7d", x"7f", x"7c", x"7e", x"7c", x"7c", x"7b", x"7c", x"7e", x"78", x"78", x"79", x"7a", x"7b", 
        x"7b", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7b", x"7a", x"7a", x"79", x"79", x"79", x"7b", x"7b", 
        x"7c", x"7c", x"7b", x"78", x"78", x"78", x"78", x"7b", x"79", x"77", x"78", x"79", x"7b", x"7c", x"7a", 
        x"79", x"79", x"79", x"79", x"7c", x"7c", x"7a", x"7b", x"79", x"77", x"77", x"7a", x"7c", x"7b", x"79", 
        x"79", x"7a", x"76", x"76", x"78", x"77", x"76", x"76", x"76", x"76", x"78", x"78", x"77", x"77", x"78", 
        x"79", x"78", x"76", x"78", x"7a", x"79", x"79", x"7a", x"77", x"78", x"7b", x"7a", x"78", x"79", x"7b", 
        x"7a", x"79", x"75", x"75", x"77", x"78", x"78", x"7a", x"7b", x"7a", x"7a", x"79", x"78", x"78", x"77", 
        x"78", x"78", x"78", x"78", x"78", x"78", x"78", x"78", x"77", x"77", x"76", x"77", x"78", x"77", x"78", 
        x"79", x"79", x"78", x"78", x"78", x"78", x"79", x"78", x"76", x"74", x"75", x"76", x"77", x"77", x"79", 
        x"78", x"76", x"76", x"76", x"77", x"78", x"7a", x"78", x"78", x"76", x"77", x"78", x"79", x"78", x"79", 
        x"73", x"75", x"76", x"77", x"76", x"73", x"75", x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"72", 
        x"72", x"72", x"72", x"71", x"73", x"75", x"75", x"74", x"75", x"75", x"77", x"76", x"74", x"75", x"75", 
        x"75", x"75", x"75", x"75", x"75", x"75", x"74", x"74", x"74", x"75", x"76", x"74", x"73", x"73", x"73", 
        x"74", x"74", x"75", x"75", x"76", x"75", x"78", x"77", x"74", x"76", x"77", x"76", x"77", x"77", x"77", 
        x"75", x"74", x"74", x"74", x"75", x"75", x"76", x"75", x"76", x"78", x"77", x"74", x"74", x"77", x"77", 
        x"76", x"77", x"77", x"76", x"78", x"78", x"77", x"76", x"75", x"74", x"74", x"76", x"79", x"77", x"76", 
        x"78", x"77", x"77", x"78", x"78", x"78", x"78", x"78", x"78", x"77", x"77", x"78", x"7a", x"77", x"77", 
        x"79", x"79", x"78", x"78", x"79", x"78", x"77", x"78", x"7a", x"7b", x"77", x"78", x"77", x"76", x"77", 
        x"79", x"78", x"78", x"77", x"78", x"78", x"77", x"7b", x"79", x"79", x"7a", x"7a", x"7a", x"79", x"7a", 
        x"7a", x"79", x"78", x"79", x"7c", x"7d", x"7b", x"7b", x"7c", x"7c", x"7b", x"7a", x"7b", x"7c", x"78", 
        x"81", x"ce", x"d8", x"cf", x"d0", x"d3", x"dd", x"db", x"ca", x"a8", x"91", x"ae", x"c9", x"d0", x"cc", 
        x"c9", x"ca", x"cc", x"cd", x"cc", x"cd", x"ce", x"cd", x"ce", x"cf", x"ce", x"cd", x"cd", x"d0", x"d1", 
        x"d0", x"cf", x"ce", x"ce", x"ce", x"ce", x"ce", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", 
        x"d0", x"d0", x"d0", x"d0", x"cf", x"ce", x"cc", x"d8", x"dc", x"d2", x"d6", x"d3", x"d0", x"d1", x"c9", 
        x"b1", x"6e", x"5e", x"5c", x"5d", x"5d", x"5e", x"5e", x"5d", x"69", x"6f", x"62", x"5e", x"5e", x"5c", 
        x"5c", x"5d", x"5e", x"5e", x"5f", x"5f", x"5e", x"5d", x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"60", x"5f", x"5c", x"61", 
        x"7c", x"b4", x"e5", x"f5", x"f8", x"f7", x"f9", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fa", x"f7", 
        x"f1", x"eb", x"da", x"c7", x"b4", x"9e", x"8e", x"86", x"7e", x"76", x"7a", x"81", x"86", x"8b", x"8f", 
        x"96", x"9e", x"aa", x"b7", x"ce", x"d9", x"d8", x"d1", x"c3", x"b8", x"b2", x"ad", x"a2", x"a1", x"ac", 
        x"d5", x"e8", x"ee", x"ec", x"ec", x"ee", x"ee", x"ed", x"eb", x"ee", x"ed", x"ec", x"ee", x"f0", x"f0", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"f0", x"f2", x"ea", x"df", x"d2", x"c2", x"ce", x"dc", x"d3", x"b4", x"8d", x"76", x"75", x"7b", x"81", 
        x"82", x"81", x"83", x"84", x"82", x"7f", x"7e", x"81", x"83", x"7f", x"7f", x"82", x"82", x"81", x"80", 
        x"80", x"7e", x"7f", x"82", x"82", x"81", x"80", x"7f", x"7d", x"7d", x"7f", x"80", x"7f", x"80", x"81", 
        x"7e", x"7f", x"7f", x"7f", x"7f", x"7e", x"7e", x"80", x"82", x"7f", x"81", x"82", x"81", x"7f", x"7e", 
        x"7f", x"7f", x"7e", x"7e", x"7c", x"7c", x"7c", x"7e", x"7f", x"7e", x"7e", x"7d", x"7d", x"7f", x"7e", 
        x"80", x"81", x"80", x"7f", x"7d", x"7d", x"7f", x"7f", x"7b", x"7c", x"7d", x"7e", x"7e", x"7e", x"7e", 
        x"7d", x"7c", x"7c", x"7e", x"7e", x"7d", x"7e", x"7f", x"7c", x"7e", x"7f", x"7d", x"7d", x"7f", x"7d", 
        x"7d", x"7f", x"7f", x"7e", x"7d", x"7d", x"7d", x"7e", x"7f", x"7f", x"7e", x"7d", x"7d", x"7d", x"7c", 
        x"7e", x"7d", x"7b", x"7c", x"7d", x"7c", x"7a", x"7c", x"7e", x"7e", x"7e", x"7c", x"7c", x"7c", x"7e", 
        x"7d", x"7d", x"7e", x"7d", x"7f", x"7c", x"7c", x"7d", x"7c", x"7b", x"7b", x"7d", x"7f", x"7d", x"7e", 
        x"7e", x"7f", x"81", x"7e", x"80", x"7e", x"7d", x"7b", x"7c", x"7d", x"7c", x"7c", x"7a", x"7a", x"7c", 
        x"7c", x"7c", x"7b", x"7b", x"7d", x"7c", x"7c", x"7b", x"7a", x"7a", x"7a", x"78", x"78", x"7a", x"7a", 
        x"7c", x"7d", x"7d", x"79", x"79", x"7a", x"79", x"7a", x"78", x"78", x"79", x"79", x"7b", x"7b", x"7a", 
        x"79", x"7a", x"7a", x"7a", x"7b", x"7a", x"79", x"7b", x"7a", x"78", x"7b", x"7c", x"7c", x"7c", x"7a", 
        x"79", x"78", x"79", x"79", x"77", x"76", x"75", x"76", x"77", x"79", x"79", x"78", x"78", x"77", x"77", 
        x"78", x"77", x"77", x"78", x"79", x"7a", x"79", x"79", x"78", x"79", x"7b", x"7a", x"79", x"79", x"7b", 
        x"7a", x"7b", x"77", x"77", x"78", x"79", x"7a", x"7b", x"7a", x"78", x"76", x"77", x"79", x"7a", x"79", 
        x"78", x"79", x"7a", x"79", x"77", x"77", x"77", x"7a", x"79", x"79", x"77", x"77", x"77", x"74", x"76", 
        x"77", x"77", x"77", x"77", x"77", x"77", x"77", x"78", x"76", x"75", x"75", x"76", x"76", x"76", x"78", 
        x"78", x"77", x"77", x"77", x"77", x"77", x"78", x"77", x"78", x"77", x"77", x"77", x"77", x"76", x"78", 
        x"74", x"75", x"75", x"76", x"76", x"75", x"77", x"75", x"74", x"74", x"74", x"75", x"75", x"75", x"74", 
        x"73", x"73", x"73", x"73", x"75", x"76", x"75", x"75", x"76", x"75", x"78", x"76", x"73", x"75", x"74", 
        x"74", x"73", x"73", x"73", x"74", x"74", x"75", x"75", x"76", x"77", x"76", x"75", x"74", x"74", x"74", 
        x"75", x"76", x"76", x"75", x"75", x"75", x"78", x"77", x"75", x"76", x"76", x"75", x"77", x"78", x"78", 
        x"77", x"74", x"72", x"73", x"73", x"74", x"75", x"75", x"75", x"76", x"75", x"73", x"75", x"78", x"77", 
        x"76", x"76", x"76", x"74", x"74", x"75", x"75", x"76", x"76", x"75", x"74", x"75", x"77", x"78", x"79", 
        x"7a", x"77", x"75", x"74", x"76", x"78", x"77", x"77", x"79", x"77", x"77", x"7a", x"79", x"76", x"75", 
        x"78", x"7a", x"79", x"79", x"79", x"79", x"78", x"78", x"7b", x"7b", x"76", x"76", x"78", x"79", x"7a", 
        x"7b", x"7a", x"79", x"77", x"77", x"78", x"78", x"7a", x"78", x"78", x"79", x"7a", x"7a", x"7a", x"7c", 
        x"7c", x"7a", x"78", x"79", x"7c", x"7e", x"7c", x"7d", x"7d", x"7b", x"7b", x"7b", x"7c", x"7d", x"78", 
        x"81", x"ce", x"d5", x"cf", x"d0", x"d6", x"e3", x"c9", x"89", x"93", x"c2", x"cd", x"cf", x"cd", x"c9", 
        x"c9", x"cb", x"cd", x"cd", x"cc", x"cd", x"ce", x"ce", x"cd", x"cc", x"cd", x"cf", x"d0", x"d0", x"d1", 
        x"d1", x"ce", x"cd", x"cd", x"ce", x"ce", x"ce", x"ce", x"cf", x"cf", x"ce", x"ce", x"cf", x"d1", x"d0", 
        x"d0", x"cf", x"cf", x"cf", x"cf", x"ce", x"cd", x"d9", x"dc", x"d1", x"d6", x"d4", x"d2", x"d2", x"cb", 
        x"b4", x"6f", x"5d", x"5c", x"5d", x"5b", x"5e", x"60", x"6a", x"9d", x"bc", x"9f", x"7b", x"62", x"5b", 
        x"5a", x"5e", x"60", x"5e", x"5f", x"61", x"5f", x"5e", x"5d", x"5e", x"5f", x"5f", x"5d", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"60", x"5e", x"5e", 
        x"5f", x"69", x"9a", x"d2", x"f3", x"f7", x"f8", x"f8", x"fa", x"fb", x"fb", x"fb", x"fa", x"f9", x"f8", 
        x"f8", x"fb", x"f9", x"f5", x"f0", x"ea", x"e5", x"e0", x"d9", x"d4", x"d6", x"dc", x"e2", x"e4", x"e6", 
        x"e8", x"ec", x"f0", x"f0", x"ee", x"e7", x"d8", x"cb", x"ba", x"b6", x"c6", x"be", x"9e", x"80", x"7f", 
        x"a0", x"ab", x"c5", x"dd", x"f0", x"f1", x"ec", x"ee", x"f2", x"ef", x"ee", x"ee", x"ed", x"ec", x"ed", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f1", x"f2", x"f0", 
        x"ec", x"ed", x"f0", x"f2", x"ed", x"e1", x"d6", x"ca", x"cd", x"dd", x"de", x"c6", x"9a", x"74", x"73", 
        x"7a", x"7f", x"83", x"83", x"83", x"82", x"80", x"7f", x"81", x"81", x"81", x"82", x"82", x"80", x"80", 
        x"7f", x"7e", x"80", x"81", x"81", x"81", x"80", x"7f", x"7e", x"7e", x"80", x"80", x"80", x"80", x"81", 
        x"7f", x"7f", x"7f", x"80", x"80", x"80", x"7f", x"7f", x"80", x"7f", x"81", x"82", x"82", x"80", x"7f", 
        x"80", x"7f", x"7f", x"7f", x"7d", x"7d", x"7d", x"80", x"80", x"7e", x"7e", x"7d", x"7d", x"7f", x"7e", 
        x"81", x"82", x"7f", x"7f", x"7f", x"7f", x"7f", x"7e", x"7d", x"7c", x"7c", x"7c", x"7d", x"7e", x"7f", 
        x"7d", x"7e", x"7f", x"80", x"7f", x"7e", x"80", x"7f", x"7d", x"7f", x"7e", x"7b", x"7e", x"80", x"7d", 
        x"7d", x"7f", x"80", x"7e", x"7d", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7f", 
        x"7f", x"7d", x"7c", x"7d", x"7d", x"7d", x"7b", x"7c", x"7e", x"7e", x"7e", x"7c", x"7c", x"7c", x"7e", 
        x"7c", x"7b", x"7c", x"7c", x"7f", x"7c", x"7b", x"7d", x"7c", x"7c", x"7b", x"7c", x"7f", x"7e", x"7d", 
        x"7d", x"7f", x"80", x"7e", x"7e", x"7e", x"7d", x"7c", x"7b", x"7b", x"79", x"79", x"7a", x"7c", x"7e", 
        x"7d", x"7d", x"7b", x"7a", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", x"7a", x"7b", x"7a", 
        x"7b", x"7b", x"7b", x"78", x"7a", x"7c", x"7a", x"7a", x"78", x"78", x"7c", x"7d", x"7a", x"78", x"77", 
        x"79", x"7c", x"7c", x"7b", x"7b", x"79", x"78", x"7b", x"7a", x"79", x"7c", x"7c", x"7a", x"7b", x"7a", 
        x"79", x"77", x"7b", x"7a", x"78", x"77", x"77", x"79", x"78", x"79", x"77", x"77", x"7a", x"7a", x"79", 
        x"78", x"78", x"7b", x"7b", x"7a", x"7c", x"7a", x"7a", x"7a", x"79", x"7a", x"79", x"77", x"77", x"77", 
        x"78", x"7a", x"78", x"77", x"78", x"78", x"78", x"7a", x"7a", x"79", x"77", x"79", x"7a", x"7b", x"7b", 
        x"77", x"77", x"7b", x"7a", x"77", x"76", x"76", x"79", x"78", x"78", x"77", x"78", x"79", x"76", x"77", 
        x"78", x"7a", x"7b", x"7b", x"7b", x"7a", x"79", x"79", x"78", x"77", x"78", x"79", x"78", x"77", x"78", 
        x"7a", x"7b", x"7b", x"7a", x"79", x"77", x"77", x"77", x"78", x"78", x"78", x"77", x"76", x"75", x"77", 
        x"76", x"75", x"74", x"74", x"75", x"77", x"78", x"74", x"73", x"73", x"73", x"73", x"73", x"73", x"74", 
        x"76", x"76", x"76", x"77", x"76", x"75", x"75", x"76", x"76", x"75", x"77", x"75", x"73", x"75", x"75", 
        x"75", x"75", x"75", x"75", x"75", x"75", x"76", x"76", x"77", x"77", x"76", x"76", x"75", x"76", x"76", 
        x"76", x"76", x"75", x"75", x"75", x"75", x"75", x"76", x"78", x"77", x"75", x"75", x"75", x"75", x"77", 
        x"77", x"76", x"75", x"76", x"75", x"73", x"76", x"76", x"75", x"77", x"76", x"74", x"77", x"78", x"77", 
        x"76", x"77", x"77", x"74", x"75", x"75", x"77", x"78", x"79", x"78", x"78", x"78", x"76", x"75", x"75", 
        x"76", x"77", x"77", x"75", x"76", x"78", x"77", x"77", x"78", x"78", x"76", x"77", x"79", x"7b", x"7a", 
        x"78", x"77", x"78", x"79", x"7a", x"79", x"79", x"79", x"7b", x"7d", x"7c", x"7c", x"7b", x"7a", x"78", 
        x"77", x"76", x"7a", x"78", x"79", x"7a", x"79", x"7b", x"79", x"78", x"79", x"7a", x"7a", x"7b", x"7c", 
        x"7c", x"7c", x"7b", x"7b", x"7c", x"7c", x"7c", x"7c", x"7d", x"7a", x"7a", x"7b", x"7c", x"7c", x"77", 
        x"7f", x"cc", x"d8", x"d2", x"d8", x"d2", x"b9", x"95", x"aa", x"c9", x"d5", x"ce", x"c8", x"ce", x"ce", 
        x"cb", x"cc", x"cd", x"cc", x"cc", x"cd", x"ce", x"cd", x"cb", x"cb", x"cc", x"ce", x"cf", x"ce", x"cf", 
        x"d0", x"ce", x"cd", x"cd", x"ce", x"cf", x"ce", x"cd", x"ce", x"ce", x"cd", x"cd", x"ce", x"d0", x"d0", 
        x"cf", x"cf", x"cf", x"cf", x"cf", x"cd", x"cc", x"d8", x"da", x"d0", x"d4", x"d3", x"d0", x"d2", x"ce", 
        x"b7", x"6f", x"5c", x"5c", x"5e", x"5b", x"5e", x"60", x"63", x"a7", x"e9", x"ee", x"df", x"c5", x"a4", 
        x"84", x"6f", x"63", x"5d", x"5d", x"5f", x"5e", x"5f", x"5d", x"5c", x"5e", x"5d", x"5d", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5a", x"5b", x"5f", 
        x"5d", x"5c", x"61", x"76", x"a1", x"d3", x"ee", x"f5", x"f8", x"fa", x"f9", x"fb", x"fa", x"fa", x"fb", 
        x"fa", x"f8", x"f7", x"f7", x"fa", x"fc", x"fc", x"fa", x"f9", x"f8", x"f8", x"f9", x"fb", x"fb", x"fb", 
        x"fa", x"f8", x"f6", x"f2", x"ec", x"e8", x"e5", x"eb", x"eb", x"e4", x"c4", x"90", x"6a", x"60", x"7a", 
        x"c7", x"db", x"bf", x"ae", x"ad", x"c7", x"e1", x"ec", x"eb", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", 
        x"f1", x"ef", x"ec", x"ec", x"f1", x"ee", x"ed", x"e9", x"dd", x"cf", x"ca", x"d9", x"e1", x"ce", x"a3", 
        x"7f", x"75", x"79", x"7e", x"85", x"87", x"83", x"82", x"83", x"81", x"80", x"80", x"80", x"80", x"80", 
        x"80", x"80", x"7f", x"7f", x"7f", x"80", x"80", x"7f", x"7f", x"80", x"80", x"80", x"80", x"80", x"80", 
        x"80", x"7f", x"7f", x"81", x"81", x"80", x"7f", x"80", x"81", x"82", x"80", x"80", x"80", x"81", x"81", 
        x"7f", x"7e", x"7f", x"80", x"80", x"7f", x"7e", x"7f", x"80", x"80", x"80", x"7e", x"7d", x"7e", x"7d", 
        x"80", x"82", x"7f", x"7f", x"80", x"80", x"7f", x"7e", x"7e", x"7d", x"7d", x"7d", x"7e", x"7f", x"7f", 
        x"7d", x"7f", x"80", x"80", x"80", x"80", x"80", x"80", x"7f", x"80", x"7e", x"7b", x"7d", x"7f", x"7e", 
        x"7f", x"7f", x"7e", x"7d", x"7d", x"7f", x"80", x"7f", x"7e", x"7e", x"7e", x"7e", x"7d", x"7f", x"80", 
        x"7f", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7f", 
        x"7d", x"7c", x"7d", x"7b", x"7d", x"7c", x"7c", x"7e", x"7e", x"7d", x"7d", x"7e", x"7f", x"7e", x"7d", 
        x"7d", x"7e", x"7e", x"7d", x"7d", x"7f", x"7e", x"7c", x"7b", x"7a", x"79", x"79", x"7a", x"7c", x"7e", 
        x"7e", x"7d", x"7b", x"7a", x"7a", x"7b", x"7b", x"7c", x"7d", x"7d", x"7d", x"7f", x"7e", x"7e", x"7c", 
        x"7c", x"7c", x"7b", x"7a", x"7c", x"7d", x"7a", x"79", x"78", x"78", x"7d", x"7d", x"7a", x"78", x"77", 
        x"7a", x"7c", x"7c", x"7b", x"7b", x"79", x"78", x"7b", x"7a", x"79", x"7b", x"7a", x"77", x"79", x"79", 
        x"79", x"79", x"7a", x"79", x"78", x"79", x"7a", x"7b", x"7a", x"7a", x"78", x"77", x"7a", x"7b", x"79", 
        x"79", x"79", x"7c", x"7b", x"7a", x"7c", x"7a", x"7a", x"7a", x"78", x"78", x"78", x"78", x"79", x"79", 
        x"79", x"79", x"7a", x"79", x"79", x"79", x"79", x"79", x"7b", x"7c", x"7d", x"7a", x"79", x"78", x"79", 
        x"79", x"7b", x"7c", x"7a", x"78", x"79", x"7c", x"7b", x"76", x"77", x"77", x"79", x"7a", x"79", x"78", 
        x"75", x"77", x"78", x"79", x"78", x"77", x"77", x"78", x"78", x"78", x"79", x"7a", x"7a", x"79", x"7b", 
        x"7b", x"79", x"79", x"79", x"79", x"7a", x"78", x"78", x"79", x"7a", x"7a", x"79", x"78", x"76", x"77", 
        x"78", x"76", x"75", x"73", x"74", x"78", x"77", x"75", x"75", x"75", x"74", x"74", x"73", x"73", x"75", 
        x"77", x"76", x"77", x"78", x"77", x"76", x"75", x"77", x"76", x"74", x"76", x"75", x"74", x"76", x"77", 
        x"78", x"78", x"78", x"78", x"78", x"76", x"76", x"77", x"77", x"77", x"76", x"75", x"77", x"78", x"78", 
        x"76", x"75", x"74", x"75", x"76", x"76", x"73", x"75", x"79", x"76", x"75", x"75", x"75", x"76", x"77", 
        x"78", x"77", x"76", x"75", x"75", x"77", x"77", x"77", x"77", x"79", x"79", x"76", x"77", x"78", x"77", 
        x"76", x"79", x"78", x"76", x"76", x"76", x"77", x"77", x"77", x"76", x"76", x"78", x"75", x"73", x"74", 
        x"74", x"77", x"78", x"79", x"7b", x"7a", x"79", x"78", x"78", x"78", x"77", x"78", x"79", x"7c", x"7b", 
        x"77", x"78", x"79", x"78", x"78", x"79", x"78", x"78", x"79", x"7a", x"7b", x"7a", x"7a", x"7a", x"79", 
        x"78", x"7a", x"7d", x"79", x"7a", x"7b", x"79", x"7a", x"7a", x"7a", x"7b", x"7b", x"7b", x"7a", x"7b", 
        x"7b", x"7e", x"7f", x"7d", x"7d", x"7c", x"7a", x"7a", x"7b", x"7b", x"7b", x"7a", x"7b", x"7b", x"76", 
        x"7e", x"c9", x"d4", x"d2", x"c5", x"9d", x"98", x"c5", x"cd", x"d1", x"c5", x"c9", x"cf", x"cd", x"c9", 
        x"cb", x"cd", x"cd", x"cd", x"cc", x"cd", x"ce", x"cb", x"cb", x"ce", x"ce", x"cd", x"cc", x"cd", x"ce", 
        x"cd", x"ce", x"cf", x"cf", x"cf", x"ce", x"cd", x"cd", x"cd", x"cd", x"cd", x"cd", x"cf", x"cf", x"cf", 
        x"cf", x"cf", x"cf", x"cf", x"ce", x"cd", x"cb", x"d6", x"d9", x"cf", x"d3", x"d1", x"cf", x"d2", x"cf", 
        x"ba", x"70", x"5b", x"5c", x"5f", x"60", x"61", x"5e", x"61", x"a8", x"ee", x"f9", x"f8", x"f8", x"f1", 
        x"df", x"c5", x"a1", x"7d", x"69", x"61", x"5a", x"60", x"61", x"5c", x"5c", x"5b", x"5d", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5e", 
        x"5e", x"5e", x"5d", x"5b", x"5d", x"77", x"a5", x"d2", x"e8", x"ef", x"f4", x"f5", x"f8", x"f9", x"fa", 
        x"fd", x"fb", x"fa", x"f9", x"f9", x"f9", x"fb", x"fc", x"fc", x"fc", x"fc", x"fb", x"f9", x"fa", x"fb", 
        x"fb", x"fa", x"fa", x"f7", x"f4", x"f6", x"f4", x"ec", x"dc", x"b9", x"7e", x"5a", x"5c", x"62", x"73", 
        x"c8", x"f3", x"f1", x"e6", x"ca", x"ad", x"a7", x"bc", x"d8", x"e7", x"ed", x"f1", x"ee", x"ea", x"ec", 
        x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"ef", 
        x"ed", x"ef", x"f0", x"f0", x"f0", x"ec", x"ed", x"f1", x"ed", x"eb", x"ec", x"d4", x"ce", x"d9", x"e5", 
        x"db", x"ae", x"86", x"74", x"74", x"79", x"7d", x"81", x"83", x"83", x"82", x"80", x"7f", x"80", x"80", 
        x"80", x"81", x"80", x"7e", x"7f", x"7f", x"80", x"7f", x"7e", x"7f", x"80", x"7f", x"80", x"7f", x"7f", 
        x"80", x"80", x"81", x"81", x"80", x"7f", x"7e", x"80", x"82", x"82", x"80", x"7e", x"80", x"82", x"81", 
        x"7e", x"7d", x"7f", x"81", x"82", x"81", x"7f", x"7f", x"81", x"82", x"82", x"80", x"7f", x"7f", x"7e", 
        x"80", x"80", x"7e", x"7e", x"7e", x"7f", x"7e", x"7e", x"7e", x"7f", x"80", x"80", x"7f", x"7f", x"7e", 
        x"7e", x"80", x"80", x"7e", x"7f", x"7f", x"7f", x"80", x"80", x"81", x"7f", x"7c", x"7f", x"7e", x"7f", 
        x"81", x"7f", x"7f", x"7f", x"80", x"80", x"80", x"80", x"7f", x"7f", x"7f", x"7f", x"7e", x"7f", x"80", 
        x"7e", x"7e", x"7f", x"7f", x"7e", x"7f", x"80", x"7f", x"7d", x"7d", x"7e", x"7d", x"7c", x"7f", x"81", 
        x"80", x"7f", x"7f", x"7c", x"7e", x"7d", x"7e", x"7f", x"7e", x"7f", x"7f", x"80", x"7f", x"80", x"7f", 
        x"7f", x"7e", x"7d", x"7e", x"7e", x"7f", x"7e", x"7d", x"7d", x"7b", x"7e", x"7d", x"7b", x"7c", x"7d", 
        x"7d", x"7d", x"7c", x"7b", x"7a", x"7a", x"7b", x"7c", x"7d", x"7e", x"7e", x"7f", x"7c", x"7d", x"7a", 
        x"7b", x"7b", x"7b", x"7b", x"7d", x"7d", x"7a", x"7a", x"79", x"79", x"7c", x"7c", x"7c", x"7b", x"7a", 
        x"7a", x"7c", x"7b", x"7a", x"7b", x"7a", x"79", x"7b", x"7a", x"78", x"7a", x"78", x"77", x"78", x"79", 
        x"7a", x"79", x"79", x"79", x"7a", x"7b", x"7b", x"7b", x"7a", x"7c", x"7b", x"79", x"79", x"79", x"79", 
        x"79", x"7a", x"7a", x"79", x"78", x"79", x"78", x"78", x"7a", x"7c", x"7a", x"7b", x"7c", x"7c", x"7b", 
        x"7b", x"7a", x"7c", x"7d", x"7a", x"7a", x"7b", x"79", x"79", x"7a", x"7b", x"7a", x"78", x"77", x"77", 
        x"78", x"79", x"7a", x"79", x"79", x"7a", x"7b", x"7b", x"78", x"78", x"78", x"79", x"7b", x"78", x"78", 
        x"78", x"7a", x"7a", x"7c", x"7b", x"7b", x"7a", x"78", x"76", x"76", x"77", x"79", x"79", x"79", x"79", 
        x"79", x"79", x"79", x"78", x"78", x"78", x"78", x"7a", x"7a", x"7c", x"7b", x"7a", x"7a", x"77", x"78", 
        x"78", x"76", x"76", x"74", x"76", x"79", x"75", x"76", x"77", x"76", x"75", x"74", x"73", x"73", x"74", 
        x"75", x"72", x"73", x"74", x"75", x"76", x"76", x"78", x"76", x"73", x"74", x"74", x"74", x"76", x"75", 
        x"76", x"77", x"77", x"77", x"76", x"74", x"74", x"76", x"78", x"78", x"76", x"75", x"75", x"79", x"79", 
        x"76", x"75", x"74", x"75", x"76", x"78", x"76", x"77", x"78", x"75", x"76", x"75", x"76", x"78", x"77", 
        x"77", x"77", x"76", x"75", x"76", x"78", x"77", x"75", x"77", x"7a", x"79", x"77", x"79", x"7a", x"78", 
        x"77", x"79", x"79", x"76", x"77", x"77", x"76", x"76", x"76", x"76", x"77", x"79", x"76", x"76", x"77", 
        x"76", x"78", x"76", x"79", x"7a", x"78", x"78", x"77", x"76", x"77", x"78", x"7a", x"7b", x"7a", x"78", 
        x"78", x"7a", x"7b", x"78", x"7a", x"7b", x"7b", x"7a", x"7a", x"7b", x"7e", x"7b", x"7a", x"7a", x"78", 
        x"77", x"7a", x"7c", x"79", x"7b", x"7c", x"78", x"78", x"79", x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", 
        x"7b", x"7d", x"7d", x"7c", x"7d", x"7d", x"7a", x"7b", x"7c", x"7d", x"7d", x"7c", x"7c", x"7c", x"77", 
        x"81", x"cf", x"cf", x"b0", x"9f", x"b3", x"d8", x"db", x"ca", x"cf", x"cc", x"cd", x"cb", x"cc", x"cd", 
        x"cc", x"cc", x"ce", x"ce", x"ce", x"cd", x"cd", x"cc", x"cd", x"ce", x"cf", x"ce", x"cd", x"cd", x"cd", 
        x"cc", x"ce", x"cf", x"cf", x"cf", x"cf", x"cf", x"cd", x"cd", x"cd", x"cd", x"cf", x"d0", x"d0", x"cf", 
        x"cf", x"cf", x"cf", x"cf", x"ce", x"cd", x"cb", x"d6", x"d9", x"cf", x"d3", x"d1", x"cf", x"d1", x"d0", 
        x"bc", x"72", x"5c", x"5d", x"5e", x"5e", x"5d", x"5f", x"61", x"a3", x"ec", x"f9", x"f9", x"f8", x"f8", 
        x"f7", x"f4", x"ea", x"d8", x"c3", x"9b", x"6d", x"61", x"63", x"60", x"5e", x"60", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"60", 
        x"5f", x"5a", x"5d", x"61", x"5f", x"5c", x"62", x"79", x"9a", x"af", x"bb", x"cd", x"e1", x"e7", x"e6", 
        x"f0", x"f8", x"fa", x"fb", x"fa", x"fa", x"fb", x"fc", x"fb", x"fa", x"fb", x"fb", x"fa", x"fa", x"fb", 
        x"fc", x"fc", x"f7", x"f3", x"ea", x"e0", x"c8", x"a6", x"89", x"6f", x"62", x"5e", x"60", x"5e", x"72", 
        x"ca", x"f0", x"ee", x"ed", x"ec", x"e9", x"db", x"c3", x"b0", x"b5", x"c1", x"d4", x"e3", x"ec", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"ef", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", 
        x"ef", x"f0", x"ef", x"ed", x"ee", x"eb", x"f0", x"f1", x"ef", x"f0", x"f0", x"ee", x"e8", x"d9", x"d2", 
        x"d6", x"dc", x"d5", x"ba", x"9b", x"7f", x"75", x"7a", x"81", x"83", x"83", x"82", x"80", x"81", x"81", 
        x"80", x"81", x"80", x"7d", x"7f", x"80", x"81", x"82", x"82", x"82", x"81", x"7f", x"80", x"7f", x"7f", 
        x"82", x"80", x"80", x"81", x"81", x"81", x"7f", x"7f", x"80", x"7f", x"7f", x"80", x"81", x"80", x"7f", 
        x"7e", x"7d", x"7f", x"82", x"83", x"81", x"80", x"7f", x"81", x"80", x"81", x"80", x"7f", x"80", x"7f", 
        x"80", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7e", x"7f", x"80", x"80", x"80", x"7f", x"7f", x"7e", 
        x"7f", x"80", x"7e", x"7d", x"7e", x"7f", x"7e", x"7e", x"7f", x"81", x"80", x"7f", x"81", x"7d", x"7d", 
        x"7f", x"7d", x"7d", x"7f", x"7f", x"7e", x"7e", x"80", x"7f", x"7e", x"7f", x"7f", x"7e", x"7e", x"7f", 
        x"7d", x"7f", x"81", x"80", x"7f", x"7f", x"7f", x"7e", x"7e", x"7f", x"80", x"7e", x"7c", x"7d", x"7f", 
        x"7d", x"7c", x"7d", x"7b", x"7e", x"7e", x"7e", x"7f", x"7d", x"7d", x"7e", x"7f", x"7f", x"80", x"80", 
        x"80", x"7d", x"7b", x"7e", x"7d", x"7d", x"7e", x"7e", x"7e", x"7b", x"7c", x"7a", x"7b", x"7b", x"7c", 
        x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7d", x"7b", x"7b", x"79", 
        x"79", x"7a", x"7b", x"7d", x"7e", x"7c", x"7a", x"7b", x"79", x"79", x"7b", x"7b", x"7c", x"7b", x"79", 
        x"79", x"7b", x"7b", x"79", x"7c", x"7b", x"7a", x"7b", x"79", x"78", x"79", x"79", x"7a", x"7b", x"7b", 
        x"7a", x"78", x"7a", x"7b", x"7c", x"7c", x"7b", x"7a", x"7a", x"79", x"7a", x"7a", x"79", x"79", x"7b", 
        x"7c", x"7b", x"7b", x"7a", x"7a", x"78", x"79", x"7a", x"7b", x"7d", x"7a", x"7b", x"7d", x"7c", x"7a", 
        x"7b", x"7b", x"7d", x"7b", x"77", x"78", x"7b", x"7b", x"7c", x"79", x"77", x"79", x"7c", x"7b", x"79", 
        x"78", x"79", x"79", x"79", x"78", x"78", x"78", x"79", x"77", x"78", x"78", x"7a", x"7c", x"7a", x"79", 
        x"77", x"77", x"77", x"78", x"79", x"7a", x"7a", x"79", x"78", x"77", x"78", x"79", x"79", x"79", x"79", 
        x"7a", x"7b", x"7b", x"7a", x"79", x"78", x"79", x"7b", x"7a", x"7c", x"7b", x"7b", x"7a", x"78", x"79", 
        x"78", x"77", x"77", x"76", x"76", x"77", x"73", x"75", x"76", x"75", x"73", x"72", x"72", x"72", x"74", 
        x"74", x"71", x"72", x"74", x"76", x"76", x"76", x"78", x"76", x"74", x"75", x"75", x"76", x"76", x"73", 
        x"75", x"74", x"73", x"74", x"74", x"73", x"73", x"76", x"78", x"77", x"76", x"75", x"76", x"79", x"78", 
        x"76", x"76", x"75", x"76", x"77", x"79", x"77", x"78", x"77", x"74", x"76", x"76", x"76", x"77", x"75", 
        x"74", x"76", x"78", x"78", x"77", x"76", x"75", x"75", x"76", x"79", x"77", x"76", x"7a", x"7a", x"78", 
        x"78", x"79", x"77", x"75", x"78", x"79", x"78", x"77", x"78", x"78", x"78", x"7c", x"79", x"77", x"77", 
        x"76", x"78", x"76", x"78", x"78", x"76", x"77", x"77", x"77", x"79", x"79", x"79", x"7c", x"7b", x"79", 
        x"7a", x"7a", x"79", x"76", x"78", x"7a", x"7a", x"7a", x"78", x"79", x"7a", x"79", x"79", x"7a", x"79", 
        x"79", x"7b", x"7c", x"7c", x"7c", x"7b", x"79", x"7a", x"7b", x"7a", x"79", x"7a", x"7b", x"7c", x"7d", 
        x"7c", x"7b", x"79", x"7a", x"7c", x"7d", x"7c", x"7c", x"7d", x"7e", x"7c", x"7b", x"7d", x"7c", x"78", 
        x"81", x"bf", x"aa", x"a3", x"ca", x"da", x"d6", x"d2", x"cb", x"d0", x"cc", x"cb", x"ce", x"d1", x"cd", 
        x"cb", x"cd", x"cf", x"cf", x"ce", x"cd", x"cc", x"cd", x"ce", x"ce", x"ce", x"d0", x"d0", x"ce", x"cd", 
        x"cd", x"ce", x"ce", x"cd", x"ce", x"d0", x"d0", x"ce", x"cd", x"cd", x"cf", x"d1", x"d2", x"d1", x"cf", 
        x"ce", x"ce", x"ce", x"cd", x"cd", x"cd", x"cb", x"d7", x"da", x"cf", x"d3", x"d3", x"d1", x"d1", x"d0", 
        x"bc", x"72", x"5d", x"5d", x"5e", x"5d", x"5d", x"61", x"60", x"a1", x"ee", x"fb", x"f8", x"ef", x"e3", 
        x"eb", x"f5", x"fa", x"fa", x"f7", x"e0", x"8d", x"63", x"5f", x"5e", x"5f", x"60", x"5c", x"5c", x"5c", 
        x"5e", x"5f", x"5d", x"5d", x"5e", x"5c", x"5d", x"5f", x"5e", x"5e", x"5d", x"5e", x"5e", x"5d", x"5d", 
        x"5d", x"5d", x"5c", x"5c", x"5d", x"5f", x"5e", x"5a", x"59", x"5e", x"66", x"77", x"91", x"9b", x"a0", 
        x"b4", x"c8", x"d4", x"e1", x"e9", x"f1", x"f7", x"f9", x"fb", x"fb", x"fb", x"f9", x"f8", x"f4", x"ed", 
        x"e3", x"dc", x"d0", x"c1", x"a7", x"89", x"6e", x"5b", x"5a", x"5b", x"5e", x"5c", x"60", x"5f", x"70", 
        x"c7", x"f0", x"ee", x"ed", x"ee", x"f0", x"f3", x"f3", x"ec", x"d1", x"b7", x"a5", x"b0", x"c8", x"dd", 
        x"e7", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"f1", 
        x"f2", x"f2", x"ef", x"ee", x"ef", x"e7", x"ed", x"f0", x"ef", x"f2", x"f2", x"f0", x"f2", x"f3", x"ea", 
        x"dd", x"d3", x"d5", x"e2", x"e3", x"cc", x"a0", x"7f", x"79", x"7b", x"7e", x"84", x"84", x"82", x"82", 
        x"80", x"80", x"81", x"80", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"80", x"82", x"80", x"7e", 
        x"81", x"81", x"80", x"81", x"83", x"81", x"81", x"7f", x"7e", x"7c", x"7f", x"81", x"81", x"80", x"7e", 
        x"7f", x"7e", x"7f", x"81", x"83", x"82", x"81", x"80", x"81", x"81", x"81", x"7f", x"7f", x"80", x"7f", 
        x"80", x"80", x"80", x"7f", x"7e", x"7e", x"7e", x"7f", x"81", x"80", x"7f", x"7f", x"7f", x"7f", x"80", 
        x"80", x"80", x"7f", x"7d", x"7e", x"7f", x"7e", x"7d", x"7e", x"80", x"81", x"81", x"82", x"7e", x"7f", 
        x"80", x"7d", x"7f", x"81", x"81", x"7e", x"7e", x"7f", x"7f", x"7e", x"7f", x"7f", x"7e", x"7f", x"7f", 
        x"7d", x"80", x"81", x"80", x"80", x"80", x"7e", x"7e", x"7e", x"7f", x"80", x"80", x"7e", x"7d", x"7f", 
        x"7e", x"7e", x"7f", x"7e", x"80", x"7f", x"7e", x"7e", x"7e", x"7d", x"7d", x"7f", x"7f", x"80", x"80", 
        x"7f", x"7d", x"7c", x"7e", x"7c", x"7b", x"7d", x"7f", x"7f", x"7a", x"79", x"78", x"7c", x"7c", x"7c", 
        x"7d", x"7c", x"7c", x"7c", x"7c", x"7d", x"7c", x"7b", x"7a", x"7b", x"7b", x"7e", x"7e", x"7d", x"7b", 
        x"7b", x"7c", x"7b", x"7d", x"7e", x"7c", x"79", x"7a", x"79", x"79", x"7a", x"7b", x"7d", x"7b", x"79", 
        x"79", x"7c", x"7c", x"7a", x"7c", x"7c", x"7b", x"7b", x"7b", x"78", x"79", x"7b", x"7c", x"7d", x"7b", 
        x"79", x"78", x"79", x"7c", x"7d", x"7c", x"7b", x"7b", x"7a", x"77", x"78", x"7a", x"7a", x"7a", x"7b", 
        x"7b", x"7c", x"7c", x"7a", x"7b", x"79", x"7a", x"7b", x"7a", x"7a", x"78", x"7a", x"7c", x"7b", x"7a", 
        x"7b", x"7c", x"7b", x"79", x"77", x"78", x"79", x"7a", x"7c", x"79", x"74", x"76", x"7a", x"7b", x"79", 
        x"7b", x"7b", x"7a", x"79", x"78", x"79", x"7a", x"7b", x"7a", x"7a", x"7a", x"79", x"7a", x"79", x"79", 
        x"77", x"77", x"79", x"79", x"7a", x"7c", x"7c", x"7b", x"7a", x"79", x"79", x"79", x"79", x"7a", x"7c", 
        x"7c", x"7b", x"7a", x"79", x"7a", x"7a", x"78", x"79", x"79", x"7b", x"7a", x"7a", x"7b", x"79", x"7a", 
        x"78", x"78", x"77", x"76", x"74", x"73", x"72", x"77", x"78", x"76", x"75", x"74", x"74", x"75", x"78", 
        x"74", x"74", x"77", x"77", x"78", x"76", x"74", x"74", x"74", x"74", x"76", x"76", x"75", x"75", x"75", 
        x"77", x"75", x"73", x"75", x"76", x"76", x"75", x"75", x"76", x"75", x"74", x"75", x"76", x"77", x"74", 
        x"75", x"78", x"79", x"77", x"77", x"78", x"76", x"75", x"76", x"75", x"74", x"76", x"77", x"78", x"76", 
        x"73", x"76", x"78", x"77", x"77", x"74", x"75", x"78", x"7a", x"7a", x"76", x"75", x"77", x"78", x"79", 
        x"79", x"78", x"77", x"77", x"78", x"79", x"78", x"77", x"78", x"78", x"76", x"79", x"79", x"78", x"79", 
        x"7a", x"79", x"77", x"78", x"79", x"78", x"78", x"78", x"7a", x"7a", x"7b", x"7a", x"7a", x"7a", x"7b", 
        x"7a", x"7a", x"78", x"78", x"7a", x"7b", x"7b", x"7a", x"79", x"77", x"7a", x"7b", x"7b", x"7c", x"7b", 
        x"7a", x"7a", x"7b", x"7f", x"7d", x"78", x"7b", x"7f", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", 
        x"7a", x"7b", x"7c", x"7e", x"7d", x"7d", x"7e", x"7c", x"7d", x"7d", x"7a", x"79", x"7e", x"7b", x"78", 
        x"78", x"a8", x"c6", x"d6", x"cd", x"d0", x"d8", x"d6", x"ca", x"cd", x"cf", x"cc", x"cc", x"cc", x"cc", 
        x"ce", x"ce", x"ce", x"ce", x"ce", x"cd", x"cc", x"cd", x"ce", x"ce", x"cf", x"d0", x"d0", x"d0", x"ce", 
        x"ce", x"ce", x"cd", x"cc", x"ce", x"cf", x"cd", x"cd", x"ce", x"cf", x"d0", x"d0", x"d0", x"d0", x"ce", 
        x"ce", x"ce", x"cd", x"cc", x"cc", x"cc", x"cb", x"d5", x"da", x"ce", x"d2", x"d2", x"d2", x"d1", x"cf", 
        x"ba", x"71", x"5c", x"5d", x"5f", x"5d", x"5d", x"61", x"61", x"a4", x"ef", x"fa", x"f6", x"d0", x"8f", 
        x"99", x"ba", x"d6", x"ec", x"f7", x"e6", x"8f", x"5a", x"5b", x"5d", x"61", x"75", x"83", x"6e", x"5f", 
        x"5a", x"5e", x"60", x"5d", x"5f", x"5e", x"60", x"60", x"5b", x"5d", x"5f", x"5f", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5d", x"5d", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5f", x"60", x"60", x"5f", 
        x"63", x"6d", x"77", x"82", x"91", x"a4", x"b2", x"ba", x"c0", x"c3", x"c1", x"ba", x"b1", x"a5", x"98", 
        x"89", x"7c", x"71", x"68", x"5f", x"5b", x"5d", x"60", x"5f", x"5d", x"5c", x"5e", x"5f", x"5e", x"71", 
        x"c5", x"f2", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f1", x"f0", x"e4", x"cc", x"b9", x"b2", 
        x"b6", x"c5", x"da", x"ed", x"f2", x"f1", x"ee", x"ed", x"f0", x"ee", x"ed", x"ee", x"ef", x"ee", x"ed", 
        x"f0", x"f0", x"ee", x"ee", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", 
        x"f2", x"f1", x"f0", x"ee", x"f0", x"ec", x"ec", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"f3", x"ef", x"e6", x"dd", x"d3", x"d6", x"de", x"d5", x"b5", x"94", x"77", x"72", x"76", x"7d", x"83", 
        x"83", x"83", x"85", x"82", x"81", x"81", x"80", x"80", x"81", x"82", x"80", x"80", x"84", x"86", x"84", 
        x"82", x"83", x"82", x"81", x"82", x"80", x"82", x"7f", x"7f", x"80", x"80", x"80", x"81", x"81", x"82", 
        x"82", x"7e", x"7e", x"80", x"82", x"82", x"82", x"80", x"81", x"82", x"81", x"80", x"7f", x"7e", x"7d", 
        x"7e", x"81", x"82", x"81", x"7e", x"7e", x"80", x"81", x"80", x"80", x"80", x"80", x"80", x"80", x"80", 
        x"80", x"80", x"80", x"7f", x"7f", x"7f", x"80", x"80", x"80", x"7f", x"7f", x"7f", x"80", x"81", x"83", 
        x"81", x"7f", x"80", x"80", x"7f", x"80", x"80", x"80", x"80", x"80", x"7e", x"7d", x"7e", x"7f", x"7c", 
        x"7c", x"80", x"7f", x"7f", x"82", x"81", x"7f", x"81", x"7e", x"7c", x"7e", x"81", x"7f", x"7e", x"7f", 
        x"80", x"80", x"7f", x"7f", x"80", x"7f", x"7d", x"7d", x"80", x"7f", x"7d", x"7d", x"7f", x"80", x"7f", 
        x"7f", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7f", x"7f", x"7e", x"7d", x"7d", x"7e", x"7e", x"7d", 
        x"7d", x"7c", x"7b", x"7b", x"7b", x"7d", x"7d", x"7c", x"7a", x"7a", x"7c", x"7e", x"7d", x"7d", x"7c", 
        x"7e", x"7e", x"7b", x"7c", x"7d", x"7c", x"7a", x"7a", x"7a", x"7b", x"79", x"7a", x"7d", x"7c", x"7a", 
        x"7b", x"7c", x"7b", x"7b", x"79", x"7b", x"7a", x"7b", x"7d", x"79", x"7b", x"7c", x"7c", x"7b", x"7a", 
        x"79", x"79", x"77", x"79", x"7b", x"7b", x"7b", x"7a", x"77", x"79", x"7a", x"7b", x"7b", x"7a", x"79", 
        x"78", x"7a", x"7b", x"79", x"78", x"79", x"7b", x"7a", x"7a", x"7a", x"79", x"7b", x"7b", x"7a", x"7b", 
        x"7b", x"7c", x"7a", x"7a", x"7e", x"7e", x"7b", x"7a", x"7a", x"7b", x"79", x"76", x"77", x"7b", x"7d", 
        x"79", x"7a", x"7b", x"7a", x"78", x"78", x"79", x"79", x"7a", x"79", x"7b", x"78", x"7b", x"7a", x"7b", 
        x"77", x"77", x"7a", x"79", x"79", x"7c", x"7a", x"7a", x"7a", x"7a", x"78", x"78", x"79", x"7a", x"7a", 
        x"7b", x"7a", x"79", x"78", x"78", x"78", x"77", x"78", x"7a", x"7c", x"79", x"78", x"7b", x"7b", x"79", 
        x"79", x"78", x"77", x"76", x"76", x"75", x"74", x"77", x"77", x"77", x"76", x"76", x"75", x"75", x"77", 
        x"75", x"75", x"76", x"76", x"78", x"75", x"73", x"74", x"74", x"74", x"75", x"75", x"75", x"75", x"74", 
        x"76", x"76", x"76", x"76", x"76", x"75", x"75", x"77", x"77", x"77", x"76", x"75", x"76", x"76", x"74", 
        x"76", x"77", x"77", x"75", x"76", x"77", x"77", x"76", x"76", x"75", x"76", x"76", x"75", x"77", x"78", 
        x"75", x"77", x"78", x"77", x"77", x"76", x"76", x"77", x"79", x"79", x"77", x"76", x"78", x"79", x"7a", 
        x"78", x"77", x"77", x"78", x"79", x"78", x"78", x"79", x"78", x"77", x"77", x"76", x"76", x"77", x"79", 
        x"7a", x"7a", x"79", x"78", x"78", x"77", x"77", x"77", x"78", x"78", x"7a", x"7b", x"7a", x"7a", x"7a", 
        x"7a", x"7b", x"7a", x"7a", x"7b", x"7b", x"7b", x"7a", x"79", x"78", x"7b", x"7c", x"7c", x"7c", x"7b", 
        x"7b", x"7b", x"7b", x"7c", x"7b", x"79", x"7a", x"7c", x"7c", x"7c", x"7c", x"7a", x"7b", x"7c", x"7c", 
        x"7c", x"7b", x"7b", x"7d", x"7e", x"7d", x"7e", x"7b", x"7c", x"7d", x"7e", x"7b", x"7e", x"7c", x"78", 
        x"79", x"c1", x"d8", x"d2", x"c9", x"cf", x"d7", x"da", x"cb", x"cd", x"cf", x"cc", x"cc", x"cd", x"cc", 
        x"cd", x"ce", x"ce", x"ce", x"ce", x"cd", x"cd", x"cd", x"ce", x"ce", x"cf", x"cf", x"cf", x"d0", x"cf", 
        x"ce", x"ce", x"cb", x"ca", x"cc", x"cd", x"cd", x"cf", x"d0", x"d0", x"d0", x"d0", x"cf", x"cf", x"d0", 
        x"cf", x"cf", x"cf", x"ce", x"ce", x"cd", x"ca", x"d5", x"db", x"d0", x"d3", x"d2", x"d1", x"d0", x"cf", 
        x"ba", x"71", x"5c", x"5d", x"5f", x"5d", x"5d", x"60", x"61", x"a3", x"f0", x"fa", x"f7", x"c9", x"6e", 
        x"5b", x"6d", x"83", x"a0", x"bf", x"cb", x"89", x"5b", x"5d", x"5d", x"63", x"95", x"ce", x"bb", x"9e", 
        x"84", x"67", x"5c", x"5f", x"60", x"5f", x"60", x"5d", x"5c", x"5e", x"5c", x"5e", x"5f", x"5d", x"5d", 
        x"5e", x"5e", x"5d", x"5c", x"5d", x"5d", x"5d", x"5e", x"5e", x"5f", x"5e", x"5d", x"5f", x"60", x"5e", 
        x"5c", x"5d", x"5e", x"5b", x"5e", x"63", x"69", x"6e", x"71", x"72", x"73", x"6f", x"67", x"60", x"5d", 
        x"5c", x"5b", x"5b", x"5b", x"5c", x"5d", x"5e", x"5e", x"5d", x"5c", x"5c", x"5e", x"5e", x"5d", x"6e", 
        x"c2", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f3", x"ee", x"d8", 
        x"c4", x"b9", x"b7", x"be", x"cf", x"e4", x"ee", x"ef", x"f0", x"f0", x"ee", x"ec", x"ed", x"ef", x"ee", 
        x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f2", x"f1", x"f0", x"ee", x"f0", x"ec", x"eb", x"f0", x"f0", x"f1", x"f1", x"f0", x"f2", x"f3", x"f0", 
        x"f1", x"f2", x"f3", x"f1", x"e5", x"dc", x"d9", x"db", x"df", x"d8", x"bb", x"99", x"7e", x"73", x"78", 
        x"7d", x"83", x"85", x"84", x"83", x"83", x"83", x"82", x"80", x"82", x"83", x"81", x"82", x"84", x"83", 
        x"83", x"84", x"82", x"81", x"83", x"82", x"82", x"80", x"7f", x"81", x"81", x"81", x"81", x"82", x"82", 
        x"81", x"80", x"80", x"80", x"81", x"81", x"81", x"81", x"81", x"82", x"81", x"81", x"80", x"80", x"80", 
        x"7f", x"7e", x"7f", x"7f", x"7f", x"7f", x"81", x"81", x"80", x"80", x"80", x"80", x"80", x"80", x"80", 
        x"81", x"81", x"80", x"81", x"81", x"80", x"7e", x"7f", x"80", x"80", x"80", x"80", x"80", x"81", x"81", 
        x"80", x"7f", x"81", x"80", x"7e", x"7f", x"80", x"80", x"81", x"80", x"7f", x"7d", x"7e", x"7e", x"7c", 
        x"7d", x"7f", x"7f", x"80", x"81", x"82", x"81", x"81", x"80", x"7e", x"7f", x"81", x"80", x"80", x"80", 
        x"81", x"7f", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7e", x"7e", x"7d", x"7d", x"7e", x"7f", x"80", 
        x"80", x"7d", x"7c", x"7e", x"7f", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7c", x"7c", x"7c", 
        x"7c", x"7c", x"7d", x"7d", x"7c", x"7d", x"7e", x"7e", x"7c", x"7b", x"7c", x"7d", x"7d", x"7d", x"7d", 
        x"7e", x"7d", x"7b", x"7a", x"7b", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7c", x"7d", x"7b", x"7a", 
        x"7b", x"7c", x"7a", x"79", x"79", x"7a", x"79", x"79", x"7b", x"79", x"7a", x"7a", x"7a", x"7b", x"7b", 
        x"7b", x"7b", x"79", x"79", x"79", x"7b", x"7a", x"79", x"78", x"79", x"7a", x"7b", x"7c", x"7b", x"7b", 
        x"7a", x"7a", x"79", x"79", x"7a", x"7b", x"7b", x"7a", x"79", x"79", x"79", x"7a", x"7b", x"7b", x"7c", 
        x"7c", x"7a", x"79", x"7b", x"7d", x"7d", x"7b", x"7c", x"7c", x"7b", x"7a", x"78", x"78", x"79", x"7b", 
        x"7a", x"7a", x"7a", x"79", x"78", x"79", x"7a", x"7b", x"7b", x"78", x"79", x"77", x"7b", x"7b", x"7e", 
        x"7a", x"7a", x"7c", x"7a", x"7a", x"7c", x"7a", x"7a", x"7b", x"7b", x"7a", x"79", x"7a", x"7b", x"7a", 
        x"7a", x"7a", x"79", x"79", x"79", x"79", x"7a", x"7b", x"7c", x"7d", x"7a", x"79", x"7c", x"7c", x"7b", 
        x"78", x"78", x"78", x"77", x"77", x"77", x"76", x"76", x"77", x"77", x"77", x"76", x"75", x"74", x"76", 
        x"76", x"76", x"76", x"75", x"78", x"74", x"73", x"76", x"76", x"76", x"76", x"77", x"77", x"77", x"76", 
        x"77", x"77", x"78", x"77", x"75", x"73", x"77", x"78", x"78", x"77", x"76", x"76", x"77", x"76", x"76", 
        x"77", x"76", x"74", x"73", x"74", x"76", x"78", x"78", x"75", x"76", x"78", x"77", x"74", x"77", x"79", 
        x"76", x"77", x"78", x"77", x"78", x"77", x"77", x"78", x"79", x"79", x"78", x"77", x"7a", x"79", x"79", 
        x"79", x"79", x"79", x"78", x"79", x"78", x"79", x"7a", x"78", x"76", x"79", x"77", x"77", x"78", x"79", 
        x"7a", x"79", x"77", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7a", x"7a", x"79", x"7a", x"7a", 
        x"7b", x"7c", x"7c", x"7b", x"7b", x"7a", x"7a", x"7b", x"7c", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", 
        x"7c", x"7c", x"7c", x"7b", x"7c", x"7e", x"7c", x"7b", x"7d", x"7d", x"7c", x"7b", x"7a", x"7b", x"7c", 
        x"7d", x"7c", x"7b", x"7d", x"7e", x"7e", x"7e", x"7b", x"7b", x"7b", x"7f", x"7c", x"7e", x"7e", x"79", 
        x"78", x"c3", x"d6", x"cd", x"d0", x"d2", x"d5", x"d9", x"cb", x"cd", x"ce", x"cc", x"cc", x"ce", x"cd", 
        x"cd", x"cd", x"cd", x"cd", x"ce", x"ce", x"ce", x"ce", x"ce", x"ce", x"cf", x"cf", x"cf", x"cf", x"cf", 
        x"cf", x"ce", x"cc", x"ca", x"cb", x"cd", x"cd", x"d0", x"d1", x"d2", x"d1", x"d0", x"cf", x"ce", x"d1", 
        x"d0", x"cf", x"cf", x"d0", x"cf", x"cd", x"ca", x"d6", x"dc", x"d1", x"d4", x"d1", x"cf", x"d0", x"cf", 
        x"ba", x"71", x"5c", x"5d", x"5f", x"5d", x"5d", x"60", x"61", x"a1", x"ef", x"fb", x"f8", x"d6", x"87", 
        x"5f", x"58", x"55", x"5c", x"6f", x"7b", x"6c", x"5c", x"62", x"5f", x"5f", x"99", x"eb", x"f6", x"ed", 
        x"d9", x"a0", x"69", x"60", x"60", x"5e", x"5e", x"5b", x"5e", x"61", x"5a", x"5e", x"5f", x"5c", x"5c", 
        x"5d", x"5f", x"5d", x"5c", x"5d", x"5d", x"5d", x"5e", x"5e", x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"60", x"5c", x"5a", x"5c", x"5e", x"5e", x"5b", x"5c", x"5d", x"5d", x"5d", x"5d", 
        x"5e", x"5f", x"5e", x"5e", x"5f", x"5d", x"5c", x"5c", x"5d", x"5d", x"5d", x"5e", x"5d", x"5c", x"6b", 
        x"bc", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"ee", x"ef", x"f3", 
        x"f4", x"ea", x"db", x"c7", x"b5", x"ab", x"bb", x"d8", x"f0", x"f5", x"f2", x"ee", x"ee", x"f0", x"ef", 
        x"ec", x"ed", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f2", x"f1", x"f0", x"ee", x"f0", x"ec", x"eb", x"f0", x"f0", x"f1", x"f1", x"f0", x"f3", x"f4", x"f2", 
        x"f0", x"ef", x"ed", x"ef", x"f1", x"f0", x"ea", x"e1", x"dc", x"d8", x"dc", x"df", x"cf", x"ac", x"82", 
        x"6b", x"72", x"83", x"84", x"86", x"86", x"84", x"82", x"83", x"84", x"83", x"84", x"85", x"83", x"81", 
        x"83", x"84", x"7f", x"7f", x"81", x"81", x"81", x"80", x"80", x"83", x"82", x"82", x"82", x"82", x"82", 
        x"82", x"82", x"82", x"81", x"80", x"80", x"81", x"82", x"83", x"83", x"82", x"82", x"81", x"80", x"7f", 
        x"7f", x"80", x"7f", x"7f", x"7f", x"80", x"80", x"80", x"81", x"81", x"81", x"81", x"81", x"81", x"81", 
        x"82", x"81", x"81", x"82", x"83", x"81", x"7e", x"7d", x"7e", x"7f", x"81", x"81", x"81", x"81", x"80", 
        x"7f", x"80", x"81", x"80", x"7e", x"7f", x"7f", x"80", x"80", x"80", x"7f", x"7f", x"7e", x"7e", x"80", 
        x"81", x"80", x"80", x"7f", x"7d", x"80", x"81", x"81", x"80", x"7f", x"80", x"81", x"81", x"81", x"82", 
        x"82", x"80", x"7e", x"7d", x"7e", x"7e", x"7e", x"7e", x"7f", x"7e", x"7e", x"7e", x"7f", x"7f", x"7e", 
        x"7e", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", x"7f", x"7e", x"7e", x"7f", x"7e", x"7d", x"7c", x"7b", 
        x"7a", x"7b", x"7c", x"7d", x"7d", x"7d", x"7e", x"7e", x"7e", x"7c", x"7b", x"7d", x"7c", x"7c", x"7e", 
        x"7d", x"7b", x"7b", x"7c", x"7e", x"7e", x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", x"7c", x"7a", x"7c", 
        x"7e", x"7c", x"7a", x"7b", x"7b", x"7c", x"7b", x"7a", x"7c", x"7c", x"7b", x"79", x"79", x"7b", x"7d", 
        x"7d", x"7d", x"7a", x"78", x"78", x"79", x"78", x"77", x"79", x"7a", x"7b", x"7c", x"7c", x"7d", x"7c", 
        x"7c", x"7a", x"7a", x"7a", x"7a", x"7b", x"7b", x"7b", x"79", x"79", x"7b", x"79", x"7b", x"7d", x"7c", 
        x"7c", x"7a", x"7a", x"7b", x"7b", x"7a", x"79", x"7b", x"7c", x"7b", x"7b", x"7b", x"79", x"78", x"7a", 
        x"7a", x"79", x"77", x"78", x"79", x"7b", x"7c", x"7d", x"7d", x"78", x"79", x"77", x"7c", x"7c", x"7e", 
        x"7c", x"7b", x"7d", x"7a", x"7a", x"7c", x"79", x"78", x"7a", x"7b", x"7a", x"78", x"78", x"79", x"7a", 
        x"79", x"79", x"79", x"7a", x"79", x"79", x"79", x"7a", x"7c", x"7d", x"7b", x"7b", x"7d", x"7e", x"7c", 
        x"77", x"77", x"77", x"77", x"77", x"77", x"77", x"77", x"76", x"76", x"76", x"76", x"75", x"76", x"77", 
        x"77", x"78", x"77", x"75", x"77", x"75", x"74", x"76", x"76", x"76", x"77", x"77", x"77", x"78", x"77", 
        x"76", x"76", x"78", x"78", x"76", x"76", x"77", x"78", x"77", x"76", x"75", x"77", x"78", x"74", x"75", 
        x"76", x"75", x"75", x"76", x"77", x"76", x"78", x"79", x"77", x"77", x"79", x"78", x"75", x"78", x"79", 
        x"76", x"77", x"77", x"78", x"79", x"77", x"77", x"79", x"7a", x"7a", x"77", x"77", x"7b", x"79", x"78", 
        x"79", x"7a", x"79", x"78", x"77", x"7a", x"7a", x"78", x"78", x"79", x"7a", x"7a", x"7b", x"7b", x"7a", 
        x"79", x"78", x"77", x"7a", x"7b", x"7b", x"7a", x"7a", x"79", x"79", x"79", x"7a", x"79", x"7a", x"7a", 
        x"7c", x"7c", x"7c", x"7b", x"7a", x"7a", x"7a", x"7b", x"7c", x"7d", x"7c", x"7b", x"7a", x"7a", x"7b", 
        x"7b", x"7c", x"7c", x"7b", x"7c", x"80", x"7e", x"7b", x"7c", x"7c", x"7c", x"7d", x"7d", x"7c", x"7c", 
        x"7c", x"7c", x"7b", x"7d", x"7e", x"7e", x"7e", x"7b", x"7c", x"7c", x"7e", x"7e", x"7f", x"7d", x"7a", 
        x"78", x"c1", x"d8", x"d1", x"d1", x"d4", x"db", x"d7", x"cb", x"cc", x"cd", x"cc", x"cd", x"cf", x"ce", 
        x"cd", x"cc", x"cc", x"cd", x"ce", x"cf", x"d0", x"cf", x"ce", x"ce", x"cf", x"cf", x"cf", x"cf", x"cf", 
        x"d0", x"cf", x"ce", x"ce", x"cd", x"cd", x"ce", x"cf", x"cf", x"d0", x"d0", x"d0", x"cf", x"cf", x"d0", 
        x"cf", x"cd", x"ce", x"ce", x"cd", x"cc", x"cb", x"d6", x"dc", x"d1", x"d3", x"d2", x"d0", x"d1", x"cf", 
        x"ba", x"71", x"5c", x"5d", x"5f", x"5e", x"5e", x"5f", x"61", x"9e", x"ee", x"fc", x"f9", x"f0", x"dc", 
        x"c1", x"a5", x"85", x"6c", x"62", x"5d", x"5f", x"5c", x"5c", x"5e", x"5e", x"94", x"ec", x"f9", x"f8", 
        x"f7", x"de", x"91", x"5e", x"5a", x"5c", x"60", x"69", x"60", x"5d", x"60", x"60", x"5e", x"5c", x"5c", 
        x"5d", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5c", x"5d", x"5e", x"60", 
        x"5f", x"5e", x"5d", x"5e", x"5e", x"5e", x"5f", x"60", x"60", x"5f", x"5e", x"5f", x"60", x"5f", x"5d", 
        x"5d", x"5f", x"5f", x"5f", x"5f", x"5e", x"5f", x"5e", x"5e", x"5e", x"5e", x"5d", x"5c", x"5c", x"69", 
        x"b6", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"ed", x"ed", x"ed", x"ed", x"ee", 
        x"ef", x"ee", x"f2", x"f0", x"e6", x"d8", x"c7", x"b8", x"b4", x"c6", x"dd", x"ed", x"f1", x"ee", x"ed", 
        x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f2", x"f1", x"f0", x"ee", x"f0", x"ec", x"eb", x"f0", x"f0", x"f1", x"f1", x"f1", x"ef", x"ed", x"f0", 
        x"f1", x"f0", x"ee", x"ee", x"f2", x"f1", x"ee", x"ef", x"ee", x"e7", x"e1", x"d8", x"d7", x"dd", x"d4", 
        x"b7", x"91", x"78", x"79", x"7d", x"80", x"82", x"84", x"82", x"81", x"84", x"85", x"85", x"83", x"82", 
        x"82", x"82", x"7f", x"80", x"82", x"81", x"80", x"81", x"81", x"82", x"81", x"81", x"81", x"82", x"83", 
        x"84", x"83", x"82", x"82", x"82", x"82", x"81", x"82", x"82", x"82", x"82", x"81", x"80", x"7f", x"7f", 
        x"7f", x"82", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", 
        x"81", x"82", x"83", x"82", x"81", x"7f", x"7e", x"7e", x"7f", x"81", x"81", x"81", x"81", x"80", x"7e", 
        x"7e", x"81", x"81", x"80", x"7f", x"7f", x"80", x"80", x"81", x"81", x"81", x"80", x"7f", x"7e", x"7f", 
        x"81", x"80", x"80", x"80", x"7d", x"80", x"80", x"7f", x"80", x"80", x"7f", x"7f", x"80", x"80", x"81", 
        x"82", x"82", x"80", x"7f", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"80", x"7f", x"7e", 
        x"7d", x"7e", x"7f", x"7e", x"7e", x"80", x"80", x"7f", x"7e", x"7e", x"7f", x"7e", x"7e", x"7d", x"7b", 
        x"7b", x"7c", x"7d", x"7e", x"7f", x"7e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7e", 
        x"7d", x"7a", x"7b", x"7e", x"7f", x"7e", x"7d", x"7d", x"7d", x"7d", x"7b", x"7b", x"7d", x"7c", x"7d", 
        x"7f", x"7e", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7a", x"7c", x"7c", x"7b", x"7a", x"7b", x"7c", 
        x"7c", x"7c", x"7b", x"79", x"79", x"7a", x"79", x"78", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", 
        x"7a", x"7b", x"7c", x"7b", x"7b", x"7a", x"7a", x"7c", x"7b", x"7b", x"7d", x"7a", x"7b", x"7d", x"7c", 
        x"7b", x"7b", x"7b", x"7c", x"7b", x"79", x"78", x"7b", x"7b", x"7a", x"7a", x"7c", x"7b", x"79", x"7a", 
        x"7b", x"7a", x"78", x"78", x"79", x"7b", x"7c", x"7d", x"7d", x"79", x"7b", x"79", x"7d", x"7b", x"7c", 
        x"7a", x"7a", x"7c", x"7a", x"7a", x"7c", x"79", x"78", x"79", x"7b", x"7a", x"79", x"78", x"79", x"7a", 
        x"79", x"79", x"7a", x"7b", x"7a", x"79", x"78", x"7a", x"7c", x"7d", x"7c", x"7b", x"7b", x"7b", x"7b", 
        x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"78", 
        x"76", x"78", x"78", x"76", x"77", x"76", x"74", x"75", x"75", x"75", x"76", x"76", x"76", x"76", x"76", 
        x"75", x"76", x"78", x"78", x"79", x"79", x"76", x"78", x"79", x"79", x"78", x"78", x"78", x"75", x"75", 
        x"76", x"75", x"76", x"78", x"79", x"77", x"78", x"79", x"79", x"79", x"79", x"78", x"76", x"78", x"79", 
        x"76", x"77", x"78", x"78", x"79", x"78", x"78", x"7a", x"7b", x"7a", x"77", x"76", x"7a", x"7b", x"7a", 
        x"78", x"76", x"78", x"79", x"78", x"7b", x"7a", x"78", x"79", x"7b", x"7a", x"7a", x"7b", x"7b", x"7a", 
        x"79", x"79", x"7a", x"79", x"79", x"79", x"79", x"79", x"79", x"78", x"78", x"79", x"7a", x"7b", x"7b", 
        x"7b", x"7a", x"7b", x"7c", x"7c", x"7a", x"7a", x"7a", x"7b", x"7b", x"7a", x"7a", x"79", x"79", x"79", 
        x"7a", x"7a", x"7b", x"7a", x"7b", x"7e", x"7c", x"79", x"7b", x"7a", x"7a", x"7c", x"7e", x"7e", x"7e", 
        x"7e", x"7f", x"7e", x"7f", x"7f", x"7f", x"7f", x"7e", x"80", x"7f", x"7d", x"7f", x"7f", x"7c", x"79", 
        x"7a", x"c3", x"da", x"d4", x"d0", x"d1", x"db", x"d7", x"cb", x"cc", x"cd", x"cc", x"ce", x"d0", x"cf", 
        x"cd", x"cc", x"cc", x"cc", x"cd", x"cf", x"d1", x"d0", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", 
        x"d0", x"cf", x"d1", x"d0", x"ce", x"ce", x"ce", x"ce", x"ce", x"ce", x"ce", x"cf", x"d0", x"d0", x"cf", 
        x"ce", x"cd", x"cd", x"cd", x"cc", x"cb", x"cc", x"d7", x"dc", x"d0", x"d3", x"d2", x"d2", x"d1", x"cf", 
        x"ba", x"71", x"5c", x"5d", x"5f", x"5e", x"5d", x"5f", x"61", x"9d", x"ee", x"fd", x"fa", x"f9", x"fb", 
        x"f2", x"e9", x"dc", x"c3", x"a7", x"7f", x"5f", x"5d", x"5d", x"60", x"5f", x"90", x"eb", x"fb", x"f9", 
        x"f8", x"f3", x"bb", x"6b", x"5b", x"5b", x"6d", x"aa", x"a0", x"82", x"68", x"5d", x"5c", x"5d", x"5e", 
        x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5e", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5f", x"5f", 
        x"5e", x"5d", x"5c", x"5d", x"5e", x"5f", x"5e", x"5d", x"5e", x"5f", x"5d", x"5e", x"5f", x"5e", x"5e", 
        x"5f", x"61", x"60", x"5e", x"5d", x"5d", x"5f", x"5f", x"5e", x"5d", x"5e", x"5d", x"5b", x"5d", x"68", 
        x"b3", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"ee", x"e4", x"d7", x"bf", x"b1", x"ba", x"d5", x"e8", x"f0", 
        x"f0", x"f0", x"ee", x"ef", x"f1", x"f2", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f2", x"f1", x"f0", x"ee", x"f0", x"ec", x"eb", x"f0", x"f0", x"f1", x"f2", x"f3", x"f0", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"f2", x"f3", x"ef", x"ee", x"f1", x"f2", x"f1", x"f0", x"e8", x"db", x"d1", x"d1", 
        x"dc", x"da", x"bd", x"98", x"7b", x"72", x"7b", x"82", x"84", x"85", x"85", x"85", x"80", x"7b", x"7b", 
        x"7d", x"80", x"83", x"86", x"85", x"83", x"80", x"82", x"83", x"82", x"80", x"80", x"80", x"82", x"83", 
        x"84", x"82", x"82", x"82", x"83", x"83", x"82", x"81", x"81", x"80", x"80", x"80", x"80", x"80", x"80", 
        x"80", x"81", x"81", x"81", x"81", x"82", x"83", x"83", x"81", x"81", x"81", x"81", x"81", x"81", x"80", 
        x"7f", x"81", x"82", x"82", x"7f", x"7e", x"7f", x"82", x"83", x"83", x"82", x"81", x"7f", x"7e", x"7d", 
        x"7f", x"80", x"80", x"7f", x"80", x"80", x"80", x"81", x"81", x"81", x"82", x"81", x"7f", x"7e", x"7e", 
        x"7f", x"80", x"80", x"80", x"80", x"82", x"80", x"7f", x"7f", x"80", x"80", x"7f", x"7f", x"7f", x"80", 
        x"81", x"81", x"80", x"7f", x"7f", x"7f", x"80", x"7f", x"7e", x"7e", x"80", x"80", x"7f", x"80", x"80", 
        x"7f", x"7e", x"7e", x"7f", x"80", x"80", x"80", x"80", x"7f", x"7f", x"7e", x"7d", x"7d", x"7c", x"7c", 
        x"7d", x"7e", x"7f", x"81", x"80", x"7e", x"7d", x"7c", x"7c", x"7d", x"7e", x"7e", x"7d", x"7d", x"7e", 
        x"7e", x"7c", x"7b", x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", x"80", x"7b", x"79", x"80", x"7f", x"7c", 
        x"7c", x"7e", x"7d", x"7c", x"7d", x"7c", x"7d", x"7c", x"7b", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", 
        x"7c", x"7a", x"7b", x"7b", x"7a", x"7b", x"7b", x"7a", x"7c", x"7c", x"7b", x"7b", x"7c", x"7b", x"7b", 
        x"7a", x"7c", x"7e", x"7c", x"7a", x"7a", x"7b", x"7c", x"7c", x"7c", x"7d", x"7b", x"7c", x"7c", x"7b", 
        x"7b", x"7a", x"7a", x"7b", x"7b", x"7a", x"7b", x"7d", x"7c", x"7a", x"7a", x"7c", x"7b", x"7a", x"7a", 
        x"7d", x"7d", x"7b", x"7a", x"79", x"79", x"79", x"7c", x"7d", x"7b", x"7c", x"7b", x"7d", x"7b", x"7b", 
        x"78", x"78", x"7b", x"79", x"7a", x"7c", x"7a", x"7a", x"7b", x"7c", x"7b", x"7a", x"7a", x"7b", x"7a", 
        x"7a", x"7a", x"7a", x"7b", x"7b", x"7a", x"79", x"7b", x"7d", x"7b", x"7a", x"79", x"77", x"78", x"79", 
        x"77", x"77", x"77", x"77", x"77", x"76", x"76", x"75", x"76", x"76", x"77", x"77", x"77", x"76", x"77", 
        x"76", x"77", x"79", x"77", x"77", x"78", x"76", x"75", x"75", x"75", x"76", x"76", x"76", x"77", x"77", 
        x"76", x"77", x"79", x"77", x"77", x"79", x"73", x"75", x"77", x"77", x"77", x"77", x"78", x"78", x"79", 
        x"77", x"76", x"77", x"79", x"78", x"78", x"78", x"79", x"7a", x"7a", x"78", x"78", x"77", x"78", x"79", 
        x"77", x"79", x"7a", x"78", x"79", x"79", x"79", x"79", x"7a", x"7a", x"77", x"77", x"7b", x"7b", x"7a", 
        x"77", x"76", x"78", x"7b", x"79", x"7a", x"7a", x"7a", x"7b", x"7c", x"7b", x"79", x"79", x"7a", x"7b", 
        x"7a", x"7a", x"7a", x"7a", x"79", x"7a", x"7b", x"7b", x"7b", x"7a", x"79", x"79", x"7a", x"7b", x"7c", 
        x"7b", x"79", x"79", x"7c", x"7c", x"7b", x"7a", x"7a", x"7a", x"7a", x"7b", x"7c", x"7d", x"7d", x"7c", 
        x"7c", x"7c", x"7b", x"7b", x"7b", x"7c", x"7b", x"7b", x"7b", x"7b", x"7c", x"7d", x"7d", x"7c", x"7c", 
        x"7d", x"7d", x"7a", x"7b", x"7a", x"79", x"7b", x"7a", x"7e", x"7e", x"7d", x"81", x"80", x"7c", x"7a", 
        x"7a", x"c3", x"d7", x"d3", x"d2", x"d1", x"d5", x"d6", x"cc", x"cc", x"cc", x"cc", x"ce", x"d1", x"cf", 
        x"ce", x"cd", x"cc", x"cc", x"cd", x"ce", x"d0", x"d1", x"d1", x"d1", x"d0", x"d0", x"d0", x"cf", x"d0", 
        x"d0", x"cf", x"d0", x"d0", x"cf", x"cf", x"d0", x"ce", x"cd", x"cd", x"cd", x"ce", x"cf", x"d1", x"cf", 
        x"ce", x"ce", x"cd", x"cc", x"cc", x"cc", x"cb", x"d7", x"dc", x"d1", x"d4", x"d4", x"d4", x"d2", x"cf", 
        x"ba", x"71", x"5c", x"5d", x"5f", x"5f", x"5e", x"5e", x"61", x"9b", x"ec", x"fd", x"fa", x"f4", x"ef", 
        x"f4", x"f8", x"f8", x"f5", x"e9", x"bd", x"6b", x"5e", x"5d", x"5f", x"60", x"92", x"eb", x"fb", x"f8", 
        x"fa", x"f9", x"de", x"86", x"5d", x"5d", x"6e", x"d3", x"e7", x"d9", x"a5", x"6c", x"5c", x"5f", x"60", 
        x"5f", x"5e", x"5e", x"5f", x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5f", x"60", x"61", x"5f", x"5e", x"5e", x"5f", x"5f", x"60", x"60", x"5e", x"5e", x"5d", x"5d", x"5c", 
        x"5c", x"5e", x"5f", x"5f", x"5d", x"5c", x"5d", x"5d", x"5e", x"5e", x"5e", x"5d", x"5b", x"5f", x"67", 
        x"b1", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"f0", x"ef", x"ee", x"ee", x"ee", x"f0", 
        x"f0", x"f0", x"ef", x"f1", x"f2", x"f1", x"ee", x"f0", x"ef", x"ea", x"df", x"c9", x"b5", x"b8", x"c7", 
        x"db", x"e6", x"ed", x"f0", x"f1", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f2", x"f1", x"f0", x"ee", x"f0", x"ec", x"eb", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", 
        x"ef", x"ef", x"f0", x"ee", x"f0", x"f2", x"f3", x"f2", x"ec", x"ef", x"f1", x"f2", x"f1", x"e9", x"df", 
        x"d9", x"d6", x"de", x"e0", x"c9", x"9b", x"7b", x"77", x"7d", x"7f", x"7d", x"7e", x"7d", x"7f", x"81", 
        x"7d", x"79", x"80", x"85", x"84", x"85", x"80", x"83", x"83", x"82", x"80", x"80", x"80", x"80", x"82", 
        x"83", x"80", x"80", x"82", x"83", x"83", x"82", x"82", x"81", x"81", x"81", x"81", x"81", x"81", x"82", 
        x"81", x"81", x"82", x"82", x"80", x"80", x"82", x"83", x"82", x"82", x"82", x"82", x"82", x"82", x"81", 
        x"80", x"81", x"82", x"81", x"81", x"81", x"81", x"83", x"83", x"82", x"81", x"80", x"80", x"80", x"7f", 
        x"80", x"7f", x"7e", x"7f", x"82", x"82", x"81", x"81", x"81", x"81", x"83", x"82", x"7f", x"7d", x"7e", 
        x"7f", x"81", x"80", x"80", x"81", x"82", x"80", x"7f", x"80", x"82", x"81", x"7f", x"80", x"81", x"81", 
        x"81", x"7f", x"7f", x"80", x"81", x"80", x"81", x"80", x"7e", x"7e", x"81", x"81", x"80", x"81", x"81", 
        x"80", x"7f", x"7e", x"80", x"81", x"80", x"81", x"81", x"81", x"80", x"7e", x"7d", x"7e", x"7e", x"7e", 
        x"7e", x"7f", x"80", x"80", x"7d", x"7f", x"7e", x"7d", x"7b", x"7c", x"7e", x"7f", x"7e", x"7e", x"7e", 
        x"7f", x"7e", x"7c", x"7c", x"7b", x"7b", x"7c", x"7d", x"7e", x"7f", x"7c", x"7b", x"7f", x"7e", x"7c", 
        x"7c", x"7c", x"7c", x"7e", x"7d", x"7b", x"7e", x"7e", x"7c", x"7d", x"7b", x"7c", x"7e", x"7e", x"7c", 
        x"7b", x"7a", x"7b", x"7b", x"7c", x"7b", x"7b", x"7c", x"7b", x"7b", x"7b", x"7b", x"7c", x"7c", x"7c", 
        x"7c", x"7d", x"7d", x"7b", x"7b", x"7c", x"7d", x"7c", x"7c", x"7b", x"7b", x"7d", x"7c", x"7c", x"7c", 
        x"7c", x"7b", x"7a", x"7b", x"7c", x"7b", x"7c", x"7e", x"7d", x"7c", x"7b", x"7b", x"7b", x"7b", x"7a", 
        x"7b", x"7d", x"7d", x"7c", x"7a", x"7a", x"7b", x"7c", x"7f", x"7c", x"7e", x"7a", x"7c", x"7b", x"7c", 
        x"79", x"79", x"7b", x"7a", x"7b", x"7d", x"7a", x"7b", x"7c", x"7b", x"7b", x"7a", x"7b", x"7c", x"79", 
        x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", x"7d", x"7c", x"79", x"79", x"7a", x"77", x"77", x"79", 
        x"79", x"79", x"78", x"78", x"78", x"78", x"78", x"75", x"75", x"77", x"78", x"78", x"76", x"75", x"78", 
        x"76", x"77", x"7a", x"77", x"77", x"79", x"79", x"78", x"77", x"78", x"78", x"78", x"79", x"78", x"78", 
        x"78", x"79", x"78", x"75", x"74", x"76", x"74", x"75", x"76", x"76", x"77", x"78", x"7a", x"79", x"79", 
        x"76", x"75", x"78", x"7a", x"78", x"78", x"77", x"78", x"7b", x"7a", x"77", x"78", x"77", x"78", x"79", 
        x"77", x"7a", x"7a", x"77", x"78", x"7a", x"78", x"78", x"79", x"78", x"79", x"78", x"7b", x"79", x"77", 
        x"76", x"77", x"78", x"79", x"7a", x"78", x"79", x"7b", x"7c", x"7b", x"7b", x"78", x"79", x"7b", x"7b", 
        x"79", x"79", x"79", x"78", x"78", x"79", x"7a", x"7a", x"79", x"79", x"79", x"79", x"7b", x"7c", x"7d", 
        x"7b", x"78", x"78", x"7a", x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", x"7c", x"7d", x"7d", x"7b", 
        x"7b", x"7a", x"7d", x"7c", x"7b", x"7c", x"7d", x"7d", x"7d", x"7c", x"7b", x"7c", x"7c", x"7c", x"7e", 
        x"7f", x"80", x"7e", x"7d", x"7c", x"7c", x"7e", x"7e", x"7f", x"7c", x"7c", x"80", x"80", x"7e", x"7c", 
        x"7b", x"c3", x"db", x"d2", x"cf", x"d4", x"d7", x"d6", x"cc", x"cc", x"cd", x"cc", x"ce", x"d0", x"cf", 
        x"ce", x"cd", x"cd", x"cd", x"cd", x"ce", x"cf", x"d1", x"d1", x"d1", x"d0", x"d1", x"d0", x"cf", x"d0", 
        x"d0", x"ce", x"cf", x"cf", x"ce", x"cf", x"d1", x"cf", x"ce", x"cd", x"cc", x"cd", x"cf", x"d0", x"cf", 
        x"d0", x"d0", x"cf", x"cd", x"cc", x"cd", x"cb", x"d6", x"dd", x"d1", x"d5", x"d4", x"d3", x"d2", x"cf", 
        x"bb", x"72", x"5c", x"5d", x"5f", x"5d", x"5d", x"5e", x"61", x"99", x"ea", x"fc", x"fa", x"e3", x"b8", 
        x"c3", x"df", x"ee", x"f6", x"f5", x"d2", x"69", x"5c", x"5e", x"5f", x"5d", x"8f", x"ec", x"fa", x"f9", 
        x"f8", x"f7", x"f0", x"b9", x"6b", x"5f", x"6c", x"d6", x"f4", x"f5", x"c5", x"74", x"5a", x"5f", x"61", 
        x"5f", x"5e", x"5d", x"5c", x"5c", x"5d", x"5d", x"5d", x"5e", x"5e", x"5d", x"5d", x"5e", x"5f", x"5d", 
        x"5d", x"5e", x"5d", x"5e", x"5d", x"5c", x"5d", x"5f", x"5e", x"5c", x"5c", x"5e", x"60", x"60", x"60", 
        x"5f", x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5e", x"5e", x"5e", x"5d", x"5b", x"5e", x"67", 
        x"af", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ed", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"f0", x"f0", x"df", x"c4", 
        x"b2", x"ba", x"cc", x"e1", x"ed", x"f1", x"f1", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", 
        x"f1", x"f1", x"ef", x"ef", x"f0", x"ec", x"ec", x"f0", x"f0", x"f1", x"f2", x"f3", x"f0", x"ef", x"ef", 
        x"ef", x"ee", x"f0", x"f1", x"f4", x"f1", x"ef", x"f2", x"f1", x"f0", x"ee", x"ed", x"f1", x"f3", x"f1", 
        x"f1", x"e8", x"d9", x"d8", x"df", x"e4", x"d6", x"b3", x"89", x"72", x"77", x"7e", x"84", x"83", x"81", 
        x"7e", x"7c", x"7b", x"7f", x"82", x"84", x"81", x"82", x"81", x"82", x"82", x"81", x"7f", x"80", x"81", 
        x"81", x"80", x"80", x"81", x"81", x"82", x"83", x"82", x"83", x"84", x"83", x"82", x"81", x"82", x"81", 
        x"81", x"82", x"83", x"82", x"7f", x"7e", x"7f", x"81", x"82", x"81", x"81", x"81", x"81", x"81", x"81", 
        x"82", x"81", x"81", x"81", x"83", x"83", x"81", x"81", x"80", x"80", x"80", x"80", x"82", x"82", x"81", 
        x"81", x"80", x"7e", x"7f", x"83", x"83", x"81", x"81", x"81", x"81", x"83", x"81", x"7e", x"7d", x"7f", 
        x"7f", x"82", x"80", x"80", x"82", x"81", x"81", x"80", x"81", x"83", x"82", x"81", x"82", x"82", x"81", 
        x"80", x"7e", x"7e", x"7f", x"81", x"80", x"81", x"80", x"7f", x"7f", x"81", x"81", x"81", x"81", x"80", 
        x"7f", x"80", x"81", x"7f", x"7f", x"80", x"81", x"82", x"81", x"80", x"7e", x"7d", x"7f", x"80", x"7f", 
        x"7f", x"7f", x"7e", x"7e", x"7d", x"7f", x"7f", x"7e", x"7c", x"7d", x"7e", x"7e", x"7e", x"7d", x"7d", 
        x"7e", x"7f", x"7b", x"7b", x"7c", x"7c", x"7d", x"7d", x"7c", x"7c", x"7e", x"7e", x"7b", x"7a", x"7c", 
        x"7e", x"7c", x"7a", x"7a", x"7a", x"79", x"7b", x"7c", x"79", x"7a", x"79", x"7b", x"7d", x"7e", x"7d", 
        x"7b", x"7b", x"7b", x"7c", x"7d", x"7b", x"7c", x"7d", x"7b", x"7a", x"7b", x"7c", x"7c", x"7d", x"7d", 
        x"7d", x"7d", x"7b", x"7b", x"7c", x"7d", x"7e", x"7d", x"7c", x"7b", x"7a", x"7d", x"7c", x"7b", x"7d", 
        x"7d", x"7e", x"7c", x"7c", x"7c", x"7b", x"7a", x"7c", x"7e", x"7e", x"7c", x"7a", x"7b", x"7b", x"79", 
        x"78", x"7a", x"7c", x"7c", x"7c", x"7c", x"7e", x"7d", x"7e", x"7d", x"7e", x"7a", x"7b", x"7c", x"7d", 
        x"7a", x"7a", x"7c", x"7b", x"7b", x"7d", x"7a", x"79", x"79", x"79", x"79", x"78", x"79", x"7b", x"7a", 
        x"7b", x"7c", x"7b", x"7a", x"7b", x"7c", x"7b", x"7c", x"7a", x"78", x"79", x"7b", x"7b", x"79", x"79", 
        x"78", x"79", x"77", x"77", x"79", x"78", x"7a", x"78", x"75", x"77", x"79", x"77", x"74", x"76", x"7a", 
        x"79", x"78", x"78", x"75", x"77", x"79", x"78", x"77", x"78", x"79", x"77", x"77", x"78", x"75", x"75", 
        x"77", x"77", x"77", x"76", x"76", x"78", x"73", x"76", x"76", x"77", x"77", x"74", x"78", x"7a", x"7a", 
        x"75", x"76", x"79", x"77", x"78", x"79", x"79", x"79", x"7a", x"79", x"79", x"79", x"77", x"78", x"7a", 
        x"79", x"78", x"78", x"78", x"78", x"79", x"77", x"78", x"7a", x"77", x"78", x"77", x"79", x"79", x"78", 
        x"77", x"77", x"78", x"7a", x"7a", x"79", x"79", x"79", x"7a", x"7a", x"7b", x"79", x"7c", x"7c", x"79", 
        x"7a", x"7d", x"7a", x"79", x"7a", x"7b", x"79", x"78", x"78", x"7a", x"7a", x"79", x"7a", x"7b", x"7c", 
        x"7b", x"7b", x"7b", x"7c", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7c", x"7c", x"7d", x"7b", x"78", 
        x"79", x"79", x"7c", x"7a", x"7a", x"7d", x"7d", x"7c", x"7d", x"7f", x"7f", x"7e", x"7d", x"7e", x"7e", 
        x"7d", x"7c", x"7c", x"7c", x"7d", x"7d", x"7f", x"7d", x"7d", x"7b", x"7c", x"7d", x"7c", x"7f", x"7d", 
        x"7b", x"c1", x"da", x"d2", x"d2", x"d3", x"d6", x"d7", x"cc", x"ce", x"cf", x"ce", x"ce", x"cf", x"ce", 
        x"cc", x"cd", x"d0", x"d0", x"cf", x"ce", x"cf", x"d0", x"cf", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", 
        x"cf", x"cf", x"cf", x"ce", x"ce", x"ce", x"ce", x"ce", x"cd", x"ce", x"ce", x"ce", x"ce", x"cf", x"d0", 
        x"d1", x"d0", x"cf", x"cd", x"cd", x"cd", x"cc", x"d5", x"dc", x"d1", x"d4", x"d1", x"d0", x"d2", x"d0", 
        x"bf", x"74", x"5c", x"5f", x"5f", x"5b", x"5d", x"5e", x"5f", x"96", x"e8", x"fa", x"fb", x"d5", x"7c", 
        x"70", x"89", x"a5", x"c6", x"da", x"c7", x"68", x"5d", x"60", x"61", x"5f", x"8d", x"eb", x"f9", x"f7", 
        x"ed", x"f3", x"f7", x"e3", x"86", x"61", x"70", x"d5", x"f7", x"fc", x"ca", x"76", x"5b", x"5c", x"5e", 
        x"5e", x"5c", x"5c", x"60", x"6b", x"68", x"61", x"5c", x"5b", x"5b", x"5d", x"5e", x"5d", x"5f", x"5c", 
        x"5c", x"63", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5f", x"5f", x"5f", 
        x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5b", x"5d", x"67", 
        x"ab", x"ee", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"f1", x"f1", x"ee", 
        x"e8", x"d6", x"c2", x"bc", x"c6", x"d5", x"e1", x"eb", x"f1", x"f1", x"f0", x"f0", x"ef", x"ee", x"ee", 
        x"f0", x"ef", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"ee", x"f0", x"f1", x"ee", x"ee", x"f0", x"f0", 
        x"ef", x"ee", x"ef", x"f0", x"f0", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"f1", x"f1", x"ed", x"ec", x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"ea", x"e0", x"d8", x"de", x"e1", x"d7", x"b7", x"94", x"7b", x"74", x"7a", x"80", 
        x"82", x"80", x"7e", x"80", x"84", x"84", x"84", x"83", x"81", x"83", x"85", x"85", x"80", x"81", x"82", 
        x"81", x"82", x"82", x"82", x"81", x"82", x"84", x"82", x"82", x"83", x"82", x"82", x"82", x"82", x"82", 
        x"82", x"83", x"82", x"82", x"81", x"81", x"81", x"82", x"83", x"82", x"82", x"82", x"82", x"80", x"7f", 
        x"81", x"80", x"80", x"81", x"82", x"81", x"80", x"81", x"7f", x"82", x"83", x"81", x"82", x"81", x"81", 
        x"82", x"81", x"80", x"80", x"82", x"82", x"82", x"81", x"81", x"81", x"82", x"81", x"7f", x"7e", x"81", 
        x"82", x"82", x"82", x"81", x"80", x"80", x"82", x"81", x"80", x"80", x"80", x"80", x"81", x"80", x"7f", 
        x"80", x"80", x"7f", x"7f", x"7f", x"7e", x"7e", x"7f", x"81", x"82", x"81", x"7f", x"7f", x"81", x"81", 
        x"81", x"81", x"80", x"7e", x"7f", x"82", x"80", x"80", x"81", x"7f", x"7f", x"80", x"7e", x"7e", x"7f", 
        x"7f", x"7f", x"80", x"80", x"81", x"80", x"7f", x"7e", x"7f", x"80", x"82", x"7d", x"7c", x"7c", x"7d", 
        x"7d", x"7d", x"7c", x"7c", x"7b", x"7b", x"7e", x"7e", x"7c", x"7c", x"7d", x"7c", x"7d", x"80", x"7d", 
        x"7c", x"7d", x"7c", x"7c", x"7b", x"7c", x"7c", x"7a", x"7b", x"7d", x"7b", x"7b", x"7b", x"7c", x"7c", 
        x"7c", x"7c", x"7d", x"7c", x"7d", x"7f", x"7e", x"7d", x"7d", x"7d", x"7d", x"7e", x"7d", x"7b", x"7a", 
        x"7a", x"7b", x"7c", x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", x"7d", x"7e", x"7d", x"7a", x"78", x"7a", 
        x"7d", x"7f", x"7c", x"7c", x"7d", x"7b", x"7a", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7b", 
        x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", x"7d", x"7b", x"7b", x"7d", x"7c", x"7b", x"7b", x"7b", x"7c", 
        x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7a", x"7b", x"7d", x"7b", x"7a", x"7b", x"7c", x"7c", 
        x"7c", x"7c", x"7d", x"7a", x"7d", x"7c", x"7a", x"79", x"78", x"78", x"7a", x"7b", x"7a", x"7a", x"7a", 
        x"78", x"7a", x"78", x"78", x"79", x"76", x"77", x"78", x"77", x"77", x"79", x"77", x"74", x"75", x"78", 
        x"79", x"79", x"79", x"78", x"77", x"76", x"76", x"76", x"78", x"7a", x"78", x"78", x"78", x"75", x"76", 
        x"78", x"78", x"79", x"79", x"78", x"7a", x"75", x"77", x"77", x"79", x"79", x"76", x"77", x"79", x"79", 
        x"76", x"77", x"7a", x"78", x"79", x"79", x"79", x"79", x"7a", x"7a", x"7a", x"7b", x"78", x"77", x"7a", 
        x"7b", x"7b", x"79", x"78", x"78", x"78", x"76", x"78", x"7a", x"77", x"78", x"77", x"79", x"78", x"77", 
        x"78", x"79", x"79", x"79", x"7a", x"7a", x"7a", x"7a", x"7a", x"7b", x"7b", x"7a", x"7d", x"7c", x"79", 
        x"7b", x"7d", x"7a", x"79", x"7b", x"7b", x"7b", x"7a", x"7b", x"7d", x"7b", x"79", x"79", x"7b", x"7c", 
        x"7d", x"7d", x"7c", x"7a", x"7d", x"7d", x"7c", x"7a", x"7c", x"7e", x"7d", x"7c", x"7e", x"7b", x"78", 
        x"7a", x"7a", x"7d", x"7b", x"7b", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7c", x"7d", x"7d", 
        x"7c", x"7c", x"7d", x"7d", x"7e", x"7e", x"7e", x"7d", x"7d", x"7c", x"7d", x"7e", x"7c", x"80", x"7e", 
        x"78", x"c4", x"dd", x"d5", x"d4", x"d3", x"d6", x"d6", x"cd", x"ce", x"cf", x"cd", x"cd", x"cf", x"ce", 
        x"ce", x"ce", x"d0", x"d0", x"ce", x"cd", x"ce", x"d0", x"d0", x"cf", x"cf", x"cf", x"d0", x"d0", x"d0", 
        x"d0", x"cf", x"ce", x"ce", x"ce", x"cf", x"cf", x"ce", x"ce", x"cf", x"cf", x"d0", x"d1", x"d1", x"d1", 
        x"d2", x"d0", x"cf", x"cd", x"cc", x"cc", x"cb", x"d5", x"dc", x"d1", x"d3", x"d1", x"d0", x"d2", x"d4", 
        x"c1", x"75", x"5d", x"5e", x"5f", x"5e", x"5e", x"5f", x"5f", x"96", x"e9", x"fa", x"fa", x"d7", x"7d", 
        x"5f", x"5d", x"5d", x"71", x"8a", x"93", x"66", x"5e", x"5e", x"61", x"5f", x"89", x"ea", x"fb", x"f5", 
        x"d4", x"db", x"f9", x"f7", x"b5", x"6c", x"6d", x"d7", x"f9", x"fd", x"ce", x"79", x"5f", x"5c", x"5f", 
        x"5c", x"5d", x"7d", x"9c", x"af", x"a9", x"97", x"83", x"6b", x"5c", x"5b", x"5c", x"5e", x"60", x"5e", 
        x"5e", x"5e", x"5d", x"5c", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5f", x"5f", x"5f", x"5f", x"5f", 
        x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5c", x"5c", x"66", 
        x"a7", x"eb", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", 
        x"f0", x"f0", x"ee", x"df", x"ca", x"be", x"bf", x"ca", x"d7", x"e4", x"ef", x"f1", x"ef", x"ee", x"ef", 
        x"ee", x"ed", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"f0", x"ee", x"ee", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"f0", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"ed", x"ec", x"f0", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"ec", x"e2", x"d9", x"dd", x"de", x"d7", x"bc", x"94", x"80", x"77", 
        x"76", x"7e", x"82", x"83", x"7e", x"80", x"84", x"82", x"86", x"87", x"85", x"84", x"83", x"82", x"82", 
        x"81", x"82", x"82", x"82", x"83", x"84", x"83", x"84", x"83", x"82", x"82", x"83", x"84", x"83", x"81", 
        x"82", x"85", x"84", x"83", x"83", x"83", x"83", x"83", x"82", x"81", x"82", x"83", x"82", x"80", x"7f", 
        x"81", x"81", x"81", x"81", x"81", x"81", x"80", x"80", x"7e", x"81", x"82", x"81", x"83", x"82", x"81", 
        x"82", x"82", x"81", x"81", x"82", x"82", x"82", x"82", x"82", x"83", x"84", x"84", x"84", x"82", x"81", 
        x"81", x"81", x"81", x"82", x"82", x"82", x"82", x"82", x"81", x"80", x"7e", x"7e", x"7e", x"80", x"81", 
        x"81", x"81", x"81", x"81", x"80", x"80", x"80", x"80", x"80", x"80", x"81", x"80", x"80", x"81", x"82", 
        x"82", x"81", x"80", x"7f", x"7f", x"80", x"7f", x"81", x"81", x"80", x"7f", x"80", x"80", x"80", x"80", 
        x"80", x"80", x"81", x"80", x"7f", x"7f", x"7f", x"7f", x"7f", x"81", x"82", x"7e", x"7e", x"7f", x"7e", 
        x"7d", x"7c", x"7d", x"7e", x"7d", x"7c", x"7d", x"7e", x"7d", x"7e", x"7d", x"7d", x"7f", x"80", x"7d", 
        x"7e", x"7f", x"7d", x"7e", x"7c", x"7d", x"7c", x"7b", x"7c", x"7f", x"7d", x"7e", x"7e", x"7c", x"7b", 
        x"7b", x"7b", x"7e", x"7e", x"7e", x"80", x"7f", x"7d", x"7f", x"7e", x"7f", x"7f", x"7e", x"7c", x"7b", 
        x"7b", x"7d", x"7e", x"7c", x"7d", x"7e", x"7f", x"7d", x"7b", x"7d", x"7e", x"7d", x"7b", x"79", x"7b", 
        x"7d", x"7d", x"7c", x"7c", x"7e", x"7d", x"7d", x"7f", x"7c", x"7c", x"7c", x"7d", x"7e", x"7d", x"7c", 
        x"7c", x"7b", x"7b", x"7d", x"7e", x"7e", x"7d", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7c", 
        x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7d", x"7b", x"7a", x"7b", x"7b", x"7c", 
        x"7a", x"7c", x"7b", x"7a", x"7c", x"7b", x"7a", x"7a", x"7b", x"7b", x"7c", x"7b", x"79", x"7a", x"7b", 
        x"77", x"79", x"78", x"79", x"7a", x"77", x"77", x"79", x"79", x"78", x"79", x"79", x"77", x"76", x"75", 
        x"78", x"78", x"78", x"7a", x"78", x"76", x"77", x"76", x"78", x"7b", x"7a", x"7a", x"79", x"77", x"78", 
        x"78", x"76", x"77", x"77", x"75", x"77", x"77", x"78", x"78", x"7a", x"7b", x"78", x"77", x"77", x"79", 
        x"77", x"79", x"7c", x"7a", x"7a", x"7a", x"7a", x"7a", x"7a", x"7a", x"7a", x"7a", x"79", x"79", x"79", 
        x"7a", x"79", x"79", x"79", x"79", x"78", x"77", x"79", x"7a", x"78", x"78", x"78", x"7b", x"7b", x"7a", 
        x"7a", x"79", x"78", x"78", x"7a", x"7a", x"7a", x"7a", x"7a", x"7b", x"7c", x"7a", x"7c", x"7c", x"7a", 
        x"7b", x"7c", x"7a", x"79", x"7a", x"7a", x"7a", x"79", x"79", x"7a", x"7a", x"79", x"7a", x"7a", x"7c", 
        x"7d", x"7e", x"7e", x"7c", x"7c", x"7c", x"7c", x"7c", x"7d", x"7d", x"7d", x"7c", x"7e", x"7d", x"7a", 
        x"7c", x"7a", x"7c", x"7b", x"7b", x"7c", x"7c", x"7c", x"7c", x"7e", x"7e", x"7d", x"7d", x"7d", x"7e", 
        x"7d", x"7f", x"80", x"7f", x"7f", x"7f", x"7f", x"7e", x"7d", x"7d", x"7f", x"7f", x"7e", x"7d", x"79", 
        x"79", x"c1", x"db", x"d2", x"d1", x"d1", x"d7", x"d7", x"cd", x"ce", x"cf", x"cd", x"cd", x"cf", x"cf", 
        x"cd", x"ce", x"cf", x"d0", x"cf", x"d0", x"d1", x"d1", x"d1", x"cf", x"ce", x"cf", x"d0", x"d1", x"d1", 
        x"d0", x"cf", x"ce", x"ce", x"ce", x"cf", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", 
        x"d1", x"d0", x"ce", x"cc", x"cc", x"cc", x"cb", x"cf", x"dd", x"d2", x"d3", x"cf", x"d5", x"de", x"be", 
        x"9b", x"69", x"58", x"5a", x"5e", x"5d", x"5d", x"60", x"5d", x"90", x"e7", x"f8", x"f8", x"d9", x"7d", 
        x"57", x"59", x"5e", x"5e", x"5e", x"5e", x"5f", x"5d", x"5b", x"5d", x"61", x"88", x"e7", x"fd", x"f4", 
        x"be", x"b4", x"eb", x"fa", x"e0", x"8c", x"6d", x"d6", x"f8", x"fa", x"d0", x"7d", x"60", x"60", x"60", 
        x"5f", x"8b", x"d0", x"ee", x"f5", x"f3", x"f0", x"e2", x"be", x"97", x"6b", x"5a", x"5b", x"61", x"5f", 
        x"5f", x"5f", x"5d", x"5d", x"5e", x"5f", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5e", x"5d", x"5d", x"64", 
        x"a2", x"e9", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", 
        x"f0", x"ef", x"ed", x"ef", x"f2", x"ec", x"dc", x"c9", x"be", x"bf", x"ca", x"da", x"e9", x"f1", x"f2", 
        x"f0", x"ed", x"ee", x"f0", x"ef", x"ee", x"ed", x"ee", x"ed", x"ed", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f1", x"f0", x"f0", x"f1", x"f2", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"ed", x"ec", x"f0", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", 
        x"f1", x"f0", x"f2", x"f1", x"f0", x"f3", x"f4", x"ec", x"e5", x"da", x"d6", x"de", x"df", x"cd", x"aa", 
        x"85", x"73", x"71", x"78", x"80", x"86", x"87", x"87", x"87", x"85", x"85", x"83", x"86", x"83", x"82", 
        x"81", x"82", x"82", x"83", x"85", x"84", x"82", x"84", x"84", x"82", x"82", x"83", x"84", x"83", x"81", 
        x"82", x"84", x"83", x"82", x"82", x"82", x"83", x"83", x"82", x"81", x"81", x"83", x"83", x"82", x"80", 
        x"81", x"82", x"82", x"81", x"80", x"81", x"82", x"81", x"80", x"81", x"82", x"82", x"83", x"83", x"83", 
        x"82", x"82", x"81", x"81", x"82", x"82", x"81", x"80", x"82", x"82", x"82", x"82", x"82", x"83", x"81", 
        x"81", x"80", x"80", x"81", x"82", x"83", x"83", x"82", x"82", x"82", x"81", x"80", x"80", x"81", x"82", 
        x"81", x"81", x"81", x"82", x"82", x"82", x"82", x"81", x"80", x"7e", x"7f", x"80", x"82", x"82", x"82", 
        x"82", x"81", x"80", x"7f", x"7f", x"7e", x"7e", x"80", x"82", x"80", x"7e", x"80", x"82", x"81", x"80", 
        x"80", x"80", x"80", x"80", x"7d", x"7e", x"80", x"80", x"7f", x"7f", x"82", x"7d", x"7d", x"7e", x"7d", 
        x"7a", x"7a", x"7b", x"80", x"7e", x"7b", x"7c", x"7e", x"7d", x"7d", x"7c", x"7b", x"7d", x"7d", x"7a", 
        x"7d", x"7e", x"7b", x"7c", x"7d", x"7f", x"7f", x"7d", x"7c", x"7d", x"7d", x"7f", x"80", x"7f", x"7f", 
        x"81", x"82", x"80", x"7e", x"7d", x"7e", x"7d", x"7c", x"7d", x"7e", x"7f", x"7f", x"7e", x"7d", x"7d", 
        x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7d", x"7d", x"7b", x"7a", x"7b", 
        x"7e", x"7d", x"7d", x"7d", x"7e", x"7f", x"80", x"80", x"7c", x"7b", x"7b", x"7d", x"7e", x"7e", x"7c", 
        x"7c", x"7c", x"7d", x"7d", x"7e", x"7d", x"7c", x"7c", x"7b", x"7a", x"7a", x"7c", x"7d", x"7d", x"7c", 
        x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7a", x"7b", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", 
        x"79", x"7c", x"7a", x"7b", x"7b", x"7b", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7a", x"7b", x"7c", 
        x"7a", x"7b", x"78", x"77", x"78", x"76", x"76", x"78", x"77", x"77", x"78", x"79", x"79", x"77", x"76", 
        x"7a", x"79", x"78", x"7a", x"77", x"76", x"78", x"78", x"78", x"79", x"79", x"7a", x"7a", x"79", x"78", 
        x"78", x"76", x"78", x"78", x"76", x"78", x"78", x"77", x"78", x"79", x"79", x"78", x"76", x"77", x"7a", 
        x"79", x"7a", x"7c", x"79", x"7a", x"7a", x"7a", x"7a", x"79", x"79", x"78", x"78", x"7a", x"7a", x"79", 
        x"78", x"78", x"79", x"7a", x"7b", x"79", x"79", x"7a", x"7a", x"79", x"78", x"79", x"78", x"79", x"7a", 
        x"79", x"78", x"79", x"7a", x"7a", x"79", x"79", x"79", x"79", x"7b", x"7b", x"79", x"7b", x"7b", x"7b", 
        x"7c", x"7d", x"7c", x"7b", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7a", x"7a", x"7b", x"7c", x"7d", 
        x"7d", x"7c", x"7d", x"7e", x"7b", x"7b", x"7d", x"7e", x"7c", x"7b", x"7d", x"7c", x"7e", x"7d", x"7c", 
        x"7d", x"7b", x"7d", x"7e", x"7d", x"7e", x"7e", x"7e", x"7d", x"7e", x"7f", x"7f", x"7f", x"7f", x"7f", 
        x"7f", x"80", x"80", x"7f", x"80", x"81", x"80", x"7f", x"7d", x"7d", x"82", x"80", x"7f", x"80", x"7d", 
        x"7b", x"c0", x"dc", x"d2", x"d1", x"d1", x"d8", x"d7", x"cd", x"cf", x"d0", x"ce", x"ce", x"cf", x"cf", 
        x"cf", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", 
        x"d1", x"d0", x"cf", x"ce", x"ce", x"cf", x"cf", x"ce", x"ce", x"cf", x"cf", x"d0", x"d0", x"d0", x"d0", 
        x"d1", x"d1", x"cf", x"cd", x"cc", x"cd", x"cc", x"d3", x"d9", x"cf", x"d6", x"d4", x"ce", x"a8", x"90", 
        x"a4", x"a7", x"8e", x"74", x"62", x"5a", x"5c", x"60", x"5c", x"8d", x"e5", x"f9", x"f7", x"e5", x"ad", 
        x"82", x"6b", x"61", x"5f", x"5d", x"5b", x"5e", x"60", x"5d", x"5e", x"60", x"85", x"e7", x"fd", x"f6", 
        x"bf", x"90", x"cd", x"f8", x"f2", x"ba", x"7c", x"cc", x"f7", x"f9", x"d3", x"7e", x"5b", x"61", x"5e", 
        x"6b", x"c0", x"f1", x"f5", x"f8", x"f9", x"f6", x"f6", x"f3", x"e2", x"be", x"8a", x"68", x"5c", x"5d", 
        x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5c", x"5b", x"5d", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5d", x"5d", x"5d", x"63", 
        x"9d", x"e8", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ed", 
        x"eb", x"ed", x"f0", x"ee", x"ec", x"ee", x"f0", x"ef", x"e7", x"da", x"ca", x"c2", x"c4", x"d0", x"de", 
        x"ec", x"f0", x"f1", x"f0", x"ee", x"ed", x"ed", x"ef", x"ee", x"ed", x"ee", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f1", x"f0", x"f0", x"f1", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"ed", x"ec", x"f0", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f3", x"f1", x"f1", x"ed", x"ec", x"ea", x"e6", x"dd", x"db", x"db", x"de", 
        x"d1", x"b8", x"96", x"76", x"73", x"7d", x"83", x"85", x"83", x"80", x"84", x"84", x"83", x"81", x"82", 
        x"80", x"81", x"83", x"84", x"83", x"81", x"81", x"82", x"84", x"84", x"83", x"83", x"83", x"83", x"81", 
        x"82", x"83", x"82", x"82", x"82", x"81", x"82", x"82", x"82", x"81", x"81", x"82", x"83", x"83", x"82", 
        x"82", x"83", x"83", x"81", x"81", x"81", x"83", x"83", x"82", x"82", x"82", x"82", x"82", x"82", x"83", 
        x"83", x"82", x"82", x"82", x"82", x"83", x"82", x"82", x"83", x"83", x"82", x"81", x"82", x"83", x"83", 
        x"82", x"81", x"80", x"81", x"82", x"82", x"80", x"7f", x"7f", x"80", x"81", x"82", x"82", x"82", x"81", 
        x"80", x"80", x"80", x"81", x"82", x"81", x"82", x"82", x"81", x"7f", x"7f", x"80", x"81", x"82", x"81", 
        x"81", x"81", x"81", x"80", x"80", x"80", x"7e", x"7f", x"80", x"7e", x"7e", x"80", x"81", x"80", x"80", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"80", x"81", x"7f", x"7d", x"7e", x"80", x"7c", x"7e", x"7f", x"7f", 
        x"7c", x"7d", x"7e", x"80", x"7d", x"7a", x"7c", x"7e", x"7d", x"7b", x"7c", x"7d", x"7c", x"7e", x"7d", 
        x"7e", x"7f", x"7c", x"7a", x"7c", x"7f", x"81", x"7d", x"7b", x"7b", x"7b", x"7e", x"7f", x"7e", x"7d", 
        x"7e", x"81", x"80", x"7d", x"7c", x"7d", x"7c", x"7b", x"7d", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", 
        x"7d", x"7b", x"7c", x"7d", x"7d", x"7b", x"7b", x"7c", x"7c", x"7b", x"7c", x"7d", x"7c", x"7c", x"7d", 
        x"7e", x"7e", x"7f", x"7e", x"7e", x"7f", x"80", x"80", x"7d", x"7c", x"7c", x"7d", x"7e", x"7d", x"7b", 
        x"7d", x"7e", x"7d", x"7d", x"7c", x"7c", x"7c", x"7d", x"7d", x"7b", x"7c", x"7d", x"7d", x"7b", x"7b", 
        x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", x"7a", x"7b", x"7c", 
        x"7a", x"7c", x"7a", x"7b", x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7d", x"7c", 
        x"7b", x"7c", x"78", x"76", x"78", x"76", x"77", x"77", x"77", x"77", x"78", x"7a", x"7b", x"79", x"78", 
        x"7a", x"79", x"77", x"78", x"77", x"76", x"78", x"78", x"78", x"77", x"79", x"7a", x"79", x"79", x"77", 
        x"78", x"77", x"79", x"79", x"77", x"7a", x"78", x"76", x"77", x"78", x"78", x"78", x"76", x"78", x"7a", 
        x"79", x"79", x"7b", x"79", x"79", x"7a", x"79", x"79", x"79", x"79", x"79", x"79", x"7a", x"7a", x"79", 
        x"79", x"7a", x"7b", x"7a", x"7a", x"79", x"79", x"7b", x"7a", x"79", x"78", x"7b", x"7c", x"7b", x"7a", 
        x"7b", x"7a", x"7a", x"7a", x"79", x"79", x"79", x"79", x"79", x"7a", x"7a", x"79", x"7a", x"7b", x"7b", 
        x"7c", x"7d", x"7d", x"7b", x"7b", x"7b", x"7c", x"7d", x"7d", x"7c", x"7b", x"7b", x"7c", x"7e", x"7e", 
        x"7d", x"7c", x"7c", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7e", x"7d", x"7b", x"7d", x"7d", x"7c", 
        x"7e", x"7b", x"7e", x"7f", x"7e", x"7d", x"7f", x"80", x"7e", x"7d", x"7d", x"7f", x"7e", x"7e", x"7e", 
        x"7f", x"7f", x"7f", x"7f", x"80", x"81", x"81", x"80", x"7f", x"7e", x"82", x"83", x"7f", x"85", x"83", 
        x"75", x"bc", x"db", x"d4", x"d2", x"d2", x"d8", x"d5", x"cc", x"cf", x"d1", x"d0", x"cf", x"d0", x"ce", 
        x"cf", x"d1", x"d1", x"d0", x"d0", x"d0", x"d1", x"d0", x"cf", x"d1", x"d1", x"d0", x"d0", x"d0", x"d0", 
        x"d0", x"d0", x"cf", x"cf", x"cf", x"cf", x"ce", x"cd", x"cd", x"ce", x"ce", x"cf", x"cf", x"d0", x"d0", 
        x"d1", x"d1", x"d0", x"ce", x"cd", x"ce", x"cf", x"d1", x"db", x"d0", x"dc", x"be", x"8f", x"92", x"b1", 
        x"db", x"eb", x"dd", x"c6", x"a8", x"87", x"70", x"60", x"56", x"87", x"df", x"fa", x"f8", x"f5", x"e8", 
        x"d4", x"bd", x"a0", x"80", x"69", x"5d", x"59", x"5f", x"5f", x"5c", x"60", x"88", x"e9", x"fe", x"f8", 
        x"c1", x"70", x"a5", x"f0", x"f9", x"e0", x"96", x"c3", x"f6", x"fa", x"d3", x"7d", x"5b", x"61", x"5d", 
        x"78", x"db", x"f8", x"f6", x"f6", x"e2", x"d6", x"e0", x"f3", x"f7", x"f2", x"d6", x"9a", x"66", x"5e", 
        x"60", x"5b", x"5e", x"60", x"5e", x"5d", x"5d", x"5d", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5e", x"5d", x"5d", x"5d", x"63", 
        x"9a", x"e9", x"f1", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ef", x"ee", x"ec", x"ee", x"ef", x"f0", x"f1", x"f2", x"ed", x"e3", x"d5", x"c7", x"bf", 
        x"c1", x"d4", x"e7", x"f0", x"f2", x"f1", x"f1", x"f0", x"f0", x"ef", x"ee", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f1", x"ed", x"ec", x"f0", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"ee", x"f0", x"ec", x"ed", x"ed", x"ee", x"f0", x"e4", x"d8", x"d6", 
        x"da", x"de", x"db", x"bc", x"95", x"7c", x"73", x"79", x"83", x"85", x"89", x"86", x"83", x"81", x"84", 
        x"83", x"82", x"84", x"85", x"81", x"80", x"81", x"81", x"82", x"83", x"82", x"83", x"84", x"84", x"83", 
        x"83", x"84", x"84", x"84", x"84", x"83", x"83", x"83", x"84", x"82", x"81", x"81", x"83", x"83", x"82", 
        x"83", x"84", x"83", x"82", x"82", x"83", x"84", x"84", x"84", x"83", x"81", x"82", x"82", x"82", x"83", 
        x"83", x"82", x"82", x"82", x"82", x"83", x"82", x"81", x"82", x"82", x"82", x"82", x"83", x"84", x"83", 
        x"82", x"81", x"80", x"80", x"81", x"81", x"80", x"7f", x"7f", x"7f", x"80", x"81", x"81", x"81", x"81", 
        x"7f", x"7f", x"7f", x"80", x"81", x"80", x"81", x"82", x"82", x"81", x"80", x"80", x"81", x"82", x"81", 
        x"81", x"81", x"81", x"81", x"82", x"82", x"7f", x"7f", x"7f", x"7e", x"7e", x"7f", x"80", x"80", x"7f", 
        x"7f", x"7f", x"7f", x"7f", x"81", x"82", x"81", x"7e", x"7c", x"7e", x"80", x"7c", x"7d", x"7f", x"7f", 
        x"7e", x"7e", x"7f", x"7f", x"7d", x"7b", x"7e", x"80", x"7d", x"7b", x"7e", x"7e", x"7b", x"7f", x"7e", 
        x"7e", x"7f", x"7d", x"7c", x"7d", x"7f", x"80", x"7d", x"7c", x"7d", x"7c", x"7d", x"7e", x"7d", x"7b", 
        x"7b", x"7d", x"80", x"7e", x"7e", x"80", x"7f", x"7e", x"7f", x"7e", x"7d", x"7d", x"7d", x"7e", x"7e", 
        x"7d", x"7d", x"7e", x"7d", x"7e", x"7e", x"7f", x"7e", x"7d", x"7c", x"7d", x"7e", x"7e", x"7e", x"7f", 
        x"7f", x"7f", x"7f", x"7e", x"7d", x"7e", x"7f", x"7e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7b", 
        x"7c", x"7d", x"7d", x"7c", x"7c", x"7c", x"7e", x"7c", x"7b", x"7b", x"7c", x"7e", x"7e", x"7d", x"7c", 
        x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7b", x"7b", 
        x"7b", x"7b", x"7a", x"7c", x"7a", x"7b", x"78", x"79", x"7b", x"7b", x"7b", x"7a", x"7a", x"7d", x"7d", 
        x"79", x"7a", x"78", x"79", x"7b", x"79", x"7b", x"77", x"78", x"79", x"78", x"78", x"7a", x"78", x"78", 
        x"77", x"78", x"77", x"77", x"78", x"79", x"78", x"79", x"78", x"77", x"7a", x"79", x"77", x"79", x"7a", 
        x"7c", x"7b", x"7b", x"7a", x"79", x"7b", x"77", x"76", x"78", x"77", x"76", x"7a", x"78", x"78", x"7a", 
        x"78", x"78", x"7a", x"79", x"7b", x"7b", x"79", x"79", x"7a", x"7a", x"7b", x"7b", x"7a", x"7a", x"7a", 
        x"7a", x"7b", x"7b", x"7a", x"7a", x"79", x"7b", x"7d", x"7b", x"7b", x"79", x"7c", x"7a", x"78", x"78", 
        x"79", x"7b", x"7b", x"7a", x"7b", x"7a", x"7a", x"7a", x"7b", x"7c", x"7c", x"7c", x"7c", x"7b", x"7b", 
        x"7b", x"7c", x"7d", x"79", x"78", x"78", x"79", x"7b", x"7b", x"7a", x"7a", x"7b", x"7c", x"7d", x"7d", 
        x"7e", x"7d", x"7b", x"7b", x"7d", x"7e", x"7d", x"7c", x"7e", x"80", x"7e", x"7b", x"7c", x"7c", x"7c", 
        x"7e", x"7c", x"7d", x"7e", x"7e", x"7c", x"7e", x"7e", x"7c", x"7b", x"7d", x"7e", x"7e", x"7e", x"7e", 
        x"7f", x"7f", x"7e", x"7e", x"7f", x"82", x"82", x"81", x"82", x"82", x"80", x"7e", x"82", x"88", x"74", 
        x"5d", x"b7", x"d9", x"d2", x"d1", x"d0", x"d9", x"d5", x"cc", x"cf", x"d1", x"cf", x"cf", x"d0", x"cf", 
        x"cf", x"d0", x"d0", x"d0", x"d0", x"d1", x"d3", x"d1", x"cf", x"d1", x"d1", x"d0", x"cf", x"d0", x"d0", 
        x"cf", x"d0", x"d1", x"d0", x"cf", x"cf", x"ce", x"ce", x"cf", x"cf", x"cf", x"ce", x"ce", x"cf", x"d1", 
        x"d2", x"d1", x"d0", x"cf", x"cf", x"cf", x"ce", x"d1", x"e2", x"ca", x"9b", x"87", x"aa", x"ce", x"d3", 
        x"dd", x"eb", x"f0", x"f0", x"e9", x"e2", x"ce", x"af", x"8b", x"91", x"c5", x"e7", x"f4", x"f7", x"fa", 
        x"f7", x"f4", x"ea", x"d9", x"c2", x"9f", x"76", x"5d", x"5c", x"5c", x"60", x"83", x"e5", x"fd", x"f9", 
        x"c5", x"69", x"81", x"dc", x"f9", x"f3", x"c3", x"cd", x"f5", x"f9", x"d2", x"7d", x"5c", x"5e", x"5f", 
        x"7e", x"e0", x"f7", x"f7", x"e7", x"96", x"73", x"82", x"aa", x"d5", x"f0", x"f5", x"c5", x"76", x"5c", 
        x"60", x"5e", x"66", x"76", x"69", x"5a", x"59", x"5f", x"62", x"5f", x"5e", x"5e", x"5e", x"5e", x"5e", 
        x"5e", x"5e", x"5d", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5e", x"5d", x"5d", x"5d", x"64", 
        x"99", x"e9", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", 
        x"ed", x"ee", x"f0", x"f0", x"ee", x"ee", x"f0", x"f3", x"f2", x"f0", x"ef", x"ef", x"ef", x"ea", x"e4", 
        x"d3", x"bd", x"b8", x"c7", x"dd", x"ec", x"f2", x"f1", x"f3", x"f1", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"f0", x"ef", x"ed", x"ed", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"ed", x"ec", x"f0", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"e9", x"e8", x"ec", x"ee", x"ed", x"e9", x"eb", x"e8", 
        x"e0", x"de", x"d6", x"e0", x"dd", x"cb", x"a8", x"82", x"71", x"7f", x"82", x"83", x"85", x"87", x"86", 
        x"87", x"84", x"83", x"84", x"83", x"83", x"84", x"83", x"84", x"85", x"83", x"84", x"84", x"84", x"82", 
        x"83", x"84", x"85", x"85", x"85", x"84", x"83", x"83", x"84", x"83", x"83", x"83", x"83", x"82", x"81", 
        x"83", x"83", x"83", x"84", x"84", x"84", x"83", x"83", x"85", x"82", x"81", x"83", x"82", x"84", x"84", 
        x"83", x"83", x"82", x"82", x"83", x"83", x"83", x"81", x"80", x"80", x"80", x"82", x"82", x"82", x"82", 
        x"82", x"82", x"81", x"81", x"81", x"81", x"82", x"82", x"82", x"82", x"81", x"80", x"80", x"82", x"81", 
        x"80", x"7f", x"80", x"81", x"82", x"80", x"81", x"81", x"82", x"83", x"82", x"80", x"81", x"82", x"81", 
        x"81", x"81", x"81", x"82", x"83", x"81", x"80", x"80", x"80", x"7e", x"7e", x"80", x"80", x"80", x"7f", 
        x"7f", x"7f", x"80", x"80", x"81", x"82", x"81", x"80", x"7e", x"7e", x"7f", x"7c", x"7c", x"7d", x"7d", 
        x"7d", x"7c", x"7d", x"7e", x"7d", x"7c", x"7e", x"7f", x"7e", x"7d", x"7f", x"7d", x"7a", x"7c", x"7b", 
        x"7c", x"7d", x"7c", x"7e", x"7e", x"80", x"7f", x"7d", x"7d", x"7f", x"7e", x"7e", x"7f", x"7f", x"7e", 
        x"7f", x"80", x"80", x"7e", x"7f", x"81", x"80", x"7f", x"80", x"7f", x"7e", x"7d", x"7d", x"7f", x"7f", 
        x"7e", x"7f", x"80", x"7e", x"7e", x"81", x"81", x"80", x"7e", x"7d", x"7e", x"7f", x"7f", x"7f", x"7e", 
        x"7e", x"7e", x"7f", x"7d", x"7b", x"7c", x"7d", x"7c", x"7c", x"7e", x"7f", x"7f", x"7d", x"7d", x"7d", 
        x"7c", x"7c", x"7d", x"7c", x"7c", x"7d", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", 
        x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7d", x"7e", x"7d", x"7c", x"7b", 
        x"7c", x"7a", x"7b", x"7c", x"7b", x"7c", x"78", x"79", x"7b", x"7b", x"7a", x"7a", x"7a", x"7c", x"7d", 
        x"7a", x"7b", x"7b", x"7b", x"7c", x"79", x"7a", x"77", x"79", x"7b", x"78", x"78", x"79", x"78", x"79", 
        x"78", x"79", x"79", x"77", x"78", x"78", x"76", x"78", x"79", x"78", x"7b", x"79", x"76", x"77", x"76", 
        x"79", x"79", x"79", x"79", x"79", x"7c", x"79", x"77", x"79", x"77", x"76", x"7b", x"7b", x"78", x"7a", 
        x"78", x"78", x"7a", x"7a", x"7d", x"7d", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7c", x"7b", x"79", 
        x"78", x"79", x"7b", x"7b", x"7b", x"7a", x"7b", x"7e", x"7c", x"7c", x"7a", x"7d", x"7b", x"7b", x"7b", 
        x"7a", x"7a", x"7b", x"7c", x"7c", x"7b", x"7b", x"7b", x"7c", x"7c", x"7d", x"7f", x"7e", x"7c", x"7b", 
        x"7b", x"7b", x"7c", x"7b", x"7a", x"7a", x"7a", x"7c", x"7b", x"79", x"79", x"7a", x"7b", x"7c", x"7d", 
        x"7e", x"7e", x"7d", x"7c", x"7b", x"7b", x"7e", x"80", x"80", x"80", x"7e", x"7b", x"7c", x"7c", x"7d", 
        x"7e", x"7c", x"7f", x"80", x"7f", x"7d", x"7f", x"80", x"7d", x"7c", x"7e", x"80", x"80", x"7f", x"80", 
        x"81", x"7f", x"7c", x"7d", x"7f", x"82", x"83", x"82", x"81", x"82", x"80", x"83", x"84", x"67", x"51", 
        x"61", x"be", x"dd", x"d3", x"d0", x"d0", x"da", x"d7", x"cd", x"cf", x"d0", x"ce", x"ce", x"d0", x"d0", 
        x"d1", x"d1", x"d1", x"d0", x"d0", x"d1", x"d2", x"d1", x"d0", x"d0", x"d0", x"cf", x"cf", x"d1", x"d1", 
        x"cf", x"d1", x"d2", x"d1", x"d0", x"cf", x"ce", x"ce", x"cf", x"cf", x"cf", x"d0", x"d0", x"d1", x"d2", 
        x"d3", x"d2", x"d0", x"cf", x"cf", x"d0", x"ce", x"d7", x"c6", x"8f", x"9d", x"c4", x"d5", x"d7", x"d1", 
        x"dc", x"ed", x"e9", x"ec", x"ed", x"ee", x"ed", x"eb", x"e2", x"d3", x"ce", x"c2", x"c4", x"d3", x"e6", 
        x"f0", x"f5", x"f8", x"f9", x"f4", x"e4", x"a1", x"64", x"5c", x"5d", x"62", x"81", x"e2", x"fb", x"f8", 
        x"c6", x"6b", x"64", x"b2", x"f1", x"f8", x"ec", x"e6", x"f8", x"fa", x"d4", x"7c", x"5a", x"5f", x"5e", 
        x"6f", x"ce", x"f8", x"f7", x"e8", x"90", x"61", x"60", x"63", x"7f", x"b7", x"ed", x"cc", x"7c", x"5c", 
        x"5b", x"5e", x"77", x"c8", x"bf", x"a1", x"80", x"6b", x"62", x"5f", x"5d", x"5d", x"5d", x"5e", x"5d", 
        x"5c", x"5d", x"5e", x"5d", x"5d", x"5d", x"5e", x"5e", x"5e", x"5e", x"5f", x"5d", x"5d", x"5d", x"63", 
        x"97", x"e9", x"ef", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ec", x"ee", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ed", x"e9", x"df", x"c9", x"b3", x"bb", x"d1", x"e2", x"ec", x"f0", x"f0", x"ef", x"f0", x"ef", x"ee", 
        x"ef", x"f0", x"ee", x"ed", x"ed", x"ee", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"ed", x"ec", x"f0", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f2", x"f4", x"f0", x"f1", x"ec", x"ea", x"eb", x"eb", x"eb", x"ed", x"ed", x"ed", 
        x"ee", x"eb", x"e6", x"e0", x"d9", x"da", x"e2", x"d4", x"b3", x"8b", x"75", x"74", x"7c", x"87", x"86", 
        x"86", x"86", x"82", x"82", x"84", x"85", x"85", x"85", x"86", x"86", x"83", x"81", x"82", x"84", x"85", 
        x"83", x"82", x"83", x"84", x"85", x"83", x"82", x"82", x"83", x"84", x"84", x"84", x"83", x"82", x"80", 
        x"83", x"83", x"83", x"84", x"85", x"84", x"82", x"82", x"83", x"81", x"81", x"83", x"83", x"85", x"85", 
        x"83", x"83", x"82", x"82", x"82", x"82", x"86", x"87", x"84", x"83", x"84", x"83", x"83", x"82", x"80", 
        x"81", x"82", x"83", x"82", x"82", x"81", x"80", x"81", x"82", x"82", x"81", x"7f", x"7e", x"82", x"82", 
        x"81", x"81", x"81", x"82", x"82", x"81", x"80", x"80", x"81", x"83", x"83", x"81", x"82", x"81", x"81", 
        x"80", x"81", x"82", x"82", x"82", x"80", x"80", x"81", x"82", x"81", x"80", x"80", x"80", x"80", x"81", 
        x"81", x"81", x"81", x"81", x"80", x"80", x"81", x"81", x"81", x"80", x"7f", x"7f", x"7e", x"7e", x"7e", 
        x"7e", x"7d", x"7d", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"80", x"7e", x"7d", x"7d", x"7c", 
        x"7f", x"80", x"7c", x"7e", x"7f", x"81", x"81", x"7f", x"7e", x"7f", x"7d", x"7d", x"7e", x"7e", x"7e", 
        x"7f", x"7f", x"7d", x"7c", x"7d", x"80", x"80", x"7f", x"7f", x"7f", x"7f", x"7e", x"7f", x"80", x"80", 
        x"7f", x"7d", x"7d", x"7f", x"7f", x"7f", x"7e", x"7f", x"7e", x"7e", x"7f", x"7f", x"80", x"7f", x"7e", 
        x"7d", x"7d", x"7e", x"7c", x"7b", x"7d", x"7e", x"7c", x"7b", x"7e", x"80", x"7f", x"7d", x"7e", x"7f", 
        x"7d", x"7d", x"7f", x"7e", x"7c", x"7b", x"7c", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", 
        x"7c", x"7c", x"7d", x"7d", x"7d", x"7d", x"7d", x"7e", x"7c", x"7c", x"7d", x"7e", x"7d", x"7b", x"7b", 
        x"7e", x"7b", x"7d", x"7d", x"7c", x"7c", x"7b", x"7b", x"7b", x"7a", x"78", x"79", x"7b", x"7c", x"7c", 
        x"7b", x"7a", x"7a", x"7c", x"7a", x"78", x"78", x"7a", x"7b", x"7c", x"7a", x"78", x"78", x"78", x"79", 
        x"79", x"7a", x"7b", x"7a", x"79", x"76", x"75", x"77", x"77", x"79", x"7b", x"7b", x"78", x"77", x"77", 
        x"79", x"7d", x"7b", x"79", x"7a", x"7a", x"7c", x"7c", x"7b", x"79", x"78", x"7a", x"7c", x"7b", x"7b", 
        x"7b", x"7a", x"7a", x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7a", x"79", x"79", x"79", 
        x"79", x"7a", x"7c", x"7b", x"7a", x"7d", x"7c", x"7c", x"7d", x"7c", x"7b", x"7a", x"7b", x"7c", x"7c", 
        x"7b", x"7b", x"7a", x"7c", x"79", x"78", x"79", x"7a", x"7a", x"7a", x"7a", x"7b", x"7c", x"7c", x"7c", 
        x"7c", x"7c", x"7c", x"7a", x"79", x"7a", x"7a", x"7b", x"7b", x"7b", x"7a", x"79", x"7b", x"7d", x"7e", 
        x"7d", x"7c", x"7c", x"7d", x"7c", x"7c", x"7d", x"7e", x"7e", x"7e", x"7d", x"7d", x"7e", x"7f", x"7e", 
        x"7e", x"7d", x"7f", x"7e", x"7d", x"7e", x"7f", x"80", x"7e", x"7d", x"80", x"81", x"80", x"81", x"82", 
        x"81", x"7f", x"7f", x"7d", x"7e", x"81", x"7d", x"7d", x"81", x"85", x"86", x"79", x"5a", x"56", x"6e", 
        x"80", x"bd", x"dc", x"d1", x"d1", x"d3", x"d8", x"d7", x"cb", x"cf", x"ce", x"d0", x"d0", x"d0", x"cf", 
        x"cf", x"d0", x"d0", x"d0", x"cf", x"cf", x"d0", x"cf", x"cf", x"d0", x"d0", x"d1", x"d2", x"d2", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d0", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"d0", x"d1", x"d0", x"d1", 
        x"d3", x"d2", x"d0", x"d0", x"d0", x"d0", x"ce", x"d4", x"d2", x"be", x"cf", x"d6", x"d3", x"d5", x"d0", 
        x"dc", x"f0", x"ea", x"ed", x"ee", x"eb", x"ec", x"ed", x"ef", x"ef", x"ec", x"e4", x"db", x"cd", x"c2", 
        x"c6", x"d5", x"e5", x"ef", x"f4", x"ef", x"ac", x"65", x"5f", x"5e", x"5f", x"7e", x"e2", x"f9", x"f6", 
        x"c8", x"6a", x"5b", x"85", x"dd", x"f7", x"fa", x"f9", x"f9", x"f8", x"d7", x"7f", x"5b", x"5f", x"5b", 
        x"69", x"b0", x"f1", x"f6", x"f5", x"cb", x"91", x"68", x"5b", x"5e", x"70", x"b4", x"c3", x"80", x"5b", 
        x"5e", x"5c", x"7a", x"df", x"f2", x"ed", x"da", x"bd", x"9b", x"78", x"68", x"62", x"5d", x"5f", x"5e", 
        x"59", x"5f", x"61", x"5d", x"5a", x"5d", x"5e", x"5d", x"5f", x"5f", x"5f", x"5d", x"5c", x"5d", x"62", 
        x"93", x"e8", x"f0", x"ec", x"ed", x"ef", x"ef", x"ed", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f3", x"f2", x"ee", x"e7", x"d5", x"c2", x"b5", x"c3", x"d7", x"e5", x"ed", x"f0", x"f2", x"ef", 
        x"ee", x"ed", x"ec", x"ed", x"ee", x"ee", x"ef", x"f0", x"ee", x"ef", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ee", x"ef", x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f0", x"ee", x"ee", x"ec", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"f1", x"f2", x"ec", x"e9", x"ec", x"ec", x"ec", x"eb", x"ec", 
        x"ed", x"ec", x"eb", x"ee", x"ea", x"e1", x"db", x"de", x"e2", x"d9", x"b9", x"92", x"79", x"7c", x"82", 
        x"7f", x"80", x"83", x"83", x"82", x"85", x"86", x"83", x"83", x"85", x"85", x"84", x"84", x"85", x"84", 
        x"82", x"81", x"82", x"83", x"84", x"84", x"84", x"85", x"87", x"85", x"82", x"80", x"81", x"82", x"82", 
        x"82", x"81", x"81", x"82", x"82", x"82", x"81", x"83", x"83", x"83", x"83", x"83", x"82", x"82", x"83", 
        x"83", x"84", x"83", x"81", x"81", x"81", x"84", x"84", x"82", x"84", x"85", x"84", x"83", x"83", x"81", 
        x"81", x"82", x"84", x"83", x"82", x"81", x"83", x"83", x"82", x"83", x"83", x"83", x"81", x"80", x"81", 
        x"82", x"82", x"81", x"81", x"82", x"82", x"81", x"81", x"82", x"83", x"83", x"82", x"82", x"80", x"80", 
        x"7f", x"81", x"82", x"80", x"80", x"80", x"81", x"81", x"81", x"82", x"82", x"80", x"81", x"82", x"82", 
        x"82", x"82", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"7e", x"7f", x"7c", 
        x"7c", x"7d", x"7e", x"7c", x"7d", x"7f", x"7f", x"7f", x"7f", x"7d", x"7e", x"80", x"80", x"80", x"80", 
        x"80", x"7f", x"7e", x"7e", x"7f", x"81", x"7e", x"7d", x"80", x"80", x"7d", x"7f", x"7f", x"7e", x"7e", 
        x"7e", x"7f", x"7f", x"7c", x"7c", x"7f", x"80", x"7f", x"7f", x"7f", x"7e", x"7e", x"7e", x"7e", x"7e", 
        x"7e", x"7b", x"7b", x"80", x"80", x"7f", x"7f", x"7e", x"7d", x"7d", x"7f", x"7f", x"7f", x"7f", x"80", 
        x"80", x"7d", x"7e", x"7e", x"7f", x"80", x"7e", x"7c", x"7d", x"7d", x"7c", x"7d", x"7f", x"7e", x"7c", 
        x"7d", x"7d", x"80", x"7f", x"7f", x"7e", x"7d", x"7d", x"7e", x"80", x"7e", x"7c", x"7d", x"7e", x"7d", 
        x"7d", x"7d", x"7d", x"7e", x"7e", x"7f", x"7f", x"7f", x"7a", x"79", x"7a", x"7b", x"7b", x"7d", x"7d", 
        x"80", x"7e", x"7f", x"7f", x"7c", x"7d", x"7b", x"7a", x"7b", x"7a", x"7a", x"7a", x"7a", x"7b", x"7b", 
        x"7b", x"7a", x"7b", x"7d", x"7a", x"78", x"79", x"7d", x"7c", x"7a", x"7a", x"7a", x"79", x"77", x"78", 
        x"7a", x"7b", x"7b", x"7b", x"79", x"75", x"77", x"7a", x"79", x"79", x"79", x"78", x"76", x"77", x"7b", 
        x"7c", x"7d", x"7b", x"78", x"77", x"77", x"7a", x"7a", x"7a", x"7a", x"7a", x"7c", x"7e", x"7a", x"79", 
        x"78", x"79", x"7a", x"7b", x"7d", x"7b", x"7b", x"7b", x"7b", x"7b", x"7b", x"7a", x"79", x"79", x"79", 
        x"78", x"7a", x"7d", x"7d", x"7c", x"7f", x"7e", x"7e", x"7d", x"7d", x"7d", x"7c", x"7b", x"7b", x"7c", 
        x"7a", x"7a", x"79", x"7a", x"79", x"78", x"79", x"7a", x"7b", x"7a", x"79", x"7b", x"7c", x"7d", x"7d", 
        x"7d", x"7c", x"7b", x"7c", x"7c", x"7d", x"7d", x"7e", x"7e", x"7f", x"7c", x"79", x"7b", x"7d", x"7d", 
        x"7e", x"7e", x"7e", x"7d", x"7e", x"7e", x"7f", x"80", x"80", x"7f", x"7e", x"7e", x"7f", x"80", x"7f", 
        x"7e", x"7e", x"7d", x"7c", x"7c", x"7d", x"7f", x"80", x"7f", x"81", x"83", x"81", x"80", x"81", x"83", 
        x"81", x"80", x"7f", x"7f", x"81", x"7d", x"7a", x"81", x"85", x"7f", x"68", x"57", x"65", x"85", x"8a", 
        x"78", x"ba", x"d9", x"d0", x"d2", x"d4", x"da", x"d9", x"cd", x"d0", x"cf", x"d0", x"d0", x"cf", x"ce", 
        x"cf", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"ce", x"d0", x"d2", x"d1", x"d2", x"d3", x"d2", x"d0", 
        x"d1", x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"d0", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"d0", 
        x"d3", x"d2", x"d0", x"d0", x"d1", x"cf", x"cc", x"d3", x"dc", x"d0", x"d5", x"d1", x"d0", x"d5", x"d0", 
        x"dc", x"f0", x"eb", x"ed", x"ee", x"ec", x"ec", x"eb", x"ec", x"ee", x"f0", x"ef", x"ef", x"ef", x"eb", 
        x"de", x"cd", x"bf", x"c2", x"ce", x"d9", x"a1", x"60", x"5c", x"60", x"5f", x"7f", x"e1", x"f9", x"f6", 
        x"c9", x"6f", x"5a", x"63", x"b5", x"f1", x"fb", x"fb", x"f9", x"fa", x"d9", x"82", x"5c", x"59", x"5c", 
        x"60", x"84", x"d6", x"f5", x"f9", x"f5", x"e0", x"b6", x"7e", x"66", x"5e", x"71", x"93", x"78", x"5a", 
        x"5d", x"61", x"77", x"de", x"f8", x"fb", x"f8", x"f4", x"eb", x"d9", x"bf", x"9b", x"75", x"62", x"5c", 
        x"5e", x"5d", x"5f", x"5e", x"5c", x"60", x"5d", x"5a", x"5f", x"5e", x"5e", x"5f", x"5d", x"5d", x"62", 
        x"8f", x"e6", x"f0", x"ec", x"ed", x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"f0", x"f1", x"ee", x"ee", x"f4", x"f3", x"ec", x"e4", x"cc", x"b7", x"b6", x"c9", x"da", x"e4", x"ec", 
        x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"f0", x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"f2", x"f0", 
        x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ec", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"ee", x"ea", x"eb", x"ed", x"ee", x"ef", x"ee", 
        x"ec", x"eb", x"ec", x"ef", x"f3", x"f3", x"ee", x"e6", x"e0", x"dc", x"e3", x"dd", x"c3", x"9c", x"84", 
        x"78", x"7c", x"80", x"83", x"87", x"86", x"83", x"84", x"84", x"81", x"82", x"83", x"81", x"7e", x"81", 
        x"84", x"84", x"84", x"84", x"85", x"85", x"85", x"85", x"84", x"83", x"82", x"82", x"83", x"83", x"84", 
        x"82", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"84", x"83", x"82", x"82", x"81", 
        x"81", x"82", x"82", x"81", x"80", x"81", x"81", x"82", x"83", x"83", x"84", x"85", x"84", x"83", x"80", 
        x"80", x"80", x"82", x"83", x"82", x"81", x"82", x"83", x"81", x"83", x"82", x"83", x"82", x"7f", x"81", 
        x"82", x"83", x"82", x"82", x"83", x"82", x"80", x"80", x"81", x"82", x"83", x"82", x"82", x"82", x"82", 
        x"82", x"82", x"83", x"82", x"82", x"80", x"82", x"81", x"81", x"82", x"82", x"80", x"80", x"81", x"81", 
        x"81", x"81", x"7f", x"7f", x"80", x"80", x"80", x"80", x"80", x"80", x"81", x"80", x"7e", x"7f", x"7c", 
        x"7c", x"7d", x"7f", x"7d", x"7d", x"80", x"7f", x"7f", x"7f", x"7d", x"7e", x"81", x"80", x"7f", x"7f", 
        x"7f", x"80", x"80", x"7f", x"7f", x"81", x"7e", x"7e", x"80", x"80", x"7e", x"7e", x"7f", x"7e", x"7e", 
        x"7e", x"7f", x"80", x"80", x"7f", x"7f", x"7f", x"80", x"7d", x"80", x"7f", x"7d", x"7b", x"7b", x"7c", 
        x"7e", x"7e", x"7e", x"81", x"80", x"80", x"80", x"7e", x"7d", x"7e", x"7d", x"7d", x"7e", x"7f", x"7f", 
        x"7f", x"7e", x"7e", x"7e", x"7f", x"7f", x"7e", x"7d", x"7f", x"7d", x"7c", x"7d", x"7e", x"7d", x"7c", 
        x"7e", x"7e", x"80", x"7f", x"7f", x"7f", x"7e", x"7d", x"7f", x"81", x"7f", x"7e", x"7e", x"7e", x"7e", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"7e", x"7d", x"7d", x"7b", x"7a", x"7b", x"7c", x"7e", x"7d", x"7e", 
        x"7f", x"7e", x"7f", x"7f", x"7c", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7a", x"79", x"7b", x"7b", 
        x"7c", x"7a", x"7b", x"7d", x"7b", x"79", x"7a", x"7c", x"7b", x"7a", x"7a", x"7a", x"79", x"78", x"78", 
        x"79", x"79", x"7b", x"7b", x"7a", x"77", x"78", x"7a", x"79", x"79", x"78", x"77", x"77", x"78", x"7a", 
        x"7c", x"7b", x"7c", x"7a", x"78", x"79", x"7a", x"7b", x"7a", x"79", x"79", x"7a", x"7c", x"7c", x"7b", 
        x"79", x"77", x"77", x"78", x"78", x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7a", x"7b", x"7c", x"7b", 
        x"79", x"7a", x"7c", x"7d", x"7b", x"7d", x"7d", x"7d", x"7c", x"7b", x"7c", x"7c", x"7b", x"7b", x"7c", 
        x"7a", x"7a", x"79", x"7a", x"7a", x"7a", x"79", x"7b", x"7c", x"7c", x"7a", x"7c", x"7c", x"7d", x"7d", 
        x"7c", x"7c", x"7b", x"7d", x"7f", x"7f", x"7d", x"7c", x"7c", x"7c", x"7c", x"7b", x"7c", x"7d", x"7e", 
        x"7f", x"80", x"7e", x"7a", x"7c", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", 
        x"7e", x"7e", x"7d", x"7c", x"7d", x"7d", x"7e", x"7f", x"7e", x"7f", x"7f", x"7d", x"7d", x"7f", x"81", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"87", x"82", x"70", x"5a", x"5e", x"7c", x"8a", x"86", x"85", 
        x"7b", x"b9", x"d9", x"d0", x"d1", x"d3", x"d8", x"d8", x"cf", x"d2", x"ce", x"cf", x"d0", x"ce", x"cd", 
        x"ce", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"ce", x"d1", x"d3", x"d3", x"d3", x"d3", x"d1", x"cf", 
        x"d1", x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"cf", x"cf", x"ce", x"ce", x"ce", x"cf", x"cf", x"d0", 
        x"d3", x"d2", x"d0", x"d0", x"d1", x"d0", x"d0", x"d2", x"da", x"ce", x"d2", x"d3", x"d1", x"d4", x"d2", 
        x"dd", x"f0", x"ec", x"ee", x"ef", x"ed", x"ed", x"ec", x"eb", x"eb", x"ed", x"f0", x"f0", x"ef", x"ed", 
        x"ef", x"f1", x"e9", x"d7", x"c8", x"ba", x"9c", x"6e", x"60", x"5a", x"59", x"7b", x"e1", x"fb", x"f6", 
        x"c8", x"70", x"5e", x"5b", x"84", x"db", x"f6", x"f8", x"fb", x"fa", x"d9", x"86", x"5a", x"59", x"5e", 
        x"5c", x"64", x"9b", x"dc", x"f9", x"f8", x"f6", x"f5", x"d3", x"a6", x"76", x"5b", x"61", x"63", x"5f", 
        x"5d", x"5d", x"75", x"da", x"f7", x"f9", x"f2", x"f1", x"f6", x"f6", x"f6", x"f0", x"d5", x"94", x"62", 
        x"5d", x"59", x"5b", x"5d", x"5e", x"60", x"5b", x"5d", x"60", x"5d", x"5e", x"60", x"5e", x"5d", x"61", 
        x"86", x"df", x"ef", x"ed", x"ee", x"f0", x"ef", x"ee", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ee", x"f0", x"ee", x"ed", x"ef", x"f2", x"f2", x"ee", x"f2", x"ec", x"db", x"c3", x"b9", x"b8", x"cb", 
        x"db", x"e9", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"f1", x"f0", x"ee", x"ed", x"f0", x"f1", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ec", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f0", x"ed", x"eb", x"e9", x"e8", x"e7", x"e8", 
        x"ea", x"ec", x"f1", x"ef", x"ee", x"ef", x"f2", x"f2", x"ee", x"e6", x"dc", x"d5", x"d9", x"e1", x"d0", 
        x"ac", x"8d", x"7e", x"75", x"79", x"82", x"86", x"86", x"82", x"80", x"83", x"84", x"82", x"80", x"82", 
        x"85", x"85", x"85", x"85", x"86", x"85", x"85", x"84", x"81", x"83", x"84", x"85", x"85", x"85", x"84", 
        x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"83", x"82", x"83", x"84", x"84", x"83", x"83", x"82", 
        x"82", x"83", x"83", x"83", x"83", x"84", x"81", x"81", x"84", x"84", x"84", x"85", x"85", x"83", x"83", 
        x"82", x"83", x"83", x"83", x"82", x"81", x"81", x"83", x"82", x"83", x"81", x"82", x"82", x"80", x"81", 
        x"83", x"83", x"84", x"84", x"84", x"82", x"7f", x"7f", x"80", x"82", x"83", x"82", x"82", x"82", x"84", 
        x"83", x"82", x"83", x"82", x"83", x"81", x"82", x"81", x"81", x"82", x"81", x"80", x"80", x"80", x"81", 
        x"80", x"80", x"7f", x"7f", x"81", x"81", x"80", x"80", x"80", x"81", x"81", x"81", x"7f", x"80", x"7e", 
        x"7e", x"7f", x"80", x"7f", x"7f", x"80", x"7f", x"7f", x"80", x"7f", x"80", x"81", x"7f", x"7e", x"7e", 
        x"7f", x"7f", x"80", x"7f", x"80", x"82", x"80", x"7f", x"81", x"80", x"7f", x"7f", x"7f", x"7f", x"7f", 
        x"7f", x"7f", x"7f", x"81", x"80", x"7e", x"80", x"82", x"7f", x"80", x"81", x"7f", x"7d", x"7d", x"7d", 
        x"7e", x"7f", x"81", x"81", x"7f", x"80", x"80", x"7e", x"7e", x"80", x"7e", x"7d", x"7e", x"7f", x"7d", 
        x"7b", x"7d", x"7e", x"7e", x"7e", x"7d", x"7e", x"7e", x"7f", x"7d", x"7c", x"7e", x"7e", x"7d", x"7c", 
        x"7e", x"7e", x"80", x"7f", x"7f", x"7f", x"7e", x"7e", x"80", x"80", x"7e", x"7d", x"7e", x"7e", x"7e", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7e", x"7e", x"7e", x"7c", x"7c", x"7d", x"7e", x"7b", x"7c", 
        x"7e", x"7d", x"7e", x"80", x"7d", x"7e", x"7f", x"7e", x"7f", x"7f", x"7e", x"7d", x"7c", x"7d", x"7c", 
        x"7c", x"7b", x"7b", x"7d", x"7b", x"7a", x"7b", x"79", x"7a", x"7b", x"7b", x"79", x"78", x"7b", x"78", 
        x"77", x"78", x"79", x"7b", x"7b", x"7a", x"79", x"7a", x"79", x"79", x"78", x"79", x"7c", x"7c", x"7b", 
        x"7d", x"7a", x"7c", x"7a", x"77", x"79", x"7a", x"7b", x"7a", x"79", x"79", x"79", x"7b", x"7b", x"7b", 
        x"7a", x"7a", x"7b", x"7c", x"7d", x"7b", x"7b", x"7b", x"7c", x"7c", x"7b", x"7a", x"7b", x"7b", x"7b", 
        x"7a", x"7c", x"7d", x"7d", x"7a", x"7a", x"7b", x"7b", x"7a", x"79", x"79", x"7b", x"7c", x"7c", x"7c", 
        x"7b", x"7d", x"7b", x"7c", x"7c", x"7b", x"7a", x"7b", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", x"7d", 
        x"7d", x"7d", x"7c", x"7d", x"7c", x"7c", x"7d", x"7d", x"7e", x"7f", x"7e", x"7d", x"7d", x"7e", x"7e", 
        x"7f", x"7f", x"7c", x"7b", x"7e", x"80", x"80", x"7e", x"7d", x"7e", x"7e", x"7f", x"7f", x"7f", x"7f", 
        x"7f", x"7f", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7e", x"7f", x"7e", x"7f", x"80", x"81", 
        x"7f", x"80", x"7e", x"7d", x"82", x"84", x"7b", x"62", x"5a", x"71", x"8b", x"8e", x"87", x"88", x"84", 
        x"78", x"ba", x"db", x"d1", x"d1", x"d2", x"d6", x"d7", x"cf", x"d2", x"ce", x"cf", x"d0", x"cf", x"ce", 
        x"ce", x"ce", x"cf", x"d0", x"cf", x"cf", x"ce", x"ce", x"d1", x"d4", x"d4", x"d4", x"d3", x"d0", x"cf", 
        x"d1", x"d2", x"d1", x"d1", x"d0", x"d0", x"cf", x"cf", x"ce", x"ce", x"ce", x"ce", x"cf", x"cf", x"d0", 
        x"d3", x"d2", x"d0", x"d0", x"d1", x"d0", x"cf", x"d0", x"dc", x"cf", x"d0", x"d3", x"d2", x"d4", x"d3", 
        x"dc", x"ef", x"ec", x"ee", x"ee", x"ec", x"ed", x"ed", x"ed", x"ec", x"ed", x"ef", x"f0", x"ee", x"ee", 
        x"ed", x"ec", x"ed", x"ef", x"ef", x"e8", x"d7", x"ba", x"a0", x"85", x"6f", x"77", x"d2", x"f0", x"f7", 
        x"cf", x"72", x"5c", x"5d", x"69", x"b4", x"ef", x"f6", x"fa", x"f8", x"dd", x"89", x"5e", x"5e", x"5e", 
        x"5e", x"5c", x"67", x"9e", x"d9", x"f1", x"f7", x"fa", x"f4", x"e9", x"bc", x"7f", x"62", x"5c", x"60", 
        x"5f", x"60", x"74", x"d5", x"f5", x"f7", x"de", x"c2", x"c8", x"e1", x"ef", x"f6", x"eb", x"a7", x"64", 
        x"5b", x"59", x"5c", x"5c", x"5f", x"61", x"5c", x"5c", x"5f", x"5d", x"5e", x"60", x"5e", x"5c", x"5f", 
        x"7f", x"dc", x"ef", x"ee", x"ef", x"f0", x"ef", x"ee", x"ef", x"ed", x"ee", x"ef", x"f0", x"f0", x"ef", 
        x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f2", x"f0", x"ee", x"f0", x"f0", x"e6", x"d8", x"c3", 
        x"bf", x"c3", x"cf", x"de", x"ea", x"f2", x"f3", x"f0", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ec", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"ee", x"eb", x"ea", x"ec", 
        x"ee", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"e9", x"dc", x"d5", x"d9", 
        x"de", x"cf", x"b5", x"95", x"7f", x"7b", x"7f", x"84", x"84", x"84", x"86", x"84", x"82", x"83", x"82", 
        x"82", x"85", x"85", x"85", x"85", x"85", x"85", x"84", x"82", x"84", x"85", x"86", x"85", x"85", x"84", 
        x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"82", x"83", x"84", x"85", x"85", x"85", x"84", x"83", 
        x"82", x"82", x"82", x"82", x"82", x"82", x"81", x"82", x"85", x"85", x"84", x"83", x"83", x"83", x"81", 
        x"80", x"80", x"82", x"83", x"83", x"82", x"82", x"84", x"83", x"82", x"80", x"82", x"82", x"81", x"81", 
        x"83", x"84", x"85", x"85", x"84", x"83", x"82", x"81", x"81", x"83", x"83", x"82", x"81", x"80", x"83", 
        x"82", x"81", x"81", x"80", x"83", x"81", x"82", x"82", x"82", x"81", x"80", x"80", x"80", x"81", x"81", 
        x"81", x"80", x"80", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"80", x"81", x"81", x"80", 
        x"7f", x"80", x"81", x"81", x"80", x"7f", x"7f", x"7f", x"7f", x"80", x"81", x"81", x"81", x"80", x"80", 
        x"80", x"80", x"80", x"80", x"81", x"81", x"81", x"81", x"80", x"80", x"80", x"7f", x"7f", x"80", x"81", 
        x"80", x"7f", x"81", x"81", x"80", x"80", x"80", x"80", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
        x"7e", x"80", x"81", x"7f", x"7e", x"7f", x"7f", x"7e", x"7f", x"81", x"80", x"80", x"7f", x"7e", x"7d", 
        x"7c", x"7d", x"7e", x"7e", x"7d", x"7d", x"7d", x"7f", x"7d", x"7c", x"7c", x"7e", x"7f", x"7f", x"7d", 
        x"7e", x"7e", x"80", x"7f", x"7f", x"7f", x"7e", x"80", x"7f", x"7e", x"7d", x"7d", x"7d", x"7e", x"7e", 
        x"7d", x"7d", x"7e", x"7f", x"80", x"80", x"7f", x"7e", x"7d", x"7c", x"7d", x"7c", x"7d", x"7d", x"7b", 
        x"7e", x"7d", x"7e", x"80", x"7e", x"7f", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", 
        x"7b", x"7a", x"7a", x"7c", x"7b", x"7a", x"7c", x"7a", x"79", x"7a", x"7b", x"7b", x"7b", x"7c", x"7a", 
        x"78", x"78", x"79", x"7b", x"7a", x"79", x"79", x"7a", x"7a", x"7a", x"79", x"7b", x"7d", x"7d", x"7a", 
        x"7a", x"78", x"7c", x"7c", x"7a", x"7b", x"7a", x"7b", x"7b", x"79", x"79", x"79", x"7b", x"79", x"79", 
        x"79", x"7a", x"7b", x"7b", x"7b", x"7b", x"7c", x"7c", x"7d", x"7d", x"7c", x"7b", x"79", x"7a", x"7b", 
        x"7b", x"7d", x"7f", x"7d", x"7b", x"7a", x"7b", x"7b", x"7b", x"7a", x"7b", x"7c", x"7c", x"7b", x"7c", 
        x"7c", x"7f", x"7d", x"7e", x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7d", x"7e", 
        x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7e", x"7e", x"7f", x"7f", x"7e", x"7e", x"7f", x"80", x"7f", 
        x"7e", x"7d", x"7c", x"7e", x"80", x"81", x"81", x"7f", x"7e", x"7f", x"7f", x"7e", x"7e", x"7e", x"7e", 
        x"7e", x"7f", x"7d", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"81", x"81", x"80", x"82", x"82", x"80", 
        x"7f", x"7d", x"7f", x"85", x"83", x"79", x"6e", x"69", x"7e", x"90", x"88", x"89", x"87", x"83", x"81", 
        x"79", x"b9", x"da", x"d2", x"d1", x"d2", x"d6", x"d8", x"cd", x"d1", x"ce", x"d0", x"d0", x"d0", x"d0", 
        x"cd", x"ce", x"cf", x"d0", x"cf", x"ce", x"cd", x"cd", x"d1", x"d3", x"d3", x"d3", x"d3", x"d1", x"cf", 
        x"d1", x"d2", x"d1", x"d1", x"d0", x"d0", x"cf", x"cf", x"ce", x"ce", x"ce", x"ce", x"cf", x"cf", x"d0", 
        x"d3", x"d2", x"d0", x"d0", x"d1", x"cf", x"cb", x"cf", x"df", x"d2", x"d0", x"d3", x"d3", x"d4", x"d3", 
        x"dc", x"ef", x"ed", x"ee", x"ee", x"ed", x"ed", x"ef", x"ef", x"ed", x"ed", x"ed", x"f0", x"f0", x"ee", 
        x"ec", x"ec", x"ed", x"ec", x"ed", x"ef", x"ec", x"f1", x"eb", x"db", x"bf", x"a9", x"b9", x"c8", x"d5", 
        x"bd", x"6e", x"59", x"5f", x"61", x"84", x"de", x"f8", x"f8", x"f9", x"e0", x"89", x"5d", x"5b", x"5d", 
        x"5e", x"65", x"5d", x"66", x"8d", x"c6", x"ec", x"fb", x"f6", x"f9", x"f0", x"c5", x"81", x"5b", x"60", 
        x"5f", x"63", x"6f", x"d5", x"f6", x"f6", x"ca", x"82", x"72", x"93", x"af", x"cd", x"df", x"a6", x"63", 
        x"59", x"5d", x"5f", x"5e", x"5e", x"5c", x"62", x"68", x"5f", x"58", x"5c", x"60", x"62", x"60", x"5e", 
        x"7b", x"db", x"ef", x"ee", x"ef", x"ef", x"ee", x"ed", x"ef", x"ed", x"ee", x"ef", x"ef", x"f0", x"ef", 
        x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", 
        x"f2", x"f0", x"ef", x"ef", x"ee", x"ed", x"ec", x"ef", x"f2", x"f1", x"ef", x"ed", x"f1", x"f5", x"ef", 
        x"e3", x"cf", x"be", x"bb", x"c5", x"d1", x"e6", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f0", x"ef", x"ee", x"ea", x"ee", x"ef", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f2", x"f1", x"ea", x"e0", 
        x"d9", x"d8", x"df", x"dc", x"bd", x"9b", x"85", x"78", x"7c", x"82", x"86", x"86", x"85", x"85", x"84", 
        x"84", x"84", x"84", x"84", x"84", x"85", x"84", x"85", x"85", x"84", x"84", x"85", x"84", x"84", x"84", 
        x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"83", x"84", x"84", x"85", x"85", x"84", x"85", 
        x"85", x"84", x"83", x"83", x"83", x"82", x"83", x"84", x"84", x"85", x"84", x"81", x"82", x"84", x"85", 
        x"83", x"82", x"83", x"84", x"83", x"82", x"81", x"83", x"82", x"83", x"82", x"83", x"84", x"82", x"82", 
        x"83", x"84", x"85", x"85", x"84", x"85", x"85", x"83", x"83", x"84", x"83", x"81", x"81", x"80", x"82", 
        x"82", x"81", x"81", x"81", x"83", x"82", x"82", x"82", x"82", x"80", x"80", x"80", x"81", x"81", x"81", 
        x"81", x"81", x"82", x"82", x"82", x"81", x"81", x"81", x"81", x"81", x"81", x"80", x"81", x"80", x"81", 
        x"7f", x"80", x"82", x"81", x"80", x"7f", x"7f", x"7f", x"7f", x"80", x"81", x"82", x"82", x"82", x"83", 
        x"82", x"80", x"80", x"81", x"81", x"80", x"82", x"81", x"80", x"80", x"81", x"80", x"7f", x"80", x"81", 
        x"80", x"80", x"82", x"81", x"81", x"82", x"7f", x"7e", x"7f", x"81", x"82", x"81", x"80", x"7f", x"7e", 
        x"7d", x"7f", x"7f", x"7d", x"7e", x"7f", x"7f", x"7f", x"7f", x"7f", x"80", x"81", x"80", x"7f", x"80", 
        x"81", x"7e", x"7f", x"7e", x"7d", x"7d", x"7e", x"7f", x"7d", x"7c", x"7c", x"7e", x"7f", x"80", x"7f", 
        x"7f", x"7e", x"80", x"7f", x"7f", x"7f", x"7e", x"7f", x"7f", x"7e", x"7f", x"7f", x"7e", x"7d", x"7d", 
        x"7d", x"7d", x"7d", x"7e", x"7e", x"7e", x"7e", x"7e", x"7b", x"7c", x"7d", x"7b", x"7e", x"80", x"7d", 
        x"7f", x"7d", x"7e", x"7e", x"7c", x"7c", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", 
        x"7b", x"79", x"79", x"7b", x"7a", x"7a", x"7c", x"7c", x"7a", x"79", x"7b", x"7c", x"7d", x"7b", x"7b", 
        x"7b", x"79", x"7a", x"7a", x"79", x"77", x"78", x"7b", x"79", x"79", x"79", x"7a", x"7b", x"7c", x"7b", 
        x"7a", x"7a", x"7b", x"7b", x"7b", x"7a", x"7c", x"7c", x"7c", x"7a", x"79", x"79", x"7a", x"79", x"7a", 
        x"7a", x"7a", x"7b", x"7b", x"7b", x"7b", x"7b", x"7c", x"7d", x"7d", x"7c", x"7b", x"7b", x"7b", x"7c", 
        x"7b", x"7c", x"7e", x"7c", x"7b", x"7b", x"7b", x"7c", x"7d", x"7d", x"7d", x"7d", x"7c", x"7b", x"7c", 
        x"7c", x"7f", x"7d", x"7e", x"7e", x"7f", x"7e", x"7d", x"7c", x"7c", x"7e", x"7e", x"7e", x"7e", x"7e", 
        x"7d", x"7c", x"7c", x"7b", x"7b", x"7c", x"7d", x"7d", x"7e", x"7f", x"7f", x"7f", x"7f", x"7f", x"7e", 
        x"7e", x"7d", x"7c", x"7d", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"7e", x"7e", x"7e", x"7e", 
        x"7e", x"7f", x"7d", x"7d", x"7f", x"7f", x"7f", x"7f", x"81", x"81", x"80", x"80", x"80", x"7f", x"7e", 
        x"81", x"84", x"89", x"7a", x"6d", x"84", x"b1", x"9d", x"8a", x"8c", x"88", x"84", x"85", x"87", x"81", 
        x"79", x"b8", x"da", x"d1", x"d0", x"d2", x"d8", x"da", x"cc", x"d1", x"d0", x"d0", x"d0", x"cf", x"d0", 
        x"cd", x"ce", x"cf", x"d0", x"cf", x"ce", x"cd", x"cd", x"d0", x"d2", x"d1", x"d2", x"d3", x"d1", x"d0", 
        x"d1", x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", 
        x"d3", x"d2", x"d0", x"d0", x"d1", x"d0", x"d1", x"d1", x"db", x"cf", x"d3", x"d5", x"d3", x"d4", x"d4", 
        x"dc", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ed", x"ec", x"ec", x"ef", x"ef", x"eb", 
        x"ec", x"ee", x"ee", x"ed", x"ed", x"ec", x"e8", x"ee", x"ee", x"ef", x"ee", x"e7", x"dd", x"d5", x"cb", 
        x"b1", x"7d", x"64", x"5c", x"5e", x"61", x"b0", x"f5", x"fa", x"fa", x"df", x"89", x"57", x"5b", x"5c", 
        x"6d", x"a3", x"84", x"61", x"63", x"6f", x"98", x"c9", x"ee", x"f9", x"f6", x"ee", x"c1", x"79", x"5e", 
        x"61", x"5f", x"6c", x"cc", x"f3", x"f8", x"d3", x"83", x"59", x"57", x"60", x"71", x"89", x"7d", x"5f", 
        x"5a", x"5e", x"5d", x"5c", x"5b", x"5b", x"88", x"b7", x"a3", x"85", x"6e", x"5f", x"5d", x"61", x"5e", 
        x"7a", x"d9", x"ee", x"ee", x"ef", x"ef", x"ed", x"ed", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"ef", x"eb", x"df", x"d0", x"c1", x"b6", x"bf", x"d6", x"ec", x"f4", x"f3", x"ef", x"ee", x"ef", 
        x"ee", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"ea", x"ee", x"ef", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f3", x"f1", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f5", x"f3", x"f1", x"ef", x"ee", x"f1", x"f3", x"f2", x"f1", x"ef", x"ef", x"f2", x"f3", 
        x"ee", x"e6", x"dd", x"d4", x"d4", x"d9", x"ce", x"b0", x"89", x"74", x"74", x"7c", x"84", x"84", x"81", 
        x"83", x"85", x"85", x"85", x"84", x"84", x"84", x"84", x"85", x"84", x"84", x"84", x"84", x"84", x"84", 
        x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"85", x"84", x"84", x"83", x"84", 
        x"84", x"83", x"83", x"83", x"83", x"81", x"83", x"86", x"84", x"84", x"83", x"82", x"82", x"84", x"84", 
        x"83", x"82", x"83", x"84", x"85", x"84", x"83", x"83", x"82", x"84", x"83", x"84", x"84", x"84", x"84", 
        x"83", x"84", x"85", x"84", x"83", x"84", x"85", x"83", x"83", x"84", x"83", x"81", x"82", x"82", x"83", 
        x"83", x"82", x"84", x"82", x"84", x"82", x"81", x"82", x"82", x"80", x"7f", x"80", x"81", x"81", x"80", 
        x"80", x"81", x"82", x"82", x"81", x"81", x"80", x"80", x"80", x"81", x"81", x"7f", x"81", x"80", x"81", 
        x"80", x"80", x"82", x"82", x"81", x"80", x"81", x"81", x"80", x"80", x"82", x"82", x"82", x"82", x"82", 
        x"82", x"80", x"80", x"81", x"81", x"7f", x"81", x"81", x"7f", x"80", x"80", x"80", x"80", x"80", x"80", 
        x"80", x"80", x"7f", x"7f", x"80", x"81", x"80", x"7f", x"82", x"80", x"7e", x"7e", x"7e", x"7f", x"81", 
        x"82", x"81", x"7e", x"7e", x"80", x"80", x"7f", x"7f", x"80", x"7d", x"7f", x"80", x"80", x"80", x"82", 
        x"82", x"80", x"7f", x"7e", x"7e", x"7f", x"7f", x"7f", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"7f", 
        x"7e", x"7e", x"80", x"7f", x"7f", x"7f", x"7e", x"7f", x"7e", x"7e", x"80", x"81", x"7e", x"7c", x"7d", 
        x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7e", x"7f", x"7e", x"7d", x"7c", x"7a", x"7c", x"7f", x"7e", 
        x"7f", x"7c", x"7c", x"7c", x"7a", x"7a", x"80", x"80", x"7e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7e", 
        x"7a", x"78", x"79", x"7a", x"7a", x"7a", x"7d", x"7d", x"7c", x"7d", x"7c", x"7b", x"7a", x"7a", x"7b", 
        x"7a", x"79", x"79", x"7a", x"79", x"77", x"78", x"79", x"77", x"78", x"79", x"7b", x"7b", x"7b", x"7c", 
        x"7a", x"7b", x"79", x"7a", x"7b", x"78", x"79", x"7b", x"7c", x"7b", x"7a", x"7a", x"7c", x"7b", x"7b", 
        x"7b", x"7b", x"7c", x"7e", x"7e", x"7c", x"7c", x"7d", x"7e", x"7d", x"7c", x"7b", x"7b", x"7b", x"7b", 
        x"7a", x"7b", x"7d", x"7c", x"7b", x"7b", x"7a", x"7b", x"7c", x"7c", x"7c", x"7c", x"7d", x"7b", x"7b", 
        x"7b", x"7d", x"7c", x"7c", x"7e", x"80", x"80", x"7d", x"7b", x"7c", x"7f", x"80", x"80", x"7f", x"7e", 
        x"7d", x"7b", x"7a", x"7c", x"7e", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7e", x"7e", x"7e", 
        x"7e", x"7f", x"7f", x"7e", x"7d", x"7e", x"7f", x"80", x"80", x"7f", x"7f", x"7e", x"7e", x"7e", x"7d", 
        x"7e", x"7f", x"7f", x"7f", x"80", x"80", x"7f", x"7f", x"80", x"80", x"7f", x"7f", x"80", x"80", x"82", 
        x"86", x"86", x"76", x"72", x"9a", x"c7", x"d1", x"9f", x"86", x"8b", x"88", x"87", x"88", x"88", x"86", 
        x"7e", x"ba", x"db", x"d2", x"d0", x"d1", x"d6", x"d9", x"cc", x"d2", x"d2", x"d1", x"cf", x"cf", x"d0", 
        x"ce", x"cd", x"cf", x"cf", x"cf", x"ce", x"cd", x"cd", x"cf", x"d0", x"d0", x"d1", x"d3", x"d2", x"d1", 
        x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"cf", x"cf", x"cf", x"d0", x"d0", x"d0", 
        x"d3", x"d2", x"d0", x"cf", x"d0", x"d0", x"d1", x"d3", x"de", x"d1", x"d4", x"d4", x"d2", x"d4", x"d4", 
        x"dc", x"ee", x"ee", x"ee", x"ed", x"ee", x"ed", x"ee", x"ee", x"ed", x"ed", x"ed", x"ee", x"ef", x"eb", 
        x"ec", x"ed", x"eb", x"ec", x"ee", x"ec", x"ed", x"ef", x"ed", x"ed", x"eb", x"ec", x"f0", x"f1", x"ea", 
        x"df", x"c9", x"ae", x"90", x"73", x"64", x"83", x"df", x"f3", x"f6", x"e3", x"8d", x"59", x"5d", x"5e", 
        x"6f", x"ca", x"c6", x"84", x"5e", x"5a", x"63", x"79", x"b1", x"e3", x"f5", x"f7", x"e8", x"9f", x"5e", 
        x"5f", x"5c", x"6b", x"c8", x"f3", x"f6", x"eb", x"c3", x"a1", x"7e", x"68", x"5c", x"5d", x"62", x"5e", 
        x"5c", x"5d", x"5d", x"5d", x"5d", x"65", x"ac", x"ef", x"e8", x"d8", x"b4", x"7c", x"5d", x"5e", x"5f", 
        x"7d", x"d8", x"ee", x"ed", x"ee", x"ee", x"ed", x"ed", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"ee", x"ef", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"ef", x"ed", x"f0", 
        x"ef", x"ee", x"f0", x"f2", x"ef", x"e7", x"d7", x"c8", x"bd", x"bf", x"ce", x"df", x"ec", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"eb", x"ef", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f0", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f1", x"ee", x"e6", x"dc", x"d8", x"d9", x"dd", x"d0", x"b3", x"91", x"79", x"76", x"7e", x"84", 
        x"86", x"88", x"86", x"86", x"86", x"84", x"84", x"84", x"84", x"84", x"84", x"85", x"84", x"84", x"84", 
        x"86", x"85", x"85", x"86", x"86", x"86", x"85", x"85", x"85", x"85", x"85", x"84", x"84", x"83", x"84", 
        x"83", x"82", x"82", x"84", x"84", x"83", x"84", x"85", x"83", x"81", x"81", x"84", x"84", x"84", x"86", 
        x"84", x"83", x"84", x"84", x"85", x"85", x"87", x"86", x"84", x"84", x"83", x"82", x"81", x"84", x"84", 
        x"83", x"83", x"84", x"83", x"81", x"83", x"83", x"82", x"82", x"83", x"83", x"81", x"82", x"82", x"83", 
        x"82", x"83", x"84", x"83", x"84", x"83", x"81", x"82", x"83", x"80", x"7f", x"80", x"80", x"80", x"7f", 
        x"7f", x"80", x"81", x"82", x"81", x"80", x"7f", x"80", x"80", x"80", x"80", x"7f", x"81", x"7f", x"81", 
        x"80", x"80", x"81", x"81", x"80", x"7f", x"83", x"82", x"80", x"81", x"82", x"82", x"81", x"81", x"81", 
        x"81", x"80", x"80", x"81", x"80", x"7e", x"80", x"81", x"7f", x"81", x"80", x"81", x"81", x"81", x"80", 
        x"80", x"80", x"7e", x"80", x"81", x"7f", x"7f", x"80", x"82", x"7f", x"7d", x"7e", x"80", x"80", x"81", 
        x"81", x"81", x"7f", x"80", x"82", x"82", x"7f", x"80", x"81", x"80", x"7f", x"7f", x"80", x"80", x"7f", 
        x"7f", x"80", x"7f", x"7e", x"7f", x"80", x"80", x"80", x"7f", x"7f", x"7f", x"7e", x"7e", x"7d", x"7e", 
        x"7e", x"7e", x"80", x"7f", x"7f", x"7f", x"7e", x"81", x"7f", x"7d", x"7e", x"7e", x"7d", x"7d", x"7e", 
        x"7e", x"7e", x"7e", x"7f", x"7f", x"80", x"7f", x"7e", x"7e", x"7c", x"7b", x"7b", x"7e", x"7e", x"7c", 
        x"7c", x"7b", x"7c", x"7d", x"7c", x"7d", x"7f", x"80", x"7f", x"7e", x"7e", x"7f", x"7f", x"7f", x"7e", 
        x"7b", x"7b", x"7c", x"7c", x"7b", x"7b", x"7e", x"7d", x"7c", x"7b", x"7b", x"7a", x"79", x"7a", x"7a", 
        x"79", x"7a", x"7b", x"7c", x"7b", x"78", x"79", x"7c", x"79", x"79", x"7b", x"7b", x"7c", x"7a", x"7b", 
        x"79", x"7c", x"7b", x"7c", x"7d", x"7a", x"79", x"79", x"7a", x"7b", x"7b", x"7a", x"79", x"7c", x"7d", 
        x"7d", x"7c", x"7b", x"7b", x"7c", x"7c", x"7c", x"7d", x"7e", x"7e", x"7e", x"7d", x"7c", x"7a", x"7b", 
        x"7b", x"7c", x"7c", x"7b", x"7c", x"7e", x"7d", x"7c", x"7c", x"7b", x"7a", x"7a", x"7b", x"7b", x"7a", 
        x"7b", x"7e", x"7d", x"7b", x"7c", x"7d", x"7e", x"7e", x"7e", x"7f", x"80", x"7d", x"7d", x"7d", x"7c", 
        x"7c", x"7c", x"7d", x"7d", x"7e", x"7f", x"7d", x"7f", x"7f", x"7b", x"7f", x"7e", x"7d", x"7e", x"7f", 
        x"7f", x"7f", x"7f", x"7e", x"7f", x"80", x"80", x"80", x"7f", x"7f", x"7e", x"80", x"81", x"7f", x"7c", 
        x"7e", x"81", x"82", x"7e", x"7e", x"7e", x"7d", x"7f", x"80", x"7e", x"80", x"81", x"80", x"84", x"87", 
        x"7a", x"68", x"80", x"bb", x"d6", x"d4", x"cc", x"9f", x"83", x"85", x"8b", x"8a", x"85", x"8c", x"86", 
        x"6a", x"ae", x"db", x"d1", x"d0", x"d1", x"d3", x"d8", x"ce", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", 
        x"cd", x"cc", x"cd", x"cf", x"ce", x"cd", x"ce", x"cf", x"ce", x"cf", x"cf", x"d1", x"d1", x"d2", x"d2", 
        x"d2", x"d1", x"d0", x"cf", x"cf", x"cf", x"cf", x"ce", x"ce", x"cf", x"cf", x"d0", x"cf", x"d0", x"d1", 
        x"d3", x"d2", x"cf", x"ce", x"cf", x"d0", x"d0", x"d1", x"dd", x"d1", x"d3", x"d4", x"d3", x"d3", x"d3", 
        x"dc", x"ef", x"ee", x"ed", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ec", 
        x"ec", x"ec", x"ec", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"ec", x"ed", x"ee", x"ef", x"ee", 
        x"ef", x"f0", x"ec", x"e3", x"cf", x"af", x"90", x"a6", x"c6", x"e2", x"e2", x"90", x"5e", x"5f", x"60", 
        x"6e", x"cf", x"f0", x"cc", x"8d", x"63", x"5d", x"5d", x"6f", x"a8", x"eb", x"f7", x"f5", x"c0", x"6a", 
        x"5c", x"5f", x"68", x"c8", x"f6", x"f9", x"f8", x"f4", x"ea", x"dd", x"c4", x"a0", x"7c", x"62", x"5c", 
        x"61", x"5e", x"5b", x"5e", x"5c", x"71", x"ca", x"f6", x"fa", x"fb", x"ee", x"a3", x"65", x"5d", x"5d", 
        x"7d", x"d8", x"ef", x"ee", x"ee", x"ef", x"ee", x"ed", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"ef", x"e6", x"d5", x"c2", x"b4", x"b8", x"d4", x"ec", 
        x"f2", x"f2", x"ef", x"ed", x"ee", x"f1", x"f2", x"ef", x"ee", x"ef", x"f0", x"f3", x"f4", x"f0", x"f2", 
        x"f3", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"eb", x"ee", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"f1", x"f1", x"eb", x"e0", x"d9", x"d6", x"dc", x"de", x"c2", x"95", x"74", x"73", 
        x"81", x"88", x"80", x"83", x"88", x"85", x"83", x"85", x"87", x"84", x"84", x"81", x"81", x"84", x"86", 
        x"86", x"85", x"84", x"85", x"86", x"87", x"86", x"84", x"84", x"84", x"83", x"84", x"84", x"86", x"86", 
        x"85", x"83", x"83", x"84", x"84", x"85", x"84", x"84", x"84", x"84", x"84", x"84", x"83", x"82", x"85", 
        x"84", x"84", x"85", x"84", x"82", x"83", x"84", x"83", x"82", x"82", x"82", x"83", x"84", x"87", x"85", 
        x"84", x"84", x"84", x"83", x"84", x"84", x"84", x"84", x"85", x"86", x"84", x"82", x"82", x"83", x"84", 
        x"83", x"84", x"83", x"83", x"84", x"85", x"83", x"82", x"84", x"85", x"83", x"81", x"81", x"83", x"82", 
        x"83", x"84", x"81", x"81", x"80", x"81", x"7e", x"80", x"84", x"81", x"81", x"80", x"7f", x"80", x"83", 
        x"82", x"81", x"82", x"82", x"80", x"7e", x"81", x"81", x"80", x"81", x"83", x"81", x"81", x"83", x"82", 
        x"80", x"80", x"82", x"83", x"81", x"80", x"81", x"82", x"82", x"82", x"81", x"80", x"7f", x"7e", x"7e", 
        x"7f", x"7f", x"81", x"81", x"80", x"7f", x"7f", x"80", x"82", x"81", x"80", x"7f", x"7e", x"7e", x"7f", 
        x"81", x"81", x"81", x"80", x"80", x"81", x"80", x"7f", x"7f", x"80", x"81", x"80", x"80", x"81", x"80", 
        x"7d", x"7f", x"7f", x"80", x"80", x"80", x"7f", x"7e", x"7f", x"80", x"80", x"80", x"80", x"7f", x"7e", 
        x"7f", x"7e", x"7f", x"7f", x"80", x"80", x"7e", x"7e", x"7f", x"7e", x"80", x"7f", x"80", x"7f", x"80", 
        x"7e", x"7e", x"7e", x"7f", x"80", x"7e", x"7e", x"7e", x"7d", x"7e", x"7d", x"7d", x"7e", x"80", x"7e", 
        x"7c", x"7b", x"7c", x"7e", x"7f", x"7f", x"7e", x"7f", x"80", x"7f", x"7e", x"7e", x"7f", x"7f", x"7e", 
        x"7d", x"7d", x"7d", x"7c", x"7c", x"7b", x"7c", x"7d", x"7b", x"7a", x"7b", x"7a", x"7a", x"7b", x"7b", 
        x"7b", x"7a", x"7b", x"7c", x"7c", x"7a", x"7a", x"7c", x"79", x"7a", x"7c", x"7b", x"7c", x"7a", x"79", 
        x"78", x"7b", x"7a", x"7b", x"7c", x"79", x"7a", x"7a", x"7a", x"7b", x"7a", x"7b", x"7b", x"7b", x"7c", 
        x"7c", x"7c", x"7c", x"7c", x"7d", x"7d", x"7c", x"7d", x"7d", x"7d", x"7c", x"7b", x"7c", x"7c", x"7c", 
        x"7c", x"7c", x"7c", x"7b", x"7c", x"7e", x"7e", x"7e", x"7d", x"7c", x"7b", x"7b", x"7b", x"7c", x"7b", 
        x"7b", x"7d", x"7e", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7d", x"7e", x"7f", x"7e", 
        x"7d", x"7e", x"80", x"7e", x"7d", x"7f", x"7d", x"7f", x"7e", x"7b", x"80", x"7e", x"7d", x"7e", x"80", 
        x"7f", x"7f", x"80", x"80", x"80", x"81", x"81", x"81", x"81", x"80", x"7b", x"7f", x"83", x"82", x"80", 
        x"7f", x"80", x"80", x"82", x"7f", x"80", x"83", x"80", x"82", x"81", x"7d", x"7f", x"85", x"81", x"71", 
        x"76", x"a2", x"cd", x"d4", x"cf", x"ce", x"cb", x"9d", x"85", x"8b", x"87", x"89", x"91", x"71", x"41", 
        x"32", x"ad", x"de", x"d3", x"d1", x"d0", x"d1", x"d5", x"ce", x"ce", x"cf", x"d0", x"d0", x"d0", x"cf", 
        x"ce", x"ce", x"ce", x"d0", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"d0", x"d1", x"d1", x"d2", x"d3", 
        x"d2", x"d1", x"d0", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"ce", x"d0", x"d0", x"d0", x"cf", 
        x"d1", x"d1", x"cf", x"cc", x"cd", x"cf", x"cf", x"d1", x"dc", x"cf", x"d1", x"d5", x"d4", x"d4", x"d2", 
        x"dc", x"ef", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", 
        x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ef", x"ee", x"ed", 
        x"ec", x"ee", x"f0", x"f2", x"ee", x"ef", x"e6", x"d7", x"c3", x"b6", x"a9", x"7f", x"63", x"5d", x"5c", 
        x"69", x"c5", x"f3", x"f2", x"e2", x"b4", x"85", x"6e", x"63", x"8c", x"e2", x"f9", x"f7", x"cc", x"72", 
        x"5d", x"5f", x"6a", x"c4", x"f3", x"f6", x"f6", x"f5", x"f7", x"f6", x"f6", x"ee", x"d0", x"88", x"5c", 
        x"5c", x"61", x"5f", x"61", x"5d", x"89", x"e0", x"f7", x"fa", x"fc", x"f9", x"c0", x"6e", x"5e", x"5d", 
        x"77", x"cf", x"ee", x"ed", x"ed", x"ee", x"ed", x"ec", x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"e3", x"d3", x"c3", x"b9", 
        x"c6", x"da", x"ea", x"f0", x"ee", x"ec", x"ef", x"f1", x"f0", x"f0", x"f4", x"f3", x"f0", x"f1", x"f2", 
        x"f2", x"f0", x"f1", x"f2", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"eb", x"ed", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f1", x"f2", x"f2", x"ee", x"e5", x"dc", x"d9", x"dd", x"df", x"cd", x"a5", 
        x"83", x"74", x"7c", x"80", x"82", x"86", x"88", x"86", x"84", x"88", x"88", x"85", x"86", x"86", x"86", 
        x"87", x"87", x"86", x"86", x"86", x"86", x"86", x"83", x"83", x"85", x"86", x"85", x"85", x"85", x"86", 
        x"85", x"84", x"84", x"84", x"85", x"85", x"84", x"83", x"84", x"85", x"85", x"84", x"83", x"84", x"85", 
        x"84", x"84", x"84", x"84", x"84", x"85", x"83", x"84", x"84", x"83", x"83", x"83", x"84", x"85", x"83", 
        x"82", x"84", x"83", x"82", x"83", x"84", x"84", x"85", x"85", x"86", x"85", x"84", x"83", x"82", x"83", 
        x"84", x"84", x"83", x"81", x"82", x"84", x"82", x"82", x"83", x"84", x"83", x"82", x"83", x"84", x"80", 
        x"82", x"83", x"81", x"83", x"80", x"82", x"80", x"81", x"82", x"80", x"82", x"83", x"81", x"81", x"84", 
        x"83", x"80", x"80", x"82", x"81", x"80", x"81", x"81", x"80", x"81", x"82", x"81", x"82", x"83", x"83", 
        x"7f", x"7f", x"82", x"81", x"81", x"81", x"81", x"82", x"81", x"80", x"80", x"80", x"81", x"82", x"82", 
        x"82", x"81", x"81", x"80", x"7f", x"7f", x"7f", x"80", x"80", x"81", x"81", x"7f", x"7f", x"7f", x"80", 
        x"81", x"82", x"81", x"80", x"80", x"81", x"80", x"7f", x"7d", x"7d", x"80", x"80", x"80", x"82", x"83", 
        x"81", x"81", x"80", x"7e", x"7e", x"7e", x"7f", x"80", x"7f", x"80", x"81", x"81", x"81", x"80", x"7f", 
        x"7f", x"7f", x"7f", x"80", x"81", x"80", x"7f", x"7d", x"7f", x"7e", x"80", x"7f", x"80", x"80", x"7f", 
        x"7d", x"7d", x"7e", x"7e", x"7f", x"7f", x"7f", x"80", x"7d", x"7d", x"7d", x"7d", x"7e", x"80", x"7f", 
        x"7d", x"7c", x"7e", x"7f", x"7e", x"7e", x"7c", x"7e", x"7e", x"7e", x"7c", x"7c", x"7e", x"82", x"83", 
        x"7e", x"7d", x"7c", x"7c", x"7c", x"7b", x"7a", x"7b", x"7a", x"79", x"7b", x"7b", x"7a", x"7b", x"7c", 
        x"7b", x"7a", x"7a", x"7b", x"7c", x"7b", x"7a", x"7a", x"79", x"7a", x"7b", x"7b", x"7c", x"7c", x"7d", 
        x"7c", x"7d", x"7c", x"7c", x"7d", x"7a", x"7b", x"7b", x"7b", x"7a", x"7b", x"7d", x"7d", x"7a", x"7a", 
        x"7c", x"7c", x"7c", x"7e", x"7f", x"7e", x"7e", x"7f", x"7f", x"7d", x"7d", x"7c", x"7b", x"7b", x"7b", 
        x"7b", x"7c", x"7d", x"7d", x"7d", x"7e", x"7d", x"7e", x"7e", x"7d", x"7d", x"7c", x"7b", x"7e", x"7d", 
        x"7c", x"7d", x"7e", x"7d", x"7c", x"7c", x"7c", x"7d", x"7d", x"7d", x"7e", x"7e", x"7f", x"7f", x"7e", 
        x"7e", x"7e", x"80", x"7f", x"7f", x"80", x"7f", x"80", x"7f", x"7c", x"7f", x"7e", x"7c", x"7e", x"7f", 
        x"7f", x"7e", x"80", x"81", x"80", x"80", x"80", x"81", x"82", x"81", x"7c", x"7e", x"82", x"83", x"81", 
        x"80", x"7f", x"84", x"7d", x"80", x"80", x"79", x"7b", x"7f", x"7d", x"83", x"88", x"7a", x"6a", x"89", 
        x"c8", x"d8", x"d3", x"ce", x"cd", x"d0", x"cd", x"9d", x"87", x"8c", x"8f", x"86", x"5a", x"2d", x"1e", 
        x"29", x"b0", x"e1", x"d5", x"d1", x"d0", x"d1", x"d5", x"ce", x"ce", x"d0", x"d1", x"d1", x"d0", x"cf", 
        x"d0", x"ce", x"ce", x"d0", x"d1", x"d0", x"d1", x"d0", x"d0", x"d0", x"d0", x"d1", x"d2", x"d2", x"d2", 
        x"d2", x"d1", x"d0", x"cf", x"cf", x"cf", x"d0", x"d0", x"cf", x"ce", x"cd", x"d0", x"d0", x"d1", x"cf", 
        x"d0", x"d1", x"d0", x"ce", x"cf", x"d0", x"cf", x"d1", x"dd", x"d0", x"d1", x"d4", x"d4", x"d4", x"d2", 
        x"dc", x"ef", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ed", x"ee", 
        x"ee", x"ed", x"ed", x"ec", x"ed", x"ee", x"eb", x"ef", x"ee", x"e9", x"da", x"bb", x"97", x"78", x"69", 
        x"68", x"a0", x"da", x"f2", x"f5", x"f2", x"e2", x"c7", x"bb", x"d1", x"f3", x"f9", x"f7", x"cb", x"72", 
        x"60", x"5e", x"66", x"be", x"f3", x"f9", x"ea", x"cc", x"d1", x"e6", x"f1", x"f5", x"e3", x"90", x"5d", 
        x"5f", x"5f", x"5d", x"5f", x"61", x"a7", x"ef", x"f8", x"f9", x"f9", x"fa", x"d9", x"7e", x"5c", x"5d", 
        x"73", x"c7", x"ed", x"ed", x"ed", x"ee", x"ed", x"ec", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ef", x"ed", x"eb", x"f1", x"f5", x"f0", x"ec", x"e2", 
        x"c9", x"b7", x"b6", x"cc", x"e2", x"eb", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f2", 
        x"f1", x"f0", x"f2", x"f1", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"eb", x"ed", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f2", x"f2", x"f0", x"ef", x"f0", x"f2", x"f3", x"f1", x"e8", x"dc", x"d7", x"db", x"e2", 
        x"d6", x"b0", x"85", x"77", x"7c", x"80", x"83", x"87", x"88", x"88", x"87", x"89", x"8a", x"85", x"89", 
        x"88", x"88", x"88", x"87", x"86", x"85", x"85", x"84", x"85", x"87", x"87", x"86", x"85", x"85", x"86", 
        x"85", x"83", x"84", x"85", x"85", x"85", x"84", x"83", x"84", x"84", x"85", x"85", x"85", x"85", x"85", 
        x"86", x"85", x"85", x"86", x"87", x"86", x"85", x"86", x"86", x"85", x"83", x"83", x"84", x"85", x"83", 
        x"84", x"86", x"85", x"84", x"85", x"83", x"83", x"83", x"84", x"84", x"85", x"86", x"84", x"82", x"84", 
        x"85", x"85", x"83", x"81", x"81", x"82", x"82", x"82", x"82", x"82", x"82", x"82", x"84", x"83", x"7f", 
        x"81", x"83", x"82", x"83", x"81", x"84", x"83", x"81", x"80", x"80", x"83", x"83", x"81", x"82", x"83", 
        x"82", x"80", x"80", x"82", x"81", x"81", x"82", x"82", x"80", x"7f", x"81", x"82", x"82", x"83", x"83", 
        x"80", x"80", x"81", x"80", x"80", x"80", x"82", x"82", x"80", x"7f", x"81", x"82", x"82", x"83", x"82", 
        x"81", x"80", x"80", x"7f", x"7e", x"7f", x"80", x"80", x"7e", x"80", x"81", x"81", x"81", x"81", x"81", 
        x"80", x"81", x"81", x"80", x"80", x"81", x"81", x"80", x"7f", x"81", x"81", x"80", x"80", x"81", x"81", 
        x"80", x"81", x"80", x"7e", x"7e", x"7f", x"7f", x"80", x"7f", x"80", x"80", x"80", x"80", x"80", x"7f", 
        x"7f", x"7f", x"7f", x"80", x"81", x"80", x"7f", x"7e", x"7f", x"7e", x"7f", x"7e", x"80", x"7f", x"7f", 
        x"7d", x"7d", x"7e", x"7e", x"7e", x"80", x"82", x"81", x"7d", x"7c", x"7d", x"7d", x"7d", x"7e", x"7e", 
        x"7e", x"7e", x"7e", x"7f", x"7e", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7d", x"7c", x"7d", 
        x"7d", x"7c", x"7b", x"7c", x"7d", x"7c", x"7a", x"7a", x"79", x"79", x"7b", x"7b", x"7b", x"7c", x"7c", 
        x"7b", x"7b", x"7b", x"7b", x"7c", x"7c", x"7a", x"7a", x"79", x"7a", x"7b", x"7b", x"7c", x"7d", x"7e", 
        x"7d", x"7e", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7c", x"7d", x"7e", x"7e", x"7b", x"7b", 
        x"7c", x"7c", x"7c", x"7e", x"7f", x"7d", x"7c", x"7d", x"7d", x"7c", x"7b", x"7b", x"7b", x"7b", x"7b", 
        x"7c", x"7c", x"7c", x"7e", x"7f", x"7f", x"7f", x"7e", x"7e", x"7d", x"7c", x"7c", x"7c", x"7f", x"7e", 
        x"7c", x"7d", x"7e", x"7e", x"80", x"80", x"7f", x"7f", x"7f", x"7e", x"7e", x"7d", x"7e", x"7e", x"7d", 
        x"7c", x"7d", x"7e", x"7f", x"7f", x"80", x"80", x"7f", x"7f", x"7d", x"7f", x"7e", x"7c", x"7e", x"7f", 
        x"7f", x"7e", x"7f", x"7f", x"7f", x"7f", x"80", x"80", x"81", x"81", x"80", x"80", x"80", x"81", x"80", 
        x"80", x"80", x"82", x"81", x"7f", x"82", x"82", x"7e", x"7f", x"81", x"7f", x"71", x"73", x"a4", x"d2", 
        x"d4", x"cf", x"cd", x"cd", x"cf", x"d0", x"cb", x"9f", x"8a", x"8c", x"70", x"3f", x"1f", x"17", x"16", 
        x"27", x"ae", x"de", x"d4", x"d2", x"d1", x"d3", x"d5", x"ce", x"ce", x"d1", x"d2", x"d2", x"d0", x"cf", 
        x"d0", x"ce", x"cd", x"d0", x"d1", x"d0", x"d0", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d2", 
        x"d2", x"d1", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"cf", x"cf", x"ce", x"d0", x"d0", x"d1", x"d0", 
        x"d2", x"d3", x"d2", x"d2", x"d1", x"d2", x"cf", x"d0", x"dd", x"d0", x"d0", x"d2", x"d4", x"d4", x"d2", 
        x"dc", x"ef", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"f0", x"f0", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ee", x"ee", 
        x"ee", x"ed", x"ed", x"ec", x"ec", x"ef", x"ee", x"f0", x"ed", x"ec", x"ee", x"ed", x"e5", x"d1", x"b4", 
        x"92", x"81", x"9b", x"c7", x"e5", x"ef", x"f5", x"f3", x"f3", x"f6", x"f3", x"f6", x"f1", x"bb", x"6d", 
        x"60", x"5f", x"68", x"bf", x"f3", x"f8", x"df", x"96", x"7c", x"98", x"b6", x"ce", x"d5", x"92", x"60", 
        x"5d", x"5e", x"5e", x"5c", x"6d", x"c4", x"f3", x"f6", x"eb", x"e1", x"f6", x"eb", x"9d", x"5f", x"5e", 
        x"6f", x"c1", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", x"f2", x"ee", x"ee", x"f0", x"ef", x"ee", x"f0", 
        x"ef", x"e8", x"d5", x"c0", x"b7", x"be", x"d5", x"e2", x"ec", x"f0", x"f1", x"f1", x"f0", x"f3", x"f1", 
        x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"eb", x"ed", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ea", x"e0", x"d8", 
        x"d9", x"de", x"d7", x"b6", x"8f", x"7b", x"7b", x"7f", x"86", x"85", x"86", x"88", x"88", x"84", x"86", 
        x"86", x"87", x"88", x"87", x"86", x"84", x"85", x"86", x"87", x"87", x"86", x"85", x"85", x"87", x"87", 
        x"86", x"84", x"84", x"86", x"87", x"85", x"84", x"85", x"86", x"86", x"87", x"86", x"86", x"84", x"83", 
        x"86", x"87", x"87", x"88", x"88", x"85", x"85", x"86", x"84", x"83", x"82", x"83", x"86", x"85", x"83", 
        x"85", x"87", x"87", x"85", x"85", x"83", x"83", x"84", x"84", x"82", x"83", x"85", x"84", x"83", x"84", 
        x"85", x"85", x"84", x"82", x"82", x"82", x"83", x"84", x"82", x"82", x"82", x"83", x"83", x"82", x"81", 
        x"84", x"85", x"83", x"80", x"83", x"84", x"83", x"82", x"82", x"81", x"82", x"81", x"80", x"81", x"82", 
        x"82", x"81", x"82", x"82", x"82", x"81", x"81", x"81", x"81", x"81", x"81", x"82", x"82", x"83", x"83", 
        x"82", x"81", x"81", x"81", x"80", x"80", x"81", x"82", x"81", x"80", x"81", x"81", x"80", x"7f", x"80", 
        x"80", x"80", x"80", x"80", x"7f", x"81", x"81", x"81", x"7f", x"7f", x"80", x"81", x"82", x"82", x"81", 
        x"80", x"81", x"82", x"81", x"81", x"81", x"81", x"81", x"80", x"7f", x"80", x"80", x"80", x"81", x"82", 
        x"81", x"7f", x"80", x"80", x"80", x"80", x"7f", x"7f", x"7f", x"80", x"80", x"80", x"80", x"80", x"80", 
        x"80", x"80", x"7f", x"80", x"81", x"80", x"7f", x"7f", x"80", x"7e", x"7d", x"7e", x"7f", x"7f", x"7f", 
        x"7e", x"7e", x"7e", x"7d", x"7e", x"80", x"82", x"81", x"7e", x"7d", x"7e", x"7f", x"7d", x"7c", x"7f", 
        x"7f", x"7f", x"7e", x"7e", x"7e", x"7d", x"7d", x"7c", x"7d", x"7d", x"7e", x"7d", x"7d", x"7c", x"7e", 
        x"7d", x"7c", x"7b", x"7d", x"7e", x"7d", x"7c", x"7b", x"79", x"7a", x"7c", x"7c", x"7b", x"7c", x"7c", 
        x"7b", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"7a", x"7a", x"7a", x"7b", x"7c", x"7c", x"7d", x"7c", 
        x"7c", x"7b", x"7b", x"7b", x"7a", x"7b", x"7a", x"7c", x"7f", x"7e", x"7d", x"7d", x"7e", x"7c", x"7d", 
        x"7e", x"7d", x"7d", x"7d", x"7e", x"7b", x"7b", x"7c", x"7c", x"7d", x"7d", x"7c", x"7c", x"7c", x"7d", 
        x"7d", x"7d", x"7d", x"7e", x"7e", x"7f", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7c", x"7f", x"7e", 
        x"7c", x"7e", x"7f", x"7e", x"7c", x"7c", x"7d", x"7f", x"81", x"82", x"82", x"7f", x"7e", x"7e", x"7d", 
        x"7d", x"7d", x"80", x"80", x"7f", x"7f", x"81", x"7f", x"7f", x"7e", x"7f", x"7e", x"7c", x"7e", x"80", 
        x"7f", x"7f", x"7f", x"7f", x"80", x"81", x"81", x"81", x"81", x"81", x"81", x"80", x"7f", x"7f", x"81", 
        x"82", x"82", x"81", x"81", x"7e", x"7b", x"7f", x"84", x"82", x"77", x"6d", x"8a", x"c9", x"dd", x"d0", 
        x"cb", x"cc", x"d2", x"d3", x"cb", x"d1", x"d5", x"a6", x"7c", x"51", x"20", x"13", x"18", x"16", x"18", 
        x"27", x"ac", x"dc", x"d4", x"d2", x"d1", x"d5", x"d5", x"ce", x"ce", x"d1", x"d2", x"d2", x"d0", x"cf", 
        x"cf", x"ce", x"cd", x"cf", x"d0", x"d0", x"d0", x"d1", x"d2", x"d1", x"d0", x"d0", x"d1", x"d2", x"d2", 
        x"d2", x"d1", x"d1", x"d0", x"d0", x"d1", x"d0", x"ce", x"cf", x"d0", x"d0", x"d2", x"d0", x"d1", x"d1", 
        x"d2", x"d3", x"d2", x"d2", x"d2", x"d2", x"cf", x"cf", x"dc", x"d1", x"d0", x"d2", x"d3", x"d4", x"d2", 
        x"dc", x"ef", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ed", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"f1", x"f1", x"ef", x"f0", x"ef", x"ef", x"ef", x"f2", 
        x"f0", x"d5", x"b1", x"a4", x"b2", x"cd", x"df", x"e9", x"f3", x"f9", x"f8", x"f2", x"cc", x"88", x"5b", 
        x"5e", x"5f", x"67", x"bd", x"f2", x"f7", x"e3", x"8e", x"58", x"5b", x"60", x"71", x"8d", x"78", x"61", 
        x"5e", x"5b", x"5e", x"5c", x"86", x"dc", x"f6", x"f4", x"c9", x"b3", x"f0", x"f6", x"c6", x"69", x"5f", 
        x"6b", x"bb", x"f0", x"f0", x"f0", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ef", x"f2", x"f3", x"f1", x"ef", x"f0", x"f0", x"ee", 
        x"ed", x"ef", x"f5", x"f4", x"e7", x"ce", x"b4", x"b3", x"c3", x"da", x"e7", x"ee", x"f3", x"f3", x"f2", 
        x"ef", x"ed", x"f0", x"f2", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"eb", x"ed", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f3", x"f3", x"f1", x"f2", x"f3", x"f4", x"f2", x"f3", x"f2", x"ef", x"f1", x"f4", x"f3", x"ee", 
        x"e4", x"d6", x"d7", x"e4", x"e9", x"c6", x"99", x"80", x"79", x"80", x"87", x"86", x"89", x"8d", x"8b", 
        x"85", x"86", x"87", x"87", x"86", x"85", x"86", x"86", x"87", x"88", x"87", x"85", x"86", x"88", x"87", 
        x"86", x"86", x"86", x"87", x"87", x"86", x"85", x"86", x"88", x"89", x"89", x"87", x"85", x"84", x"84", 
        x"85", x"84", x"84", x"86", x"87", x"85", x"84", x"84", x"83", x"83", x"83", x"85", x"86", x"84", x"82", 
        x"84", x"87", x"86", x"84", x"84", x"84", x"84", x"85", x"85", x"83", x"83", x"83", x"84", x"85", x"84", 
        x"83", x"83", x"83", x"84", x"84", x"83", x"85", x"85", x"84", x"82", x"83", x"85", x"82", x"81", x"83", 
        x"85", x"86", x"84", x"80", x"84", x"82", x"82", x"83", x"84", x"83", x"81", x"81", x"82", x"81", x"81", 
        x"81", x"82", x"82", x"82", x"82", x"81", x"80", x"80", x"82", x"83", x"83", x"83", x"83", x"83", x"83", 
        x"83", x"81", x"82", x"83", x"81", x"81", x"81", x"83", x"83", x"82", x"80", x"80", x"80", x"81", x"81", 
        x"82", x"82", x"82", x"81", x"81", x"82", x"82", x"82", x"81", x"80", x"80", x"82", x"82", x"82", x"81", 
        x"80", x"81", x"83", x"82", x"82", x"83", x"82", x"81", x"80", x"80", x"80", x"81", x"81", x"81", x"81", 
        x"82", x"80", x"80", x"80", x"80", x"80", x"7f", x"7f", x"80", x"80", x"80", x"7f", x"7f", x"80", x"80", 
        x"80", x"80", x"80", x"81", x"82", x"81", x"7f", x"81", x"80", x"7e", x"7d", x"7f", x"7f", x"7f", x"7f", 
        x"80", x"80", x"7f", x"7d", x"7d", x"7f", x"81", x"80", x"7f", x"7f", x"80", x"81", x"7e", x"7c", x"80", 
        x"80", x"7f", x"7e", x"7e", x"7f", x"80", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"80", x"80", 
        x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7a", x"7b", x"7e", x"7d", x"7b", x"7c", x"7c", 
        x"7c", x"7c", x"7c", x"7b", x"7b", x"7c", x"7d", x"7b", x"7b", x"7a", x"7b", x"7d", x"7c", x"7c", x"7c", 
        x"7d", x"7c", x"7d", x"7d", x"7c", x"7d", x"7b", x"7d", x"7f", x"7d", x"7b", x"7c", x"7d", x"7c", x"7d", 
        x"7e", x"7d", x"7c", x"7c", x"7d", x"7c", x"7b", x"7c", x"7d", x"7d", x"7d", x"7d", x"7d", x"7e", x"7e", 
        x"7e", x"7d", x"7d", x"7e", x"7d", x"7d", x"7d", x"7e", x"7e", x"7e", x"7f", x"7f", x"7e", x"7f", x"7e", 
        x"7d", x"7f", x"80", x"7e", x"7d", x"7d", x"7d", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", x"80", x"7f", 
        x"7e", x"7f", x"81", x"80", x"7e", x"7e", x"81", x"7f", x"7f", x"80", x"7f", x"7f", x"7d", x"7f", x"80", 
        x"80", x"7f", x"81", x"82", x"83", x"83", x"83", x"82", x"81", x"80", x"7e", x"7f", x"7f", x"80", x"81", 
        x"82", x"83", x"84", x"81", x"80", x"83", x"85", x"7d", x"6c", x"7f", x"ac", x"d2", x"d2", x"cc", x"cf", 
        x"cf", x"d0", x"cf", x"cb", x"d4", x"da", x"bf", x"74", x"33", x"1c", x"16", x"19", x"1d", x"1a", x"19", 
        x"28", x"af", x"dc", x"d4", x"d1", x"d1", x"d6", x"d5", x"ce", x"ce", x"cf", x"d0", x"d0", x"d0", x"cf", 
        x"cf", x"cd", x"cd", x"cf", x"d0", x"cf", x"d0", x"d2", x"d2", x"d0", x"cf", x"cf", x"d0", x"d1", x"d2", 
        x"d2", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"cf", x"cf", x"d0", x"d0", x"d2", x"d0", x"d1", x"d1", 
        x"d1", x"d1", x"d0", x"d0", x"d0", x"cf", x"d0", x"ce", x"db", x"d1", x"d1", x"d1", x"d3", x"d4", x"d2", 
        x"dc", x"ef", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ed", x"ef", x"ef", x"ef", x"f0", x"ef", x"ed", x"ee", x"f2", x"f1", x"ee", x"ef", x"f0", x"f2", x"f0", 
        x"eb", x"eb", x"ef", x"e5", x"db", x"d2", x"ca", x"ca", x"cb", x"c6", x"c0", x"b0", x"88", x"63", x"5f", 
        x"61", x"5e", x"65", x"b4", x"f2", x"fc", x"e5", x"94", x"58", x"58", x"5e", x"5a", x"5f", x"5d", x"5c", 
        x"5e", x"5f", x"5e", x"5c", x"a3", x"eb", x"f9", x"f0", x"a8", x"8c", x"e7", x"f7", x"e0", x"7c", x"5e", 
        x"6b", x"ba", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"f0", x"ee", x"ef", x"f1", x"f0", x"ee", 
        x"ef", x"f0", x"ee", x"ed", x"ef", x"f0", x"ec", x"dc", x"cb", x"be", x"bd", x"c5", x"d2", x"e8", x"f2", 
        x"f5", x"f2", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"eb", x"ed", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f3", x"f3", x"f3", x"f0", x"ef", x"f2", x"f3", x"f0", x"ed", x"f0", x"f4", 
        x"f1", x"ed", x"e6", x"de", x"dd", x"e0", x"dd", x"d0", x"af", x"8d", x"7c", x"78", x"7f", x"87", x"8a", 
        x"87", x"87", x"88", x"87", x"87", x"87", x"87", x"86", x"87", x"88", x"88", x"87", x"86", x"87", x"86", 
        x"86", x"87", x"87", x"87", x"86", x"86", x"86", x"87", x"88", x"89", x"8a", x"88", x"85", x"86", x"87", 
        x"85", x"83", x"83", x"84", x"87", x"87", x"85", x"84", x"84", x"86", x"87", x"86", x"86", x"87", x"86", 
        x"86", x"88", x"87", x"86", x"87", x"84", x"83", x"84", x"84", x"85", x"86", x"87", x"86", x"85", x"84", 
        x"83", x"83", x"83", x"84", x"84", x"84", x"85", x"86", x"84", x"84", x"84", x"85", x"84", x"82", x"84", 
        x"84", x"84", x"84", x"82", x"83", x"80", x"82", x"84", x"84", x"84", x"81", x"83", x"85", x"84", x"81", 
        x"81", x"83", x"82", x"81", x"82", x"82", x"80", x"80", x"83", x"84", x"83", x"83", x"84", x"82", x"82", 
        x"83", x"82", x"81", x"83", x"81", x"81", x"81", x"83", x"82", x"82", x"83", x"83", x"84", x"84", x"83", 
        x"82", x"81", x"81", x"82", x"82", x"82", x"81", x"81", x"82", x"81", x"81", x"82", x"82", x"82", x"81", 
        x"80", x"81", x"83", x"82", x"82", x"83", x"82", x"81", x"80", x"80", x"80", x"82", x"83", x"81", x"81", 
        x"83", x"82", x"81", x"80", x"7f", x"7f", x"80", x"81", x"81", x"80", x"7f", x"7f", x"7f", x"80", x"81", 
        x"80", x"80", x"80", x"81", x"82", x"81", x"80", x"80", x"7e", x"7d", x"7c", x"7f", x"7e", x"7d", x"7d", 
        x"80", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"80", x"81", x"80", x"80", x"82", x"80", x"7d", x"80", 
        x"81", x"80", x"7e", x"7e", x"7f", x"82", x"80", x"80", x"81", x"81", x"7f", x"7f", x"80", x"81", x"80", 
        x"7e", x"7f", x"7f", x"7e", x"7d", x"7c", x"7d", x"7d", x"7c", x"7d", x"7f", x"7d", x"7b", x"7b", x"7c", 
        x"7d", x"7c", x"7b", x"7a", x"7b", x"7d", x"7f", x"7c", x"7b", x"7a", x"7c", x"7f", x"7b", x"7b", x"7c", 
        x"7d", x"7b", x"7c", x"7c", x"7c", x"7f", x"7c", x"7d", x"7e", x"7b", x"79", x"7a", x"7d", x"7c", x"7d", 
        x"7e", x"7d", x"7d", x"7d", x"7e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7d", x"7e", x"7e", 
        x"7e", x"7e", x"7d", x"7d", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"7e", x"7f", x"7f", x"7f", x"7e", 
        x"7d", x"80", x"80", x"7e", x"7e", x"7e", x"7f", x"7f", x"80", x"80", x"80", x"7f", x"7f", x"7f", x"7e", 
        x"7e", x"7f", x"80", x"7f", x"7d", x"7d", x"81", x"7e", x"7e", x"81", x"7f", x"80", x"7e", x"80", x"81", 
        x"81", x"80", x"82", x"83", x"83", x"82", x"81", x"80", x"80", x"80", x"80", x"80", x"80", x"81", x"80", 
        x"81", x"82", x"81", x"82", x"84", x"83", x"76", x"72", x"8f", x"c1", x"d6", x"d0", x"cc", x"cf", x"d4", 
        x"d1", x"cf", x"d3", x"d5", x"d2", x"ac", x"5d", x"26", x"13", x"17", x"19", x"1a", x"1f", x"1a", x"16", 
        x"27", x"b2", x"dd", x"d3", x"d0", x"d1", x"d9", x"d8", x"ce", x"cd", x"ce", x"cf", x"cf", x"d0", x"d0", 
        x"cf", x"ce", x"cf", x"d1", x"d0", x"cf", x"d1", x"d2", x"d2", x"d0", x"ce", x"ce", x"cf", x"d1", x"d2", 
        x"d2", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d0", x"d0", x"d0", x"cf", x"d1", x"d1", x"d2", x"d3", 
        x"d2", x"d1", x"d0", x"d0", x"cf", x"cf", x"d0", x"cd", x"da", x"d0", x"d2", x"d2", x"d2", x"d4", x"d2", 
        x"dc", x"ef", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ed", x"ed", x"eb", x"ef", x"f0", x"ef", x"f0", x"ed", x"ec", x"ef", x"f0", x"eb", x"ef", 
        x"ef", x"ed", x"ef", x"ee", x"f0", x"f2", x"eb", x"de", x"cb", x"b4", x"9e", x"7c", x"63", x"5f", x"69", 
        x"65", x"5e", x"63", x"b2", x"f1", x"fa", x"ed", x"bb", x"87", x"6d", x"62", x"5d", x"5b", x"5e", x"5e", 
        x"5d", x"60", x"5e", x"64", x"c0", x"f4", x"fa", x"e6", x"92", x"72", x"d6", x"f4", x"f0", x"97", x"61", 
        x"6d", x"b6", x"ee", x"ee", x"ef", x"ef", x"ee", x"ed", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f0", x"f0", x"f2", x"ef", x"f1", x"f1", x"ee", x"ef", 
        x"f1", x"f0", x"ee", x"ee", x"ee", x"ee", x"f2", x"f4", x"f0", x"e6", x"d3", x"c2", x"b8", x"c0", x"cb", 
        x"de", x"f1", x"f3", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"eb", x"ed", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", 
        x"f0", x"ee", x"f2", x"f2", x"eb", x"e2", x"e2", x"e6", x"e2", x"d2", x"b3", x"8f", x"7d", x"7b", x"83", 
        x"8a", x"8a", x"89", x"88", x"89", x"88", x"88", x"86", x"86", x"87", x"87", x"87", x"87", x"88", x"86", 
        x"86", x"88", x"89", x"87", x"85", x"87", x"87", x"87", x"88", x"89", x"89", x"88", x"87", x"88", x"87", 
        x"86", x"87", x"88", x"86", x"85", x"87", x"89", x"87", x"85", x"87", x"88", x"88", x"87", x"89", x"88", 
        x"87", x"88", x"87", x"86", x"88", x"88", x"86", x"84", x"84", x"85", x"86", x"86", x"86", x"85", x"84", 
        x"84", x"84", x"84", x"83", x"84", x"84", x"85", x"85", x"84", x"84", x"84", x"85", x"84", x"82", x"85", 
        x"84", x"83", x"85", x"82", x"80", x"7f", x"85", x"85", x"82", x"83", x"82", x"83", x"85", x"84", x"81", 
        x"82", x"84", x"84", x"82", x"83", x"83", x"81", x"81", x"82", x"82", x"81", x"83", x"84", x"82", x"82", 
        x"84", x"83", x"81", x"81", x"80", x"80", x"81", x"82", x"81", x"80", x"83", x"83", x"83", x"83", x"82", 
        x"81", x"81", x"81", x"81", x"82", x"80", x"7e", x"7f", x"83", x"82", x"81", x"82", x"82", x"82", x"81", 
        x"81", x"82", x"83", x"82", x"82", x"83", x"83", x"82", x"81", x"7e", x"7f", x"82", x"84", x"82", x"81", 
        x"82", x"81", x"81", x"81", x"80", x"80", x"80", x"80", x"80", x"80", x"7f", x"7f", x"7f", x"80", x"81", 
        x"80", x"80", x"80", x"81", x"81", x"81", x"80", x"80", x"7e", x"7e", x"7d", x"81", x"7f", x"7d", x"7c", 
        x"7f", x"7e", x"7f", x"80", x"80", x"80", x"7f", x"81", x"82", x"80", x"7f", x"81", x"82", x"80", x"7f", 
        x"80", x"81", x"80", x"7f", x"80", x"82", x"80", x"81", x"81", x"80", x"7e", x"7e", x"7f", x"79", x"77", 
        x"7e", x"7e", x"7e", x"7c", x"7b", x"7b", x"7d", x"7e", x"7c", x"7c", x"7d", x"7c", x"7a", x"7c", x"7e", 
        x"7d", x"7c", x"7b", x"79", x"7b", x"7d", x"7e", x"7e", x"7d", x"7b", x"7b", x"7c", x"79", x"79", x"7c", 
        x"7b", x"7b", x"7d", x"7c", x"7b", x"7f", x"7d", x"7e", x"7d", x"7e", x"7b", x"7d", x"7d", x"7e", x"7d", 
        x"7c", x"7c", x"7e", x"7e", x"7d", x"7e", x"7e", x"7e", x"7e", x"7f", x"7e", x"7d", x"7d", x"7d", x"7e", 
        x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"7f", x"7d", x"7e", x"80", x"7d", x"7e", x"7f", 
        x"80", x"80", x"7f", x"7d", x"7f", x"80", x"81", x"81", x"80", x"80", x"7f", x"7d", x"7d", x"7e", x"7f", 
        x"7f", x"7e", x"7f", x"7d", x"7e", x"7e", x"80", x"7f", x"7f", x"81", x"80", x"81", x"7f", x"7f", x"82", 
        x"81", x"7f", x"80", x"80", x"81", x"7f", x"7e", x"7f", x"80", x"80", x"83", x"82", x"82", x"82", x"80", 
        x"81", x"80", x"84", x"8a", x"7a", x"64", x"86", x"b7", x"d6", x"d2", x"ce", x"cf", x"d0", x"ce", x"ce", 
        x"ce", x"d1", x"df", x"bc", x"6e", x"30", x"1a", x"18", x"17", x"19", x"1a", x"1b", x"17", x"16", x"19", 
        x"26", x"ad", x"db", x"d1", x"d1", x"d3", x"d8", x"d8", x"ce", x"cd", x"ce", x"cf", x"d0", x"d0", x"d0", 
        x"ce", x"ce", x"d1", x"d2", x"d1", x"cf", x"d1", x"d1", x"cf", x"cf", x"cf", x"d0", x"cf", x"d1", x"d2", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"d1", x"d3", 
        x"d2", x"d2", x"d0", x"cf", x"ce", x"cd", x"d0", x"cf", x"da", x"d0", x"d1", x"d1", x"d1", x"d3", x"d0", 
        x"da", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ed", 
        x"ed", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ed", x"ee", x"f0", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ed", x"ef", 
        x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"ec", x"e1", x"cb", x"af", x"92", x"73", 
        x"65", x"61", x"67", x"b2", x"f0", x"f9", x"f8", x"f1", x"e3", x"c9", x"ae", x"8f", x"6e", x"62", x"5d", 
        x"60", x"5e", x"5b", x"78", x"d7", x"f5", x"f8", x"d6", x"7b", x"5c", x"b3", x"ed", x"f7", x"b9", x"63", 
        x"6d", x"b6", x"ec", x"ee", x"f1", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ee", x"ef", x"f2", x"f0", x"ee", 
        x"ef", x"f1", x"f1", x"ef", x"ee", x"ef", x"f2", x"f0", x"f0", x"f1", x"f2", x"ee", x"e5", x"d4", x"c3", 
        x"b6", x"ba", x"ce", x"e5", x"f4", x"f2", x"f1", x"ef", x"ee", x"ef", x"f1", x"f0", x"ef", x"f0", x"f2", 
        x"f1", x"f0", x"f4", x"f3", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ec", x"ed", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f2", x"f2", x"f0", x"ef", 
        x"ef", x"f0", x"f1", x"f1", x"f1", x"f3", x"ef", x"e7", x"df", x"e3", x"e3", x"de", x"c5", x"9f", x"81", 
        x"76", x"7d", x"86", x"8c", x"89", x"85", x"86", x"87", x"87", x"87", x"87", x"88", x"89", x"8a", x"87", 
        x"87", x"88", x"87", x"86", x"87", x"88", x"87", x"87", x"88", x"86", x"85", x"86", x"86", x"86", x"86", 
        x"85", x"86", x"88", x"87", x"85", x"85", x"87", x"87", x"85", x"86", x"88", x"86", x"87", x"87", x"87", 
        x"86", x"86", x"87", x"88", x"87", x"87", x"86", x"85", x"84", x"84", x"85", x"85", x"87", x"86", x"86", 
        x"87", x"83", x"83", x"83", x"83", x"87", x"86", x"86", x"85", x"84", x"84", x"84", x"85", x"85", x"85", 
        x"85", x"86", x"85", x"86", x"82", x"81", x"83", x"83", x"81", x"83", x"83", x"83", x"82", x"83", x"85", 
        x"84", x"82", x"82", x"81", x"81", x"82", x"81", x"82", x"83", x"83", x"82", x"83", x"84", x"84", x"85", 
        x"84", x"82", x"81", x"81", x"82", x"82", x"83", x"83", x"82", x"81", x"81", x"81", x"80", x"80", x"81", 
        x"81", x"82", x"80", x"81", x"82", x"81", x"80", x"80", x"82", x"83", x"83", x"83", x"83", x"83", x"83", 
        x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"82", x"81", x"80", x"80", x"81", x"83", x"82", x"81", 
        x"81", x"80", x"82", x"82", x"80", x"80", x"81", x"80", x"82", x"82", x"82", x"81", x"80", x"81", x"81", 
        x"82", x"82", x"81", x"80", x"81", x"82", x"82", x"82", x"80", x"80", x"80", x"82", x"7f", x"80", x"80", 
        x"81", x"7f", x"7f", x"80", x"81", x"81", x"7f", x"7f", x"81", x"80", x"81", x"82", x"81", x"80", x"7f", 
        x"80", x"81", x"80", x"80", x"7f", x"7f", x"83", x"82", x"7f", x"7f", x"7c", x"78", x"78", x"80", x"87", 
        x"80", x"80", x"80", x"7d", x"7c", x"7c", x"7d", x"7d", x"7b", x"7a", x"7c", x"7c", x"7b", x"7e", x"80", 
        x"7d", x"7c", x"7c", x"7b", x"7d", x"7c", x"7b", x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", x"7d", x"7e", 
        x"7c", x"7d", x"7e", x"7c", x"7c", x"7e", x"7d", x"7e", x"7d", x"80", x"7d", x"7e", x"7d", x"7f", x"7e", 
        x"7c", x"7c", x"7f", x"7f", x"7c", x"7b", x"7d", x"7f", x"80", x"80", x"7f", x"7d", x"7c", x"7e", x"7e", 
        x"7e", x"7f", x"7f", x"7f", x"80", x"7f", x"7d", x"7e", x"80", x"7e", x"7e", x"7e", x"7d", x"7e", x"7f", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7c", x"7d", x"7f", x"80", 
        x"7f", x"7f", x"7e", x"7e", x"7e", x"7f", x"80", x"7f", x"7f", x"80", x"80", x"81", x"81", x"80", x"83", 
        x"81", x"7f", x"80", x"80", x"81", x"7f", x"7f", x"81", x"83", x"82", x"80", x"83", x"82", x"80", x"80", 
        x"81", x"8a", x"86", x"6e", x"75", x"a2", x"c9", x"d5", x"d0", x"cd", x"ce", x"ce", x"d1", x"d1", x"d1", 
        x"d7", x"c8", x"93", x"48", x"21", x"18", x"16", x"19", x"1b", x"18", x"18", x"19", x"16", x"15", x"18", 
        x"24", x"ad", x"dc", x"d1", x"d2", x"d3", x"d5", x"d6", x"ce", x"cd", x"cf", x"d0", x"d0", x"d0", x"cf", 
        x"ce", x"cf", x"d1", x"d3", x"d1", x"cf", x"d1", x"d1", x"ce", x"ce", x"d0", x"d1", x"d0", x"d1", x"d2", 
        x"d0", x"d0", x"d1", x"d1", x"d2", x"d3", x"d2", x"d0", x"d0", x"cf", x"cf", x"d0", x"d2", x"d3", x"d3", 
        x"d2", x"d2", x"d1", x"d0", x"cf", x"cf", x"d0", x"cf", x"db", x"d0", x"d2", x"d2", x"d2", x"d3", x"cf", 
        x"d9", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f1", x"f0", x"ef", x"ee", x"f0", x"f2", x"f2", x"f0", x"eb", x"df", x"c5", 
        x"ae", x"95", x"7d", x"9b", x"d1", x"e7", x"f1", x"f6", x"fb", x"f7", x"ed", x"e1", x"ca", x"a2", x"6d", 
        x"5d", x"5e", x"60", x"9b", x"e9", x"f7", x"f9", x"e4", x"af", x"88", x"a8", x"e5", x"fa", x"d5", x"76", 
        x"6d", x"b2", x"eb", x"ee", x"f1", x"f0", x"ef", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"f2", x"f3", x"f2", x"e9", 
        x"df", x"d0", x"c0", x"ba", x"c1", x"d9", x"e7", x"f0", x"f2", x"f0", x"f0", x"f0", x"f1", x"f1", x"f3", 
        x"f2", x"ef", x"f0", x"ee", x"ee", x"f0", x"ef", x"f0", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"ed", x"ed", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f0", x"ef", x"ee", x"ee", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"ed", x"ea", x"e5", x"e4", x"e6", x"e0", x"cc", 
        x"a8", x"8c", x"7a", x"7e", x"86", x"89", x"89", x"87", x"87", x"88", x"88", x"87", x"88", x"88", x"88", 
        x"88", x"87", x"85", x"86", x"88", x"88", x"86", x"85", x"87", x"86", x"85", x"86", x"87", x"87", x"88", 
        x"87", x"87", x"87", x"87", x"86", x"85", x"85", x"85", x"84", x"85", x"87", x"87", x"89", x"86", x"87", 
        x"86", x"86", x"88", x"89", x"86", x"83", x"84", x"85", x"85", x"86", x"86", x"87", x"88", x"86", x"86", 
        x"87", x"83", x"84", x"85", x"83", x"85", x"85", x"85", x"85", x"86", x"86", x"86", x"86", x"86", x"82", 
        x"84", x"86", x"84", x"85", x"85", x"83", x"82", x"81", x"82", x"83", x"84", x"83", x"81", x"82", x"86", 
        x"85", x"80", x"80", x"82", x"82", x"82", x"82", x"82", x"83", x"83", x"83", x"83", x"83", x"82", x"82", 
        x"82", x"82", x"83", x"84", x"84", x"83", x"82", x"82", x"82", x"81", x"81", x"82", x"83", x"84", x"83", 
        x"82", x"81", x"80", x"81", x"82", x"82", x"81", x"81", x"82", x"84", x"84", x"84", x"83", x"82", x"81", 
        x"81", x"81", x"82", x"82", x"82", x"82", x"82", x"82", x"82", x"81", x"81", x"81", x"82", x"83", x"83", 
        x"82", x"80", x"83", x"82", x"7f", x"7f", x"81", x"80", x"82", x"82", x"82", x"81", x"81", x"81", x"81", 
        x"82", x"81", x"80", x"7f", x"7f", x"7f", x"80", x"82", x"80", x"80", x"82", x"82", x"7f", x"80", x"81", 
        x"7f", x"80", x"81", x"82", x"82", x"80", x"80", x"83", x"83", x"7f", x"7f", x"80", x"7f", x"80", x"80", 
        x"81", x"81", x"81", x"81", x"81", x"80", x"85", x"7e", x"78", x"7d", x"85", x"87", x"8c", x"92", x"96", 
        x"7e", x"7f", x"7f", x"7f", x"7f", x"80", x"82", x"7e", x"7a", x"7a", x"7c", x"7d", x"7c", x"7f", x"7f", 
        x"7c", x"7c", x"7e", x"7c", x"7d", x"7c", x"7b", x"7c", x"7d", x"7c", x"7d", x"7d", x"7e", x"7e", x"7d", 
        x"7b", x"7c", x"7d", x"7d", x"7c", x"7e", x"7c", x"7d", x"7d", x"7f", x"7d", x"7e", x"7d", x"7e", x"7e", 
        x"7c", x"7c", x"7e", x"7f", x"7c", x"7c", x"7e", x"7e", x"7d", x"7d", x"7d", x"7e", x"7f", x"7f", x"7f", 
        x"7e", x"7f", x"7e", x"7e", x"80", x"81", x"7c", x"7d", x"80", x"81", x"7e", x"7c", x"7f", x"7e", x"7e", 
        x"7d", x"7e", x"80", x"81", x"80", x"7f", x"7e", x"7e", x"7e", x"7f", x"80", x"7d", x"7e", x"7f", x"80", 
        x"80", x"7f", x"7f", x"7e", x"7e", x"7f", x"80", x"7f", x"7f", x"80", x"81", x"82", x"83", x"81", x"82", 
        x"81", x"81", x"82", x"81", x"83", x"81", x"80", x"83", x"84", x"83", x"83", x"84", x"80", x"82", x"87", 
        x"88", x"7c", x"69", x"89", x"bc", x"d5", x"d1", x"d0", x"cf", x"cc", x"cb", x"cb", x"d1", x"d4", x"da", 
        x"ad", x"5e", x"26", x"1a", x"1d", x"19", x"1a", x"1d", x"18", x"18", x"17", x"19", x"16", x"17", x"17", 
        x"25", x"af", x"de", x"d3", x"d2", x"d2", x"d4", x"d6", x"ce", x"ce", x"cf", x"d0", x"d0", x"cf", x"ce", 
        x"d0", x"cf", x"d1", x"d2", x"d1", x"cf", x"d2", x"d2", x"cf", x"cf", x"d0", x"d0", x"cf", x"d0", x"d2", 
        x"d3", x"d2", x"d2", x"d1", x"d2", x"d3", x"d2", x"d2", x"d1", x"d0", x"d0", x"d1", x"d3", x"d4", x"d2", 
        x"d1", x"d0", x"d0", x"cf", x"d0", x"d0", x"ce", x"ce", x"da", x"d1", x"d2", x"d4", x"d4", x"d4", x"cf", 
        x"d9", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f2", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ed", x"ef", x"f1", x"f1", 
        x"ee", x"e3", x"d0", x"be", x"af", x"a0", x"b7", x"d7", x"ee", x"f4", x"f8", x"f9", x"f5", x"d0", x"80", 
        x"59", x"5d", x"67", x"b9", x"f3", x"fa", x"fa", x"f3", x"ec", x"de", x"dd", x"f0", x"fc", x"e8", x"98", 
        x"6e", x"ae", x"ea", x"ee", x"f1", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f2", x"f2", x"ef", x"f3", 
        x"f5", x"f2", x"ea", x"de", x"cd", x"b1", x"b2", x"c6", x"e4", x"f2", x"f2", x"f0", x"f1", x"f2", x"f2", 
        x"ee", x"ef", x"f6", x"f2", x"f0", x"f1", x"ef", x"f0", x"f1", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"ed", x"ed", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"ef", x"ee", x"ef", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f4", x"f1", x"ec", x"ea", x"e5", x"e0", 
        x"e7", x"da", x"b9", x"8a", x"72", x"75", x"86", x"88", x"85", x"84", x"87", x"8c", x"8d", x"89", x"84", 
        x"82", x"84", x"87", x"88", x"89", x"88", x"87", x"86", x"89", x"88", x"87", x"88", x"87", x"87", x"8a", 
        x"89", x"89", x"87", x"87", x"86", x"87", x"89", x"87", x"86", x"85", x"84", x"86", x"86", x"86", x"87", 
        x"88", x"87", x"88", x"87", x"84", x"83", x"85", x"86", x"86", x"85", x"85", x"86", x"88", x"87", x"87", 
        x"87", x"83", x"83", x"83", x"83", x"85", x"85", x"85", x"85", x"86", x"86", x"86", x"86", x"85", x"82", 
        x"83", x"85", x"83", x"83", x"86", x"86", x"83", x"82", x"83", x"85", x"87", x"84", x"81", x"82", x"85", 
        x"84", x"81", x"81", x"83", x"83", x"82", x"81", x"81", x"82", x"83", x"84", x"84", x"82", x"81", x"80", 
        x"81", x"82", x"83", x"86", x"85", x"83", x"82", x"82", x"82", x"82", x"81", x"83", x"84", x"86", x"84", 
        x"83", x"81", x"83", x"82", x"82", x"82", x"82", x"82", x"82", x"83", x"83", x"82", x"82", x"82", x"81", 
        x"81", x"81", x"82", x"82", x"82", x"82", x"82", x"82", x"82", x"82", x"82", x"82", x"83", x"83", x"83", 
        x"83", x"80", x"82", x"82", x"80", x"80", x"80", x"7f", x"81", x"81", x"81", x"81", x"81", x"81", x"81", 
        x"82", x"82", x"80", x"80", x"7f", x"7f", x"7e", x"80", x"80", x"80", x"81", x"81", x"7f", x"80", x"80", 
        x"7f", x"80", x"82", x"82", x"81", x"80", x"81", x"83", x"84", x"81", x"81", x"81", x"7f", x"81", x"80", 
        x"81", x"81", x"82", x"82", x"7b", x"73", x"75", x"81", x"8c", x"92", x"94", x"94", x"a0", x"b7", x"c3", 
        x"7e", x"7e", x"7e", x"7d", x"7c", x"7c", x"7d", x"7e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7d", x"7e", 
        x"7c", x"7c", x"7e", x"7e", x"7f", x"7f", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7b", 
        x"7a", x"7b", x"7d", x"7e", x"7f", x"80", x"7c", x"7d", x"7d", x"7e", x"7d", x"7d", x"7d", x"7d", x"7f", 
        x"7d", x"7c", x"7e", x"7f", x"7c", x"7d", x"7e", x"7e", x"7c", x"7b", x"7c", x"7f", x"80", x"80", x"80", 
        x"7f", x"7f", x"7e", x"7e", x"7f", x"80", x"7d", x"7d", x"81", x"82", x"7f", x"7d", x"80", x"7f", x"7d", 
        x"7c", x"7c", x"7c", x"7e", x"80", x"7f", x"7e", x"7e", x"7e", x"7f", x"80", x"7e", x"7e", x"7f", x"80", 
        x"81", x"80", x"80", x"80", x"80", x"81", x"81", x"81", x"81", x"81", x"81", x"82", x"83", x"81", x"81", 
        x"81", x"82", x"83", x"82", x"84", x"83", x"81", x"83", x"83", x"81", x"80", x"84", x"82", x"83", x"83", 
        x"75", x"73", x"ae", x"cc", x"d4", x"cf", x"ce", x"cf", x"ce", x"cf", x"cc", x"d3", x"db", x"c4", x"82", 
        x"34", x"1b", x"18", x"19", x"1b", x"19", x"1a", x"1b", x"1a", x"18", x"16", x"17", x"19", x"1b", x"18", 
        x"27", x"b0", x"de", x"d2", x"d2", x"d1", x"d4", x"d6", x"cd", x"cd", x"cf", x"d0", x"d0", x"cf", x"cf", 
        x"d1", x"d1", x"d1", x"d2", x"d0", x"cf", x"d2", x"d3", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"d2", 
        x"d4", x"d3", x"d3", x"d2", x"d1", x"d0", x"d0", x"d0", x"d1", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", 
        x"d2", x"d0", x"ce", x"cd", x"cd", x"ce", x"cd", x"cd", x"da", x"d1", x"d2", x"d4", x"d4", x"d4", x"cf", 
        x"d9", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"ef", x"ed", x"ec", x"ef", x"ef", x"ee", x"ec", 
        x"ed", x"f0", x"f0", x"eb", x"e5", x"d6", x"b6", x"9f", x"9e", x"b6", x"d6", x"e5", x"ed", x"d2", x"83", 
        x"59", x"5b", x"77", x"d1", x"f6", x"f9", x"f5", x"eb", x"ee", x"f4", x"f6", x"f7", x"f9", x"f0", x"b5", 
        x"6e", x"a7", x"e9", x"ef", x"f0", x"ee", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"ee", x"ee", x"f0", x"f1", x"f2", x"f2", x"f1", x"ef", 
        x"ed", x"ee", x"f1", x"f2", x"ee", x"e5", x"d7", x"c1", x"b3", x"ba", x"cf", x"e5", x"ec", x"ee", x"f0", 
        x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"ee", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"ed", x"ed", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f3", x"f0", x"ea", 
        x"e5", x"e6", x"e7", x"dd", x"c0", x"9a", x"78", x"7a", x"83", x"88", x"87", x"87", x"89", x"89", x"89", 
        x"87", x"88", x"87", x"85", x"84", x"88", x"89", x"88", x"89", x"88", x"88", x"88", x"87", x"86", x"89", 
        x"89", x"88", x"87", x"85", x"86", x"87", x"88", x"86", x"88", x"86", x"85", x"88", x"85", x"85", x"87", 
        x"87", x"87", x"88", x"88", x"85", x"85", x"88", x"89", x"87", x"84", x"82", x"84", x"85", x"84", x"85", 
        x"86", x"85", x"86", x"87", x"87", x"87", x"86", x"86", x"85", x"85", x"85", x"85", x"87", x"85", x"83", 
        x"84", x"85", x"83", x"82", x"86", x"86", x"84", x"83", x"83", x"86", x"87", x"85", x"82", x"82", x"84", 
        x"84", x"82", x"83", x"84", x"83", x"83", x"83", x"83", x"83", x"83", x"84", x"85", x"85", x"85", x"84", 
        x"83", x"83", x"84", x"85", x"84", x"83", x"83", x"83", x"83", x"84", x"84", x"84", x"84", x"84", x"84", 
        x"84", x"84", x"85", x"83", x"82", x"82", x"83", x"83", x"83", x"82", x"82", x"82", x"82", x"82", x"83", 
        x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", 
        x"83", x"81", x"82", x"82", x"82", x"81", x"81", x"80", x"80", x"80", x"81", x"81", x"81", x"81", x"82", 
        x"82", x"83", x"83", x"83", x"82", x"82", x"81", x"81", x"81", x"81", x"81", x"81", x"80", x"80", x"81", 
        x"81", x"82", x"81", x"7f", x"7f", x"80", x"82", x"83", x"84", x"83", x"83", x"82", x"7f", x"82", x"80", 
        x"81", x"80", x"7d", x"7b", x"82", x"8b", x"98", x"9c", x"9f", x"ab", x"bc", x"c6", x"d2", x"d4", x"d2", 
        x"7d", x"7e", x"7e", x"7d", x"7b", x"7b", x"7b", x"7c", x"7e", x"7e", x"7d", x"7e", x"7e", x"7d", x"80", 
        x"7e", x"7d", x"7d", x"7c", x"7f", x"7f", x"7e", x"7e", x"7e", x"7f", x"7e", x"7e", x"7e", x"7d", x"7c", 
        x"7c", x"7c", x"7c", x"7e", x"7f", x"7f", x"7d", x"7d", x"7e", x"7e", x"7e", x"7d", x"7d", x"7e", x"7f", 
        x"7e", x"7d", x"7e", x"80", x"7e", x"7b", x"7d", x"7f", x"80", x"7f", x"7d", x"7d", x"7f", x"80", x"80", 
        x"7f", x"7f", x"7e", x"7e", x"7d", x"7e", x"7f", x"7f", x"7f", x"80", x"81", x"81", x"81", x"80", x"7f", 
        x"7f", x"7e", x"7d", x"7e", x"7e", x"7f", x"7e", x"7e", x"7e", x"7f", x"7f", x"7e", x"7e", x"80", x"81", 
        x"81", x"81", x"80", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"80", x"80", x"81", x"81", x"7f", 
        x"80", x"83", x"83", x"83", x"84", x"82", x"81", x"82", x"82", x"81", x"84", x"89", x"87", x"79", x"6b", 
        x"94", x"d2", x"d9", x"d4", x"d1", x"cd", x"cd", x"cf", x"cf", x"d1", x"d6", x"d3", x"a5", x"53", x"1f", 
        x"1b", x"1c", x"1e", x"1b", x"1a", x"1d", x"1b", x"19", x"1b", x"18", x"19", x"1b", x"1a", x"19", x"14", 
        x"25", x"ac", x"dd", x"d1", x"d0", x"d1", x"d4", x"d8", x"cd", x"cc", x"ce", x"d0", x"d0", x"d0", x"d0", 
        x"d2", x"d1", x"d1", x"d2", x"d0", x"cf", x"d1", x"d2", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"d0", 
        x"d0", x"d1", x"d2", x"d2", x"d1", x"d0", x"cf", x"cf", x"d0", x"d1", x"d1", x"d1", x"d2", x"d3", x"d5", 
        x"d4", x"d2", x"d0", x"cf", x"cf", x"d0", x"cf", x"cf", x"db", x"d1", x"d2", x"d4", x"d3", x"d3", x"cf", 
        x"d9", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f1", x"f0", x"ef", x"ee", x"f0", x"ee", x"ec", x"ed", 
        x"ee", x"ed", x"ef", x"f1", x"ef", x"ef", x"ed", x"ea", x"d6", x"b4", x"9f", x"9f", x"b4", x"b7", x"87", 
        x"60", x"60", x"97", x"e6", x"f4", x"f4", x"d5", x"a3", x"b7", x"d4", x"e8", x"f2", x"f7", x"f5", x"d8", 
        x"82", x"98", x"e7", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ee", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"ee", x"ee", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", 
        x"f4", x"f5", x"f1", x"ef", x"f2", x"f0", x"f1", x"f1", x"e4", x"cd", x"b8", x"ad", x"bf", x"d7", x"e8", 
        x"ee", x"f1", x"f5", x"f4", x"f3", x"f2", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"ed", x"ed", x"f0", x"ef", x"f0", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"ef", x"ef", x"ef", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f0", x"ef", x"f0", x"f4", 
        x"f3", x"ed", x"e4", x"e1", x"e6", x"e2", x"ce", x"a2", x"83", x"77", x"81", x"88", x"88", x"8a", x"8b", 
        x"89", x"87", x"86", x"85", x"84", x"86", x"88", x"86", x"87", x"85", x"86", x"88", x"89", x"87", x"87", 
        x"88", x"88", x"87", x"86", x"87", x"89", x"89", x"87", x"89", x"87", x"86", x"87", x"85", x"85", x"87", 
        x"86", x"85", x"87", x"89", x"87", x"87", x"89", x"8a", x"88", x"84", x"83", x"84", x"86", x"88", x"88", 
        x"86", x"86", x"86", x"85", x"85", x"85", x"85", x"85", x"85", x"86", x"86", x"86", x"86", x"85", x"85", 
        x"85", x"84", x"83", x"82", x"85", x"85", x"84", x"83", x"83", x"85", x"86", x"84", x"83", x"83", x"84", 
        x"84", x"84", x"85", x"83", x"83", x"84", x"85", x"85", x"84", x"83", x"84", x"85", x"85", x"85", x"85", 
        x"84", x"84", x"83", x"82", x"83", x"84", x"85", x"85", x"85", x"84", x"85", x"85", x"85", x"84", x"84", 
        x"85", x"85", x"86", x"84", x"83", x"82", x"83", x"83", x"83", x"83", x"84", x"84", x"83", x"83", x"82", 
        x"82", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"81", x"81", x"81", x"82", x"82", x"82", 
        x"82", x"83", x"83", x"83", x"83", x"83", x"82", x"81", x"80", x"80", x"81", x"81", x"81", x"81", x"82", 
        x"81", x"81", x"82", x"83", x"83", x"83", x"83", x"82", x"81", x"82", x"81", x"81", x"81", x"81", x"80", 
        x"7f", x"81", x"83", x"81", x"80", x"80", x"80", x"7f", x"81", x"81", x"82", x"7f", x"7c", x"7e", x"76", 
        x"77", x"81", x"8d", x"95", x"9a", x"a3", x"b1", x"c1", x"cd", x"d6", x"d9", x"d2", x"cf", x"d0", x"d0", 
        x"7e", x"80", x"80", x"80", x"7e", x"7e", x"7e", x"7c", x"7c", x"7e", x"7d", x"7e", x"80", x"7f", x"81", 
        x"80", x"7e", x"7d", x"7b", x"7c", x"7c", x"7c", x"7f", x"7f", x"7f", x"80", x"80", x"80", x"80", x"7e", 
        x"7e", x"7d", x"7d", x"7e", x"7e", x"7e", x"7d", x"7d", x"7f", x"7e", x"7f", x"7d", x"7d", x"7e", x"7f", 
        x"7f", x"7e", x"7f", x"81", x"7f", x"7e", x"7e", x"7f", x"7f", x"7e", x"7e", x"7f", x"7f", x"80", x"7f", 
        x"7f", x"7f", x"7f", x"7f", x"7d", x"7d", x"80", x"80", x"7f", x"7f", x"82", x"82", x"80", x"80", x"81", 
        x"82", x"82", x"81", x"81", x"7f", x"7f", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", x"80", x"80", x"81", 
        x"80", x"81", x"82", x"82", x"82", x"81", x"81", x"81", x"81", x"80", x"80", x"7f", x"80", x"81", x"7f", 
        x"81", x"83", x"82", x"83", x"84", x"82", x"80", x"83", x"83", x"83", x"86", x"7e", x"73", x"7e", x"b1", 
        x"d2", x"d4", x"cd", x"cf", x"d0", x"d2", x"d0", x"d2", x"d4", x"d5", x"be", x"7a", x"32", x"1d", x"1c", 
        x"1b", x"1f", x"1c", x"19", x"1a", x"1a", x"18", x"16", x"16", x"18", x"1c", x"1c", x"16", x"12", x"0b", 
        x"22", x"aa", x"dc", x"d2", x"d1", x"d1", x"d5", x"d9", x"ce", x"cd", x"cf", x"d1", x"d1", x"d0", x"d0", 
        x"d1", x"d1", x"d2", x"d2", x"d0", x"ce", x"d0", x"d1", x"cf", x"cf", x"d0", x"d0", x"cf", x"d0", x"d1", 
        x"d0", x"d1", x"d2", x"d1", x"d0", x"d0", x"cf", x"d1", x"d0", x"cf", x"cf", x"d0", x"d2", x"d4", x"d3", 
        x"d1", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"dc", x"d1", x"d2", x"d3", x"d2", x"d3", x"cf", 
        x"d9", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"ef", x"f1", 
        x"f2", x"ef", x"ef", x"ef", x"f0", x"f0", x"ec", x"ee", x"f1", x"eb", x"e6", x"d3", x"b8", x"a3", x"8a", 
        x"77", x"70", x"a3", x"e2", x"f1", x"f1", x"b7", x"61", x"6a", x"7d", x"95", x"bc", x"eb", x"f7", x"e8", 
        x"9f", x"91", x"e6", x"f0", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"ee", x"ef", x"f2", x"f3", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ea", x"da", x"c6", x"ba", x"ba", 
        x"c9", x"dd", x"e8", x"ef", x"f4", x"f3", x"f1", x"ef", x"f0", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ed", x"ed", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"ef", x"ef", x"ef", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f0", x"eb", x"e5", x"e3", x"e2", x"e0", x"d0", x"af", x"8d", x"7e", x"7d", x"84", x"8a", 
        x"8b", x"87", x"88", x"88", x"89", x"88", x"89", x"88", x"87", x"85", x"85", x"87", x"87", x"87", x"88", 
        x"88", x"88", x"89", x"88", x"89", x"8a", x"8b", x"89", x"88", x"86", x"85", x"86", x"86", x"86", x"87", 
        x"85", x"85", x"87", x"89", x"87", x"85", x"86", x"88", x"87", x"86", x"86", x"87", x"86", x"87", x"86", 
        x"86", x"88", x"88", x"87", x"88", x"87", x"86", x"85", x"85", x"85", x"84", x"85", x"84", x"84", x"86", 
        x"85", x"83", x"84", x"83", x"84", x"85", x"84", x"83", x"84", x"84", x"85", x"84", x"84", x"84", x"85", 
        x"85", x"85", x"85", x"84", x"84", x"85", x"86", x"86", x"85", x"84", x"83", x"83", x"83", x"83", x"83", 
        x"83", x"84", x"83", x"82", x"83", x"84", x"85", x"85", x"85", x"85", x"84", x"85", x"86", x"86", x"86", 
        x"85", x"84", x"85", x"85", x"84", x"83", x"83", x"82", x"82", x"82", x"83", x"83", x"84", x"84", x"84", 
        x"84", x"84", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"81", x"81", x"81", x"82", x"82", x"82", 
        x"83", x"84", x"82", x"82", x"83", x"82", x"81", x"82", x"82", x"81", x"82", x"82", x"82", x"82", x"82", 
        x"80", x"7f", x"80", x"80", x"81", x"82", x"83", x"82", x"82", x"83", x"81", x"81", x"82", x"82", x"80", 
        x"7f", x"80", x"81", x"81", x"81", x"81", x"81", x"81", x"7e", x"7b", x"7b", x"7a", x"7c", x"87", x"92", 
        x"96", x"9f", x"ac", x"b8", x"c4", x"cf", x"d6", x"d5", x"cf", x"cf", x"d4", x"d3", x"d3", x"d2", x"d1", 
        x"7f", x"80", x"81", x"80", x"7e", x"7d", x"7d", x"7c", x"7e", x"7f", x"7e", x"7f", x"81", x"7f", x"7f", 
        x"7e", x"7d", x"7e", x"7c", x"7e", x"7d", x"7d", x"80", x"7f", x"7f", x"7e", x"7d", x"7d", x"7c", x"7d", 
        x"7e", x"7d", x"7d", x"80", x"82", x"80", x"7e", x"7d", x"80", x"7e", x"7f", x"7d", x"7e", x"7e", x"80", 
        x"80", x"7f", x"80", x"82", x"81", x"81", x"80", x"7e", x"7d", x"7d", x"7f", x"81", x"80", x"80", x"7f", 
        x"7f", x"80", x"80", x"80", x"7f", x"7f", x"81", x"7f", x"7f", x"80", x"83", x"81", x"7e", x"7e", x"80", 
        x"80", x"81", x"81", x"80", x"80", x"7f", x"7e", x"7d", x"7d", x"7f", x"80", x"81", x"80", x"81", x"81", 
        x"80", x"81", x"82", x"83", x"82", x"81", x"81", x"81", x"81", x"80", x"80", x"80", x"80", x"83", x"82", 
        x"83", x"85", x"82", x"82", x"83", x"81", x"81", x"84", x"87", x"83", x"75", x"6f", x"98", x"cc", x"d8", 
        x"d6", x"d2", x"d0", x"d1", x"d4", x"d4", x"d0", x"d6", x"d1", x"98", x"4d", x"1e", x"1a", x"1c", x"1d", 
        x"1c", x"1c", x"19", x"15", x"18", x"19", x"17", x"19", x"1b", x"18", x"1a", x"16", x"0c", x"08", x"03", 
        x"21", x"aa", x"dd", x"d3", x"d3", x"d2", x"d6", x"d9", x"d1", x"d0", x"d1", x"d1", x"d1", x"cf", x"ce", 
        x"cf", x"d0", x"d2", x"d3", x"d0", x"ce", x"ce", x"cf", x"ce", x"ce", x"d0", x"d1", x"d0", x"d1", x"d3", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d1", x"d1", x"d1", x"d2", x"d3", x"d4", x"d2", 
        x"d1", x"d1", x"d0", x"cf", x"cf", x"cf", x"cf", x"d0", x"dc", x"d2", x"d3", x"d3", x"d2", x"d3", x"cf", 
        x"d9", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"ee", x"f1", x"ef", x"f1", 
        x"f0", x"ee", x"ee", x"f0", x"ef", x"ed", x"ef", x"ee", x"ef", x"f0", x"ee", x"f1", x"f1", x"ec", x"d5", 
        x"b1", x"96", x"99", x"b1", x"c8", x"ce", x"9e", x"61", x"62", x"5e", x"5b", x"75", x"c9", x"f6", x"f3", 
        x"be", x"9a", x"e5", x"f1", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"f0", x"f1", x"f1", x"f1", 
        x"f2", x"f1", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"f1", x"f3", x"ea", x"d3", 
        x"c0", x"ba", x"be", x"d2", x"e2", x"ed", x"f4", x"f3", x"ee", x"ef", x"f1", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ed", x"ed", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f2", x"f0", x"ef", x"ef", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"ef", x"ee", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"f2", x"f2", x"f0", x"f2", x"f4", x"f0", x"e4", x"dd", x"e0", x"e6", x"dc", x"ba", x"91", x"79", x"7b", 
        x"84", x"89", x"8a", x"89", x"89", x"89", x"89", x"89", x"88", x"86", x"86", x"88", x"87", x"86", x"89", 
        x"88", x"87", x"88", x"88", x"87", x"87", x"87", x"88", x"86", x"87", x"87", x"87", x"88", x"86", x"87", 
        x"87", x"86", x"88", x"89", x"86", x"84", x"85", x"85", x"86", x"87", x"87", x"88", x"88", x"89", x"88", 
        x"86", x"88", x"87", x"85", x"87", x"87", x"86", x"85", x"85", x"85", x"84", x"84", x"82", x"83", x"87", 
        x"84", x"81", x"84", x"84", x"84", x"85", x"85", x"85", x"85", x"85", x"85", x"85", x"86", x"86", x"85", 
        x"85", x"84", x"83", x"85", x"86", x"86", x"84", x"84", x"84", x"84", x"82", x"81", x"83", x"85", x"86", 
        x"86", x"84", x"84", x"83", x"83", x"84", x"84", x"84", x"85", x"85", x"84", x"84", x"85", x"85", x"85", 
        x"84", x"84", x"84", x"84", x"85", x"83", x"82", x"81", x"81", x"81", x"81", x"82", x"82", x"83", x"84", 
        x"84", x"83", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"83", x"83", x"83", 
        x"84", x"85", x"80", x"80", x"82", x"81", x"80", x"82", x"83", x"83", x"83", x"82", x"82", x"82", x"82", 
        x"82", x"81", x"80", x"80", x"81", x"82", x"83", x"83", x"83", x"84", x"81", x"81", x"83", x"83", x"81", 
        x"81", x"82", x"82", x"82", x"81", x"7e", x"7b", x"7a", x"7b", x"80", x"89", x"8f", x"9a", x"ab", x"b5", 
        x"bb", x"c3", x"cd", x"d6", x"d8", x"d4", x"d1", x"d2", x"cf", x"cf", x"d1", x"d0", x"d0", x"d0", x"d1", 
        x"7e", x"7e", x"81", x"82", x"80", x"80", x"81", x"7f", x"80", x"80", x"7f", x"7f", x"7f", x"7d", x"7d", 
        x"7c", x"7c", x"7e", x"7e", x"7f", x"7f", x"7d", x"7e", x"7e", x"7d", x"7c", x"7d", x"7d", x"7a", x"7c", 
        x"7d", x"7d", x"7d", x"7f", x"82", x"81", x"7e", x"7e", x"7f", x"7d", x"7f", x"80", x"81", x"7f", x"7f", 
        x"7f", x"7f", x"7f", x"80", x"82", x"81", x"7f", x"7f", x"7f", x"7f", x"80", x"80", x"80", x"80", x"7f", 
        x"7f", x"80", x"80", x"80", x"80", x"7e", x"7f", x"80", x"7f", x"80", x"82", x"80", x"80", x"7e", x"7e", 
        x"7f", x"80", x"80", x"7f", x"81", x"7f", x"7d", x"7c", x"7c", x"7e", x"7f", x"81", x"7f", x"80", x"82", 
        x"80", x"82", x"84", x"82", x"80", x"80", x"7f", x"7f", x"80", x"81", x"81", x"81", x"83", x"84", x"84", 
        x"84", x"87", x"82", x"81", x"80", x"80", x"85", x"85", x"76", x"6e", x"88", x"ba", x"d5", x"d7", x"d3", 
        x"d1", x"d0", x"ce", x"ce", x"d1", x"d7", x"d3", x"b0", x"5e", x"28", x"17", x"1b", x"1c", x"1a", x"1a", 
        x"1b", x"1b", x"1c", x"1c", x"17", x"17", x"18", x"18", x"18", x"16", x"0f", x"09", x"03", x"04", x"03", 
        x"21", x"ab", x"de", x"d3", x"d4", x"d4", x"d7", x"d8", x"d1", x"d1", x"d2", x"d1", x"d0", x"d0", x"cf", 
        x"d0", x"d1", x"d1", x"d1", x"d0", x"cf", x"d0", x"d1", x"d0", x"ce", x"cf", x"d0", x"d0", x"d1", x"d1", 
        x"d1", x"d1", x"d0", x"d1", x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", x"d1", x"d2", x"d2", x"d3", x"d4", 
        x"d4", x"d4", x"d2", x"d0", x"cf", x"d0", x"ce", x"ce", x"dc", x"d2", x"d3", x"d4", x"d3", x"d4", x"d0", 
        x"d8", x"ee", x"f0", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ed", x"ee", 
        x"f0", x"ed", x"ed", x"f0", x"ee", x"ed", x"f1", x"f0", x"f0", x"f0", x"ee", x"f0", x"f0", x"f1", x"f4", 
        x"f3", x"ec", x"da", x"be", x"ab", x"a0", x"86", x"6c", x"67", x"68", x"64", x"61", x"a7", x"ee", x"f5", 
        x"d7", x"af", x"e4", x"f2", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", 
        x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ee", x"ef", x"f0", x"f1", x"f2", x"f2", 
        x"f1", x"f0", x"ef", x"f0", x"f2", x"f2", x"f0", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"f2", x"f5", 
        x"f2", x"e6", x"cf", x"c2", x"bf", x"c4", x"d4", x"e5", x"f1", x"f3", x"f2", x"f0", x"f0", x"f0", x"f1", 
        x"f2", x"f2", x"f1", x"ef", x"f0", x"f1", x"ef", x"ee", x"f0", x"ef", x"ef", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f2", x"f3", x"f0", x"ea", x"e1", x"df", x"e3", x"de", x"c6", x"a5", 
        x"89", x"77", x"7a", x"86", x"8a", x"87", x"86", x"88", x"89", x"88", x"8a", x"8c", x"89", x"87", x"8a", 
        x"88", x"86", x"87", x"89", x"88", x"85", x"88", x"89", x"87", x"88", x"88", x"85", x"87", x"87", x"88", 
        x"89", x"88", x"88", x"88", x"86", x"86", x"85", x"86", x"87", x"88", x"87", x"86", x"85", x"87", x"88", 
        x"86", x"88", x"89", x"88", x"87", x"85", x"86", x"85", x"85", x"87", x"87", x"85", x"84", x"83", x"87", 
        x"85", x"82", x"85", x"84", x"85", x"85", x"86", x"86", x"86", x"85", x"84", x"85", x"85", x"85", x"85", 
        x"85", x"85", x"83", x"85", x"85", x"85", x"85", x"83", x"85", x"86", x"83", x"82", x"85", x"87", x"87", 
        x"86", x"85", x"85", x"85", x"83", x"85", x"86", x"84", x"83", x"84", x"83", x"84", x"85", x"84", x"84", 
        x"84", x"86", x"86", x"86", x"85", x"83", x"81", x"81", x"82", x"83", x"82", x"82", x"82", x"83", x"84", 
        x"84", x"82", x"81", x"82", x"82", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"82", 
        x"83", x"84", x"82", x"80", x"82", x"82", x"80", x"83", x"85", x"83", x"83", x"82", x"81", x"80", x"82", 
        x"84", x"82", x"81", x"82", x"82", x"83", x"84", x"83", x"82", x"84", x"84", x"83", x"83", x"83", x"84", 
        x"84", x"81", x"7f", x"7e", x"7e", x"80", x"83", x"8c", x"94", x"9f", x"af", x"bb", x"c3", x"c9", x"d2", 
        x"d5", x"d5", x"d3", x"d2", x"d3", x"d2", x"d3", x"d3", x"d2", x"d0", x"cf", x"d0", x"d2", x"d1", x"d2", 
        x"84", x"80", x"83", x"83", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", x"7e", x"7d", x"7c", x"7b", x"7d", 
        x"7e", x"7e", x"7f", x"7f", x"7f", x"7f", x"7d", x"7e", x"7f", x"7e", x"7e", x"7f", x"7e", x"7c", x"7d", 
        x"7e", x"7e", x"7d", x"7e", x"7f", x"80", x"7e", x"7f", x"7e", x"7d", x"7d", x"80", x"82", x"7e", x"7d", 
        x"7e", x"7f", x"7f", x"80", x"81", x"80", x"80", x"80", x"7f", x"7e", x"7e", x"7f", x"80", x"80", x"80", 
        x"80", x"80", x"80", x"80", x"7f", x"7c", x"7e", x"82", x"7f", x"7e", x"81", x"80", x"81", x"7f", x"7f", 
        x"80", x"82", x"80", x"7d", x"7f", x"7d", x"7c", x"7c", x"7e", x"7f", x"80", x"83", x"80", x"81", x"82", 
        x"80", x"82", x"83", x"82", x"81", x"81", x"81", x"80", x"80", x"83", x"82", x"82", x"83", x"83", x"83", 
        x"7f", x"85", x"82", x"81", x"85", x"85", x"82", x"71", x"79", x"9e", x"cb", x"d8", x"d2", x"cf", x"d2", 
        x"d1", x"cf", x"d1", x"d2", x"d9", x"c5", x"81", x"41", x"1f", x"1f", x"1e", x"1c", x"1c", x"1a", x"17", 
        x"18", x"19", x"18", x"18", x"17", x"18", x"17", x"15", x"13", x"0d", x"05", x"02", x"03", x"06", x"07", 
        x"21", x"ab", x"de", x"d2", x"d5", x"d5", x"d8", x"d8", x"cf", x"d0", x"d1", x"cf", x"cf", x"d1", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", x"d1", x"d2", x"d1", x"cf", x"ce", x"cf", x"cf", x"cf", x"d0", 
        x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d0", x"d1", x"d2", x"d2", x"d3", 
        x"d4", x"d3", x"d1", x"cf", x"cf", x"d0", x"cd", x"ce", x"dc", x"d2", x"d3", x"d4", x"d4", x"d4", x"d1", 
        x"d7", x"ec", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", 
        x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ed", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f0", x"f0", x"f1", x"f0", x"e7", x"d5", x"bb", x"a1", x"8f", x"92", x"88", x"6c", x"90", x"e0", x"f5", 
        x"e8", x"c6", x"e3", x"f1", x"ee", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f2", x"f2", x"e9", x"db", x"cb", x"c2", x"c3", x"ce", x"dc", x"e9", x"f0", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f0", x"ed", x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f3", x"f1", x"e8", x"de", x"da", x"dc", x"d6", 
        x"c9", x"ac", x"8f", x"7d", x"7a", x"84", x"89", x"8a", x"8a", x"8b", x"8a", x"89", x"89", x"8b", x"8d", 
        x"8b", x"88", x"89", x"8b", x"8a", x"88", x"89", x"87", x"87", x"87", x"87", x"88", x"8a", x"88", x"88", 
        x"89", x"89", x"87", x"87", x"87", x"87", x"86", x"86", x"89", x"89", x"88", x"87", x"85", x"87", x"87", 
        x"86", x"86", x"88", x"87", x"85", x"86", x"88", x"85", x"84", x"87", x"87", x"84", x"86", x"84", x"87", 
        x"85", x"84", x"87", x"85", x"86", x"86", x"86", x"86", x"85", x"85", x"84", x"84", x"84", x"84", x"84", 
        x"85", x"85", x"83", x"85", x"84", x"85", x"86", x"84", x"85", x"85", x"83", x"83", x"85", x"85", x"84", 
        x"83", x"84", x"85", x"85", x"82", x"83", x"85", x"83", x"83", x"84", x"82", x"84", x"86", x"85", x"84", 
        x"84", x"86", x"87", x"86", x"84", x"83", x"83", x"85", x"87", x"86", x"83", x"82", x"82", x"83", x"85", 
        x"85", x"84", x"83", x"83", x"84", x"84", x"83", x"83", x"83", x"84", x"84", x"83", x"82", x"81", x"81", 
        x"81", x"83", x"83", x"81", x"82", x"83", x"81", x"83", x"83", x"7f", x"81", x"81", x"82", x"80", x"83", 
        x"83", x"80", x"80", x"85", x"88", x"85", x"83", x"82", x"82", x"83", x"85", x"84", x"81", x"82", x"81", 
        x"7d", x"7e", x"83", x"88", x"8f", x"96", x"a1", x"af", x"bb", x"c4", x"ca", x"d2", x"d5", x"d3", x"d1", 
        x"d0", x"d2", x"d3", x"d1", x"d0", x"d1", x"d2", x"d0", x"d2", x"d1", x"cf", x"d1", x"d1", x"d1", x"d2", 
        x"84", x"80", x"80", x"80", x"7d", x"7e", x"7e", x"7e", x"7f", x"7f", x"7e", x"7d", x"7d", x"7c", x"7d", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"80", x"80", x"7f", x"7e", x"7e", x"7d", x"7d", x"7d", 
        x"7f", x"7f", x"7e", x"7e", x"7f", x"80", x"7e", x"7f", x"7e", x"7d", x"7c", x"7d", x"7e", x"7c", x"7e", 
        x"7f", x"7e", x"80", x"82", x"80", x"7f", x"80", x"80", x"7f", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"80", x"82", x"7f", x"7d", x"7e", x"7d", x"80", x"7e", x"7e", 
        x"7f", x"80", x"7e", x"7c", x"7f", x"7e", x"7d", x"7d", x"7e", x"80", x"81", x"80", x"7f", x"81", x"81", 
        x"80", x"83", x"84", x"82", x"82", x"83", x"83", x"82", x"82", x"83", x"83", x"83", x"82", x"82", x"85", 
        x"82", x"84", x"82", x"84", x"8a", x"78", x"69", x"8c", x"be", x"d5", x"d3", x"d3", x"d1", x"d2", x"cf", 
        x"ce", x"d1", x"dd", x"d9", x"a7", x"52", x"25", x"1b", x"21", x"1d", x"1b", x"1c", x"1d", x"1b", x"17", 
        x"16", x"17", x"17", x"18", x"18", x"18", x"14", x"0e", x"08", x"03", x"01", x"03", x"06", x"07", x"08", 
        x"20", x"a9", x"e0", x"d5", x"d5", x"d3", x"d6", x"d8", x"cf", x"d0", x"d1", x"cf", x"cf", x"d1", x"d1", 
        x"d1", x"d1", x"d1", x"d2", x"d1", x"d0", x"cf", x"d0", x"d0", x"cf", x"ce", x"cf", x"cf", x"cf", x"cf", 
        x"d0", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", 
        x"d4", x"d2", x"d1", x"cf", x"cf", x"d0", x"ce", x"cf", x"dc", x"d2", x"d3", x"d4", x"d3", x"d4", x"d2", 
        x"d6", x"ec", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ee", 
        x"ee", x"ed", x"ee", x"ee", x"ef", x"f0", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"ea", x"da", x"d7", x"c2", x"97", x"8b", x"b2", x"d4", 
        x"e9", x"e1", x"e9", x"f0", x"ec", x"ee", x"ed", x"ed", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f3", x"f2", 
        x"ee", x"ec", x"ef", x"f0", x"f1", x"ef", x"e7", x"d8", x"c8", x"be", x"bf", x"ce", x"e9", x"f2", x"f6", 
        x"f2", x"f0", x"f1", x"ef", x"ef", x"f2", x"f2", x"ec", x"ed", x"ef", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"f2", x"f3", x"ef", x"e7", x"dd", x"cf", 
        x"cb", x"d4", x"d6", x"bc", x"91", x"7b", x"78", x"84", x"8d", x"8c", x"89", x"8b", x"8c", x"8c", x"8d", 
        x"89", x"88", x"89", x"88", x"88", x"88", x"87", x"87", x"87", x"87", x"88", x"8b", x"8a", x"88", x"88", 
        x"88", x"87", x"86", x"86", x"87", x"88", x"88", x"87", x"86", x"86", x"87", x"87", x"85", x"86", x"87", 
        x"86", x"86", x"88", x"89", x"86", x"87", x"89", x"86", x"85", x"88", x"88", x"85", x"85", x"84", x"86", 
        x"85", x"84", x"86", x"84", x"85", x"86", x"86", x"85", x"83", x"84", x"85", x"86", x"85", x"84", x"84", 
        x"85", x"86", x"85", x"85", x"84", x"85", x"85", x"83", x"83", x"83", x"81", x"83", x"84", x"84", x"84", 
        x"83", x"84", x"85", x"85", x"83", x"83", x"84", x"84", x"85", x"86", x"84", x"85", x"86", x"85", x"84", 
        x"84", x"84", x"86", x"86", x"86", x"85", x"85", x"86", x"86", x"87", x"86", x"84", x"84", x"85", x"85", 
        x"85", x"84", x"84", x"83", x"82", x"82", x"81", x"81", x"82", x"83", x"83", x"83", x"82", x"82", x"82", 
        x"82", x"83", x"84", x"82", x"82", x"83", x"82", x"84", x"83", x"81", x"83", x"84", x"83", x"81", x"82", 
        x"82", x"81", x"83", x"84", x"82", x"80", x"82", x"82", x"81", x"82", x"84", x"81", x"7c", x"78", x"7f", 
        x"8a", x"8f", x"97", x"a4", x"b2", x"c0", x"cb", x"d1", x"d6", x"d7", x"d3", x"d1", x"d1", x"d1", x"d1", 
        x"d1", x"d2", x"d4", x"d2", x"d1", x"d1", x"d3", x"d2", x"d2", x"d2", x"d0", x"d2", x"d1", x"d2", x"d1", 
        x"82", x"7f", x"7f", x"7f", x"80", x"80", x"7f", x"7f", x"7f", x"7f", x"7e", x"7e", x"7e", x"7d", x"7d", 
        x"7e", x"7e", x"7e", x"7e", x"7e", x"7e", x"7f", x"80", x"7e", x"7f", x"7f", x"7e", x"7e", x"7f", x"7d", 
        x"7f", x"80", x"80", x"80", x"80", x"80", x"7f", x"7f", x"7e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7e", 
        x"7f", x"7e", x"81", x"82", x"80", x"80", x"81", x"81", x"80", x"7e", x"7e", x"7e", x"7f", x"7f", x"7f", 
        x"7f", x"7f", x"7f", x"7f", x"7e", x"7e", x"7f", x"80", x"7f", x"7f", x"80", x"7e", x"7d", x"7d", x"7e", 
        x"80", x"82", x"81", x"7f", x"82", x"81", x"80", x"80", x"80", x"81", x"81", x"81", x"82", x"82", x"80", 
        x"80", x"81", x"81", x"7f", x"80", x"81", x"82", x"82", x"83", x"83", x"85", x"85", x"80", x"81", x"83", 
        x"81", x"85", x"8a", x"84", x"6c", x"7d", x"ac", x"ce", x"d6", x"d1", x"d1", x"d0", x"d0", x"d1", x"d0", 
        x"d5", x"db", x"b6", x"6f", x"34", x"20", x"1f", x"1d", x"1e", x"1b", x"1b", x"1d", x"1e", x"1c", x"1a", 
        x"1a", x"19", x"18", x"1b", x"18", x"11", x"09", x"03", x"02", x"03", x"04", x"08", x"09", x"09", x"08", 
        x"21", x"a9", x"e0", x"d5", x"d4", x"d1", x"d6", x"d8", x"cf", x"d0", x"d1", x"cf", x"cf", x"d1", x"d1", 
        x"d1", x"d1", x"d2", x"d1", x"d1", x"cf", x"ce", x"cf", x"d0", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", 
        x"d0", x"d0", x"d1", x"d1", x"d2", x"d3", x"d3", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", 
        x"d3", x"d2", x"d1", x"d0", x"d0", x"d0", x"cf", x"d0", x"dd", x"d3", x"d3", x"d3", x"d3", x"d4", x"d2", 
        x"d6", x"ec", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", 
        x"ee", x"ed", x"ee", x"ee", x"ef", x"f0", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f0", x"f0", 
        x"f0", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f0", x"ee", x"ef", x"f1", x"ef", x"ec", x"ef", x"f3", x"f3", x"e8", x"e1", x"d5", x"c0", x"ad", 
        x"ac", x"b3", x"cc", x"e0", x"ec", x"f0", x"ee", x"ee", x"f2", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ed", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f0", x"ee", x"ee", x"ef", x"f2", x"f3", x"f1", x"ee", x"e7", x"da", x"c9", x"bd", x"c3", x"d4", 
        x"ea", x"f3", x"f3", x"f1", x"f2", x"f2", x"f0", x"ee", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f0", x"ef", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f1", x"ef", x"ee", x"ee", x"e8", 
        x"e3", x"d6", x"cf", x"d5", x"d8", x"c4", x"a0", x"82", x"7d", x"80", x"87", x"89", x"8a", x"89", x"88", 
        x"8c", x"8f", x"8e", x"8a", x"88", x"8a", x"88", x"89", x"88", x"88", x"8a", x"8c", x"8a", x"89", x"8a", 
        x"8a", x"88", x"87", x"87", x"89", x"89", x"8a", x"89", x"86", x"85", x"86", x"87", x"87", x"88", x"88", 
        x"88", x"88", x"89", x"88", x"87", x"87", x"89", x"87", x"86", x"88", x"88", x"86", x"85", x"85", x"86", 
        x"86", x"85", x"86", x"85", x"86", x"86", x"85", x"84", x"84", x"85", x"85", x"87", x"85", x"85", x"85", 
        x"86", x"86", x"86", x"84", x"83", x"85", x"85", x"84", x"85", x"85", x"83", x"83", x"83", x"83", x"83", 
        x"84", x"87", x"87", x"83", x"83", x"85", x"86", x"86", x"86", x"86", x"85", x"85", x"85", x"85", x"85", 
        x"84", x"83", x"80", x"81", x"83", x"85", x"85", x"85", x"85", x"84", x"83", x"83", x"84", x"85", x"86", 
        x"85", x"84", x"82", x"82", x"82", x"82", x"82", x"83", x"83", x"83", x"83", x"83", x"83", x"84", x"84", 
        x"84", x"83", x"83", x"83", x"84", x"84", x"83", x"83", x"85", x"83", x"84", x"84", x"83", x"81", x"84", 
        x"86", x"85", x"84", x"84", x"82", x"81", x"83", x"85", x"82", x"7d", x"7c", x"82", x"8b", x"95", x"9c", 
        x"a7", x"b5", x"c3", x"ce", x"d4", x"d5", x"d3", x"d2", x"d1", x"d3", x"d2", x"d1", x"d1", x"d2", x"d3", 
        x"d3", x"d4", x"d4", x"d3", x"d2", x"d2", x"d3", x"d2", x"d3", x"d3", x"d1", x"d2", x"d2", x"d2", x"d3", 
        x"81", x"81", x"80", x"81", x"82", x"82", x"80", x"7f", x"7f", x"7f", x"7e", x"7e", x"7e", x"7e", x"7e", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"80", x"80", x"7e", x"7f", x"7f", x"7e", x"7f", x"7f", x"7e", 
        x"7f", x"81", x"80", x"80", x"80", x"80", x"80", x"7e", x"7e", x"7e", x"7e", x"7f", x"80", x"81", x"7f", 
        x"7d", x"7f", x"81", x"80", x"80", x"82", x"83", x"82", x"82", x"81", x"80", x"7f", x"7f", x"7f", x"7f", 
        x"7f", x"7f", x"7f", x"7f", x"7e", x"7d", x"7e", x"7f", x"80", x"81", x"81", x"81", x"7e", x"7e", x"7f", 
        x"81", x"82", x"82", x"81", x"82", x"82", x"82", x"81", x"80", x"81", x"82", x"7f", x"80", x"81", x"80", 
        x"82", x"83", x"83", x"84", x"84", x"83", x"83", x"83", x"83", x"83", x"85", x"86", x"84", x"81", x"83", 
        x"87", x"84", x"76", x"6c", x"97", x"c1", x"d2", x"d2", x"cd", x"cf", x"d0", x"d1", x"d3", x"d4", x"d8", 
        x"cc", x"96", x"44", x"26", x"20", x"21", x"1f", x"21", x"1f", x"1c", x"1c", x"1c", x"1b", x"1a", x"1a", 
        x"1a", x"19", x"17", x"14", x"0d", x"05", x"02", x"04", x"06", x"08", x"08", x"09", x"09", x"08", x"08", 
        x"21", x"ab", x"df", x"d2", x"d3", x"d2", x"d6", x"d7", x"cf", x"d0", x"d1", x"cf", x"cf", x"d1", x"d1", 
        x"d2", x"d2", x"d1", x"d0", x"cf", x"cf", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"cf", x"cf", x"d0", 
        x"d0", x"d0", x"d0", x"d1", x"d2", x"d3", x"d3", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d4", 
        x"d3", x"d1", x"d1", x"d1", x"d0", x"d0", x"cf", x"d0", x"de", x"d3", x"d3", x"d3", x"d3", x"d4", x"d2", 
        x"d6", x"ec", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"f0", x"f0", 
        x"f0", x"f0", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", x"eb", x"ee", x"eb", x"e6", x"e0", 
        x"d8", x"c4", x"af", x"ab", x"b2", x"cd", x"e4", x"ed", x"f0", x"ef", x"f0", x"f0", x"ef", x"ee", x"ed", 
        x"ee", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ed", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f2", x"f4", x"f0", x"ee", 
        x"f0", x"f1", x"f0", x"f0", x"f2", x"f3", x"f0", x"ec", x"ee", x"f3", x"f1", x"eb", x"e2", x"d5", x"c3", 
        x"bd", x"ca", x"df", x"ee", x"ef", x"f1", x"ef", x"ea", x"ec", x"ee", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f2", x"ee", x"e7", x"db", x"d1", x"d5", x"d6", x"c8", x"a8", x"8a", x"7e", x"80", x"87", x"8a", x"89", 
        x"8a", x"89", x"89", x"8a", x"8a", x"89", x"8a", x"8c", x"8a", x"89", x"8a", x"8a", x"88", x"89", x"8a", 
        x"8a", x"88", x"87", x"88", x"89", x"86", x"87", x"88", x"87", x"86", x"88", x"89", x"88", x"87", x"87", 
        x"87", x"87", x"86", x"86", x"86", x"87", x"88", x"86", x"86", x"87", x"87", x"86", x"85", x"86", x"86", 
        x"86", x"86", x"85", x"86", x"89", x"86", x"83", x"84", x"86", x"86", x"84", x"86", x"86", x"85", x"86", 
        x"87", x"87", x"85", x"85", x"86", x"86", x"87", x"86", x"86", x"86", x"86", x"86", x"85", x"85", x"85", 
        x"86", x"86", x"85", x"83", x"84", x"86", x"86", x"87", x"87", x"86", x"86", x"84", x"84", x"85", x"86", 
        x"86", x"84", x"85", x"86", x"88", x"88", x"87", x"85", x"83", x"82", x"82", x"83", x"83", x"84", x"84", 
        x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"84", x"84", x"83", x"83", x"83", x"84", x"84", x"85", 
        x"85", x"83", x"83", x"85", x"85", x"84", x"83", x"83", x"83", x"80", x"82", x"82", x"82", x"80", x"83", 
        x"84", x"83", x"83", x"84", x"83", x"80", x"7b", x"7b", x"84", x"8e", x"95", x"9b", x"a6", x"b4", x"c3", 
        x"cf", x"d6", x"d8", x"d8", x"d8", x"d5", x"d2", x"d2", x"ce", x"cf", x"d2", x"d2", x"d2", x"d3", x"d3", 
        x"d3", x"d4", x"d4", x"d4", x"d3", x"d2", x"d4", x"d2", x"d4", x"d3", x"d1", x"d3", x"d2", x"d2", x"d2", 
        x"7f", x"82", x"81", x"82", x"83", x"82", x"80", x"80", x"7f", x"7e", x"7e", x"7e", x"7f", x"7f", x"80", 
        x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"7f", x"7f", x"7f", x"80", x"7f", x"80", x"80", x"7e", 
        x"7f", x"80", x"7f", x"7f", x"7f", x"80", x"80", x"7f", x"7e", x"7e", x"80", x"82", x"82", x"82", x"7f", 
        x"7e", x"7f", x"80", x"7f", x"81", x"83", x"84", x"82", x"82", x"82", x"82", x"80", x"7f", x"7f", x"7f", 
        x"7f", x"7f", x"7f", x"7f", x"7f", x"80", x"7f", x"7e", x"80", x"81", x"80", x"81", x"81", x"80", x"80", 
        x"80", x"80", x"80", x"80", x"81", x"82", x"82", x"82", x"81", x"81", x"82", x"82", x"84", x"82", x"81", 
        x"82", x"82", x"81", x"82", x"82", x"82", x"82", x"83", x"83", x"83", x"82", x"80", x"81", x"85", x"87", 
        x"83", x"6b", x"73", x"ad", x"d3", x"d6", x"d1", x"ce", x"cf", x"ce", x"d0", x"d5", x"d7", x"dc", x"b4", 
        x"6a", x"2c", x"1f", x"21", x"20", x"1b", x"1d", x"1f", x"1b", x"1a", x"1b", x"19", x"19", x"1b", x"1d", 
        x"1b", x"14", x"0d", x"06", x"02", x"01", x"04", x"08", x"08", x"08", x"07", x"07", x"08", x"07", x"08", 
        x"22", x"a9", x"dd", x"d1", x"d3", x"d3", x"d7", x"d7", x"cf", x"d0", x"d1", x"cf", x"cf", x"d1", x"d1", 
        x"d2", x"d2", x"d0", x"cf", x"cf", x"cf", x"d0", x"cf", x"cf", x"d0", x"d1", x"d0", x"d0", x"d0", x"d1", 
        x"d1", x"d0", x"d0", x"d0", x"d1", x"d3", x"d3", x"d2", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", 
        x"d2", x"d2", x"d2", x"d2", x"d0", x"cf", x"ce", x"d0", x"de", x"d3", x"d3", x"d4", x"d4", x"d4", x"d2", 
        x"d6", x"ec", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", 
        x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"e7", x"e9", x"f0", x"f2", x"ef", 
        x"ef", x"eb", x"e5", x"d9", x"c1", x"ab", x"a9", x"b8", x"d2", x"e5", x"ed", x"f2", x"f1", x"ef", x"f0", 
        x"f2", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f0", 
        x"f1", x"f1", x"ef", x"f1", x"f3", x"f2", x"f2", x"f3", x"f2", x"ee", x"f0", x"f2", x"ef", x"ed", x"e9", 
        x"dc", x"cd", x"c2", x"c4", x"d8", x"e6", x"f0", x"f1", x"f2", x"ef", x"ee", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f3", x"f0", x"ef", x"f1", x"f1", x"f1", x"ed", 
        x"f0", x"f1", x"ef", x"ef", x"e9", x"d9", x"ca", x"ce", x"da", x"d7", x"b3", x"87", x"77", x"7c", x"85", 
        x"8b", x"8e", x"8d", x"8c", x"8a", x"87", x"8b", x"8c", x"8c", x"8a", x"89", x"88", x"87", x"88", x"89", 
        x"89", x"87", x"86", x"86", x"87", x"85", x"86", x"87", x"87", x"87", x"88", x"88", x"88", x"87", x"87", 
        x"89", x"88", x"88", x"88", x"88", x"87", x"87", x"86", x"86", x"86", x"87", x"86", x"86", x"88", x"86", 
        x"87", x"88", x"86", x"87", x"89", x"87", x"85", x"85", x"88", x"87", x"85", x"85", x"86", x"86", x"87", 
        x"88", x"87", x"85", x"85", x"87", x"87", x"87", x"89", x"87", x"87", x"87", x"86", x"87", x"88", x"89", 
        x"88", x"85", x"84", x"85", x"86", x"85", x"84", x"87", x"88", x"87", x"86", x"84", x"84", x"86", x"87", 
        x"87", x"85", x"84", x"85", x"87", x"87", x"87", x"86", x"85", x"84", x"84", x"85", x"84", x"83", x"81", 
        x"81", x"83", x"86", x"85", x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"85", x"85", x"86", 
        x"85", x"84", x"84", x"86", x"86", x"85", x"85", x"83", x"82", x"82", x"86", x"86", x"86", x"82", x"82", 
        x"84", x"84", x"81", x"7d", x"7f", x"86", x"8d", x"94", x"9e", x"aa", x"b6", x"c4", x"d0", x"d7", x"d6", 
        x"d1", x"d4", x"d4", x"d3", x"d2", x"d2", x"d3", x"d4", x"d1", x"d3", x"d6", x"d6", x"d4", x"d3", x"d3", 
        x"d5", x"d4", x"d4", x"d4", x"d4", x"d3", x"d3", x"d2", x"d3", x"d3", x"d1", x"d3", x"d2", x"d2", x"d3", 
        x"81", x"85", x"82", x"80", x"81", x"80", x"7f", x"80", x"7f", x"7e", x"7e", x"7e", x"7f", x"80", x"81", 
        x"80", x"80", x"80", x"80", x"80", x"80", x"7f", x"7f", x"80", x"7f", x"80", x"81", x"81", x"7f", x"7f", 
        x"80", x"7f", x"7f", x"7f", x"7f", x"81", x"7f", x"7e", x"7e", x"80", x"81", x"81", x"80", x"80", x"81", 
        x"80", x"80", x"80", x"80", x"81", x"83", x"82", x"81", x"81", x"82", x"82", x"81", x"80", x"80", x"80", 
        x"80", x"80", x"80", x"80", x"80", x"82", x"80", x"7d", x"81", x"82", x"80", x"82", x"82", x"81", x"7f", 
        x"7e", x"7e", x"7f", x"80", x"7f", x"80", x"82", x"82", x"81", x"82", x"84", x"82", x"83", x"81", x"82", 
        x"85", x"83", x"85", x"82", x"7f", x"7f", x"81", x"83", x"84", x"82", x"81", x"7f", x"82", x"85", x"73", 
        x"6d", x"96", x"cd", x"d7", x"ce", x"d0", x"cc", x"ce", x"d1", x"cf", x"d2", x"da", x"c1", x"80", x"38", 
        x"1e", x"1b", x"1e", x"1e", x"1c", x"1d", x"1f", x"1d", x"1e", x"1c", x"1b", x"1a", x"1a", x"1b", x"1b", 
        x"13", x"09", x"02", x"02", x"02", x"05", x"08", x"08", x"07", x"06", x"05", x"06", x"08", x"09", x"09", 
        x"21", x"a4", x"dc", x"d4", x"d5", x"d3", x"d6", x"d7", x"cf", x"d0", x"d1", x"cf", x"cf", x"d1", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"cf", x"cf", x"d1", x"d2", x"d1", x"d1", x"d1", x"d2", 
        x"d2", x"d1", x"d0", x"d0", x"d1", x"d2", x"d3", x"d2", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", 
        x"d2", x"d2", x"d3", x"d2", x"d0", x"ce", x"ce", x"cf", x"dd", x"d3", x"d4", x"d5", x"d5", x"d5", x"d2", 
        x"d6", x"ec", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"f0", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"ef", x"ee", x"ee", x"ef", x"ef", x"ec", x"ee", x"ee", x"ed", x"f0", x"f1", x"ed", x"ef", 
        x"ef", x"ef", x"f0", x"ee", x"ef", x"ed", x"e3", x"c6", x"ad", x"a9", x"ba", x"d4", x"e2", x"eb", x"ee", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f1", x"f0", x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", 
        x"f3", x"f2", x"ef", x"f0", x"ef", x"f1", x"f2", x"f0", x"ef", x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", 
        x"f3", x"f0", x"e7", x"d5", x"c1", x"c1", x"c9", x"d8", x"e9", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f3", x"ef", 
        x"ef", x"ef", x"f1", x"ef", x"eb", x"ef", x"ed", x"e1", x"d0", x"ce", x"dd", x"dc", x"bb", x"93", x"7b", 
        x"7d", x"81", x"87", x"8a", x"8c", x"8b", x"8b", x"8a", x"8b", x"8b", x"89", x"88", x"88", x"87", x"88", 
        x"89", x"88", x"86", x"86", x"87", x"89", x"87", x"87", x"88", x"88", x"87", x"86", x"8a", x"8c", x"8a", 
        x"8b", x"89", x"86", x"86", x"88", x"87", x"87", x"87", x"87", x"87", x"87", x"87", x"87", x"89", x"86", 
        x"87", x"89", x"87", x"88", x"88", x"88", x"88", x"88", x"87", x"87", x"87", x"87", x"86", x"86", x"86", 
        x"87", x"87", x"86", x"85", x"87", x"86", x"86", x"88", x"87", x"86", x"87", x"86", x"86", x"87", x"87", 
        x"87", x"86", x"85", x"87", x"88", x"86", x"85", x"87", x"88", x"87", x"86", x"86", x"86", x"86", x"86", 
        x"85", x"84", x"86", x"86", x"86", x"86", x"85", x"85", x"84", x"84", x"85", x"87", x"86", x"84", x"83", 
        x"82", x"83", x"85", x"85", x"85", x"85", x"84", x"83", x"83", x"85", x"85", x"85", x"85", x"85", x"86", 
        x"86", x"86", x"84", x"86", x"84", x"83", x"86", x"84", x"82", x"80", x"84", x"86", x"85", x"81", x"80", 
        x"7b", x"7f", x"89", x"90", x"9a", x"a5", x"ac", x"b2", x"c2", x"d2", x"d9", x"d7", x"d3", x"d2", x"d3", 
        x"d3", x"d4", x"d4", x"d3", x"d2", x"d4", x"d4", x"d2", x"d4", x"d5", x"d4", x"d2", x"d5", x"d8", x"d3", 
        x"d5", x"d5", x"d4", x"d5", x"d5", x"d3", x"d3", x"d1", x"d2", x"d3", x"d1", x"d3", x"d2", x"d3", x"d3", 
        x"7f", x"81", x"80", x"7f", x"82", x"81", x"82", x"80", x"7f", x"7e", x"7e", x"7e", x"7e", x"7f", x"7f", 
        x"80", x"80", x"7f", x"7f", x"80", x"7f", x"7f", x"80", x"81", x"81", x"80", x"80", x"7f", x"7e", x"80", 
        x"80", x"7f", x"7f", x"7e", x"7f", x"80", x"7d", x"7d", x"7f", x"81", x"81", x"80", x"7e", x"7f", x"82", 
        x"83", x"81", x"81", x"81", x"81", x"82", x"81", x"80", x"80", x"81", x"82", x"82", x"81", x"7f", x"80", 
        x"80", x"80", x"80", x"81", x"82", x"81", x"80", x"7e", x"82", x"84", x"82", x"82", x"82", x"81", x"80", 
        x"80", x"80", x"80", x"81", x"81", x"82", x"83", x"83", x"81", x"81", x"82", x"82", x"84", x"82", x"83", 
        x"84", x"81", x"83", x"85", x"81", x"82", x"84", x"85", x"84", x"82", x"84", x"87", x"7d", x"6e", x"82", 
        x"b5", x"d3", x"d4", x"ce", x"cb", x"d0", x"cf", x"cd", x"d4", x"d7", x"ce", x"a4", x"57", x"20", x"1c", 
        x"20", x"1d", x"1d", x"1f", x"1e", x"1b", x"1b", x"1b", x"1d", x"1b", x"1c", x"1b", x"18", x"14", x"0e", 
        x"05", x"02", x"02", x"04", x"06", x"07", x"07", x"07", x"06", x"06", x"07", x"08", x"09", x"09", x"0a", 
        x"20", x"a3", x"dd", x"d5", x"d5", x"d2", x"d6", x"d8", x"cf", x"d0", x"d1", x"cf", x"cf", x"d1", x"d1", 
        x"d0", x"d1", x"d1", x"d1", x"d2", x"d2", x"d0", x"cf", x"cf", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", 
        x"d2", x"d1", x"d0", x"d0", x"d1", x"d2", x"d3", x"d2", x"d1", x"d0", x"d0", x"d0", x"d0", x"d2", x"d2", 
        x"d1", x"d2", x"d2", x"d2", x"d0", x"cd", x"cd", x"cd", x"dc", x"d2", x"d4", x"d5", x"d5", x"d5", x"d1", 
        x"d5", x"ed", x"ef", x"ee", x"ef", x"ee", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ee", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"ef", x"f0", x"f2", x"f0", x"ee", x"ef", x"f0", x"ea", x"ec", x"f0", x"ef", x"f0", 
        x"ed", x"f0", x"f0", x"f0", x"ef", x"ee", x"f2", x"f1", x"ee", x"e0", x"c8", x"b1", x"b3", x"c1", x"d0", 
        x"da", x"e4", x"ed", x"f2", x"f2", x"f0", x"ef", x"ee", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f3", x"f4", x"f2", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f3", x"f3", 
        x"f0", x"ef", x"f2", x"f4", x"ee", x"e1", x"ce", x"c2", x"c7", x"d3", x"dd", x"e8", x"ee", x"f3", x"f2", 
        x"f0", x"ef", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"f0", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", 
        x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"f0", x"ee", x"e3", x"d6", x"d4", x"d8", x"d7", x"c1", 
        x"a3", x"85", x"7c", x"82", x"88", x"89", x"8a", x"89", x"8a", x"8b", x"89", x"89", x"8a", x"88", x"89", 
        x"8a", x"89", x"89", x"89", x"89", x"89", x"87", x"87", x"88", x"89", x"89", x"89", x"89", x"88", x"87", 
        x"89", x"89", x"86", x"86", x"88", x"88", x"89", x"88", x"88", x"87", x"88", x"88", x"87", x"89", x"87", 
        x"88", x"89", x"86", x"88", x"87", x"89", x"89", x"88", x"87", x"87", x"89", x"88", x"87", x"85", x"85", 
        x"86", x"86", x"86", x"86", x"88", x"87", x"86", x"88", x"85", x"83", x"88", x"89", x"86", x"84", x"84", 
        x"84", x"83", x"84", x"86", x"87", x"86", x"85", x"87", x"87", x"85", x"86", x"86", x"86", x"86", x"85", 
        x"84", x"84", x"85", x"86", x"86", x"85", x"86", x"88", x"88", x"86", x"86", x"87", x"87", x"86", x"85", 
        x"87", x"85", x"83", x"84", x"85", x"87", x"87", x"85", x"85", x"86", x"84", x"85", x"86", x"85", x"84", 
        x"86", x"87", x"85", x"86", x"84", x"83", x"86", x"87", x"84", x"80", x"80", x"80", x"81", x"82", x"86", 
        x"92", x"a0", x"ad", x"b5", x"bc", x"c9", x"d4", x"d9", x"da", x"d7", x"d4", x"d2", x"d4", x"d4", x"d5", 
        x"d6", x"d5", x"d4", x"d3", x"d2", x"d3", x"d7", x"d7", x"d4", x"d4", x"d5", x"d4", x"d3", x"d2", x"d2", 
        x"d6", x"d5", x"d5", x"d4", x"d5", x"d4", x"d4", x"d2", x"d2", x"d1", x"d1", x"d3", x"d3", x"d4", x"d4", 
        x"83", x"81", x"81", x"82", x"82", x"80", x"81", x"80", x"80", x"80", x"7f", x"7f", x"7e", x"7d", x"7e", 
        x"80", x"81", x"7f", x"7e", x"80", x"7f", x"7e", x"7d", x"7f", x"81", x"80", x"80", x"81", x"80", x"81", 
        x"80", x"80", x"80", x"80", x"80", x"7e", x"7d", x"7d", x"80", x"82", x"80", x"7e", x"7e", x"7f", x"81", 
        x"83", x"83", x"81", x"82", x"84", x"83", x"81", x"81", x"80", x"81", x"82", x"83", x"83", x"7f", x"81", 
        x"82", x"80", x"80", x"81", x"85", x"80", x"80", x"81", x"84", x"85", x"84", x"83", x"83", x"83", x"83", 
        x"84", x"84", x"82", x"80", x"7f", x"80", x"81", x"83", x"83", x"85", x"85", x"83", x"84", x"82", x"83", 
        x"84", x"82", x"82", x"86", x"82", x"83", x"83", x"83", x"84", x"86", x"82", x"76", x"74", x"a3", x"d0", 
        x"d3", x"cf", x"d0", x"ce", x"ce", x"d1", x"d1", x"d5", x"d2", x"ba", x"78", x"37", x"1c", x"1e", x"1e", 
        x"1e", x"1e", x"1d", x"1b", x"1c", x"1e", x"1b", x"19", x"1e", x"1c", x"19", x"16", x"0f", x"06", x"02", 
        x"03", x"03", x"03", x"06", x"08", x"08", x"08", x"06", x"06", x"08", x"0a", x"08", x"07", x"0e", x"12", 
        x"28", x"a6", x"dd", x"d3", x"d2", x"d4", x"d4", x"d9", x"cf", x"d0", x"d0", x"cf", x"d0", x"d2", x"d2", 
        x"d1", x"d2", x"d1", x"cf", x"d1", x"d2", x"d0", x"cf", x"d1", x"d0", x"d0", x"d0", x"d0", x"d1", x"d1", 
        x"d3", x"d2", x"d1", x"d1", x"d2", x"d3", x"d4", x"d4", x"d2", x"d1", x"d2", x"d0", x"ce", x"d1", x"d2", 
        x"d0", x"d3", x"d2", x"d0", x"d1", x"cf", x"cd", x"ca", x"d9", x"d2", x"d2", x"d4", x"d3", x"d2", x"d2", 
        x"d4", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f2", x"f1", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ea", x"ed", x"f1", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f1", x"f0", x"e9", x"dc", x"ca", x"b6", 
        x"b5", x"bd", x"ca", x"d8", x"e6", x"f1", x"f3", x"ef", x"ee", x"f0", x"ef", x"f1", x"f0", x"f1", x"f3", 
        x"f0", x"ef", x"f0", x"f2", x"f2", x"f2", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f0", x"f2", x"ef", x"e5", x"da", x"cb", x"c3", x"ca", x"d5", x"e4", x"ec", 
        x"f0", x"f0", x"ef", x"f0", x"f2", x"f1", x"f0", x"ee", x"ef", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"ee", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"ee", x"e4", x"d8", x"d1", x"da", 
        x"da", x"c9", x"a4", x"8a", x"80", x"7f", x"84", x"8a", x"8e", x"8c", x"8a", x"89", x"8a", x"8b", x"8a", 
        x"89", x"89", x"8a", x"8b", x"8b", x"8a", x"88", x"8a", x"8a", x"8a", x"8b", x"8d", x"8b", x"87", x"87", 
        x"89", x"89", x"87", x"86", x"89", x"89", x"8a", x"89", x"8a", x"88", x"89", x"89", x"87", x"86", x"88", 
        x"8a", x"87", x"85", x"86", x"87", x"88", x"87", x"86", x"88", x"8a", x"88", x"88", x"88", x"87", x"86", 
        x"86", x"86", x"86", x"86", x"88", x"87", x"86", x"88", x"86", x"85", x"87", x"88", x"87", x"86", x"85", 
        x"84", x"83", x"84", x"86", x"83", x"84", x"84", x"86", x"87", x"85", x"85", x"84", x"85", x"87", x"86", 
        x"85", x"86", x"83", x"86", x"87", x"83", x"85", x"87", x"85", x"85", x"87", x"87", x"87", x"87", x"88", 
        x"8a", x"87", x"83", x"84", x"84", x"87", x"89", x"87", x"85", x"86", x"84", x"86", x"87", x"84", x"84", 
        x"87", x"84", x"85", x"86", x"87", x"85", x"83", x"82", x"81", x"82", x"85", x"8b", x"95", x"a3", x"ae", 
        x"b5", x"be", x"cc", x"d6", x"db", x"d9", x"d6", x"d4", x"d5", x"d5", x"d5", x"d5", x"d5", x"d5", x"d5", 
        x"d4", x"d5", x"d3", x"d4", x"d3", x"d4", x"d8", x"d9", x"d3", x"d2", x"d4", x"d4", x"d2", x"d2", x"d3", 
        x"d6", x"d5", x"d6", x"d3", x"d5", x"d5", x"d5", x"d3", x"d3", x"d5", x"d7", x"d8", x"d8", x"d0", x"c4", 
        x"82", x"81", x"83", x"83", x"80", x"7f", x"82", x"82", x"81", x"7f", x"7e", x"7e", x"7e", x"7f", x"7f", 
        x"80", x"81", x"7f", x"7f", x"80", x"80", x"7f", x"7e", x"7e", x"80", x"7e", x"7f", x"81", x"7f", x"7e", 
        x"7e", x"7f", x"81", x"81", x"7f", x"7d", x"7f", x"7f", x"7f", x"80", x"81", x"80", x"80", x"7f", x"80", 
        x"81", x"81", x"81", x"81", x"82", x"82", x"82", x"82", x"82", x"82", x"81", x"81", x"82", x"81", x"82", 
        x"82", x"81", x"81", x"81", x"83", x"81", x"82", x"83", x"83", x"83", x"83", x"83", x"82", x"81", x"81", 
        x"82", x"82", x"81", x"80", x"82", x"82", x"81", x"80", x"81", x"83", x"84", x"86", x"85", x"82", x"84", 
        x"86", x"82", x"81", x"83", x"83", x"85", x"81", x"85", x"85", x"73", x"6d", x"8c", x"c2", x"da", x"d6", 
        x"ce", x"d0", x"cf", x"d1", x"d4", x"d5", x"d9", x"cc", x"92", x"4b", x"1c", x"1e", x"23", x"20", x"1b", 
        x"1c", x"1e", x"1c", x"19", x"1a", x"1f", x"1e", x"1b", x"1a", x"14", x"0e", x"07", x"02", x"00", x"02", 
        x"05", x"05", x"05", x"06", x"06", x"07", x"06", x"06", x"07", x"09", x"07", x"07", x"12", x"23", x"27", 
        x"35", x"a4", x"dc", x"d4", x"d5", x"d5", x"d4", x"d8", x"d0", x"d1", x"d2", x"cf", x"cf", x"d0", x"cf", 
        x"d1", x"d2", x"d2", x"d0", x"d1", x"d2", x"d0", x"d0", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"d1", 
        x"d3", x"d2", x"d0", x"d0", x"d2", x"d4", x"d5", x"d4", x"d2", x"d1", x"d2", x"d0", x"ce", x"d2", x"d3", 
        x"d1", x"d2", x"d1", x"d0", x"d2", x"d0", x"ce", x"cb", x"db", x"d4", x"d4", x"d3", x"d1", x"d1", x"d3", 
        x"d4", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f2", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"eb", x"ed", x"f1", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"f1", x"f5", x"f4", x"e9", 
        x"e3", x"cb", x"b8", x"b0", x"b7", x"c4", x"d6", x"e7", x"f0", x"f2", x"f0", x"f2", x"ef", x"ee", x"f2", 
        x"f0", x"ef", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"ee", x"f0", x"ef", x"ea", x"d6", x"cb", x"c1", x"c5", 
        x"d3", x"e6", x"f0", x"f3", x"f2", x"ef", x"ee", x"f0", x"f3", x"f1", x"f2", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"ee", 
        x"f0", x"f1", x"ef", x"f1", x"f1", x"ef", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"ef", x"e8", x"db", 
        x"d7", x"d5", x"da", x"d2", x"b5", x"8f", x"7c", x"7c", x"84", x"8d", x"8e", x"8a", x"87", x"89", x"8a", 
        x"8b", x"8b", x"8a", x"89", x"8b", x"8c", x"8c", x"8c", x"8b", x"8a", x"8a", x"8b", x"8b", x"88", x"87", 
        x"88", x"89", x"87", x"88", x"89", x"88", x"89", x"88", x"89", x"88", x"89", x"88", x"88", x"86", x"86", 
        x"87", x"86", x"86", x"87", x"88", x"89", x"87", x"86", x"87", x"89", x"88", x"87", x"87", x"88", x"88", 
        x"87", x"87", x"86", x"86", x"88", x"87", x"84", x"86", x"85", x"85", x"87", x"87", x"87", x"88", x"87", 
        x"86", x"86", x"86", x"86", x"84", x"87", x"86", x"86", x"85", x"83", x"87", x"86", x"85", x"85", x"86", 
        x"88", x"89", x"83", x"86", x"88", x"85", x"86", x"87", x"84", x"85", x"86", x"86", x"85", x"86", x"87", 
        x"88", x"85", x"84", x"87", x"86", x"85", x"86", x"86", x"84", x"83", x"85", x"86", x"86", x"84", x"85", 
        x"86", x"83", x"83", x"80", x"7b", x"7e", x"84", x"89", x"8d", x"96", x"a5", x"b3", x"bf", x"c8", x"cf", 
        x"d9", x"db", x"d9", x"d7", x"d5", x"d4", x"d5", x"d4", x"d5", x"d6", x"d6", x"d5", x"d5", x"d5", x"d5", 
        x"d4", x"d5", x"d3", x"d6", x"d5", x"d4", x"d7", x"d7", x"d4", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", 
        x"d6", x"d6", x"d7", x"d5", x"d5", x"d3", x"d4", x"d8", x"dd", x"db", x"ce", x"be", x"b3", x"a6", x"96", 
        x"82", x"82", x"83", x"84", x"81", x"7f", x"82", x"81", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
        x"80", x"81", x"80", x"7f", x"80", x"80", x"81", x"82", x"81", x"83", x"80", x"82", x"83", x"81", x"7f", 
        x"7f", x"7f", x"80", x"80", x"7e", x"7d", x"7e", x"7e", x"7d", x"7d", x"7f", x"81", x"80", x"81", x"81", 
        x"82", x"83", x"83", x"83", x"83", x"82", x"82", x"82", x"83", x"82", x"81", x"80", x"82", x"82", x"82", 
        x"82", x"82", x"82", x"81", x"82", x"82", x"83", x"84", x"83", x"82", x"82", x"82", x"81", x"80", x"80", 
        x"81", x"81", x"81", x"81", x"84", x"85", x"85", x"85", x"84", x"83", x"83", x"80", x"84", x"85", x"85", 
        x"85", x"84", x"82", x"80", x"83", x"88", x"8a", x"7e", x"6e", x"81", x"b3", x"d3", x"d3", x"d0", x"d4", 
        x"cb", x"ce", x"d0", x"d2", x"d9", x"d8", x"ac", x"5f", x"2d", x"19", x"20", x"22", x"20", x"20", x"20", 
        x"1e", x"1e", x"1d", x"1d", x"1d", x"1c", x"19", x"16", x"13", x"09", x"03", x"01", x"02", x"05", x"06", 
        x"05", x"05", x"06", x"05", x"05", x"06", x"08", x"07", x"07", x"07", x"0e", x"19", x"27", x"32", x"30", 
        x"38", x"a2", x"db", x"d4", x"d6", x"d7", x"d5", x"d8", x"d0", x"d2", x"d3", x"d0", x"d0", x"d0", x"ce", 
        x"cf", x"d1", x"d3", x"d1", x"cf", x"cf", x"d0", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", 
        x"d3", x"d2", x"d0", x"d0", x"d2", x"d3", x"d4", x"d3", x"d2", x"d1", x"d2", x"d0", x"ce", x"d2", x"d3", 
        x"d1", x"d2", x"d1", x"cf", x"d2", x"d1", x"d0", x"cf", x"e0", x"d8", x"d7", x"d6", x"d3", x"d3", x"d4", 
        x"d6", x"ee", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f2", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ea", x"ed", x"f2", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"ee", 
        x"f1", x"f0", x"e9", x"de", x"d2", x"c5", x"bc", x"ba", x"bf", x"d3", x"e4", x"ef", x"f1", x"f0", x"ee", 
        x"ee", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ed", x"f0", x"f1", x"f2", x"f3", x"ee", x"e3", x"d2", 
        x"c5", x"c1", x"c7", x"d3", x"e5", x"f2", x"f3", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"ee", 
        x"ef", x"f1", x"ef", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", 
        x"ea", x"e0", x"d7", x"d7", x"d7", x"d2", x"bf", x"9f", x"80", x"7d", x"86", x"8d", x"8c", x"8c", x"8b", 
        x"8b", x"8c", x"8c", x"8a", x"89", x"89", x"8a", x"8a", x"8a", x"88", x"88", x"8a", x"8b", x"89", x"88", 
        x"88", x"89", x"88", x"89", x"8a", x"88", x"88", x"87", x"89", x"88", x"88", x"87", x"87", x"87", x"88", 
        x"88", x"87", x"86", x"86", x"88", x"8a", x"89", x"87", x"87", x"88", x"88", x"86", x"86", x"87", x"88", 
        x"88", x"87", x"87", x"86", x"87", x"86", x"85", x"87", x"87", x"86", x"89", x"89", x"89", x"88", x"88", 
        x"87", x"86", x"86", x"87", x"86", x"87", x"86", x"86", x"86", x"84", x"86", x"87", x"87", x"86", x"88", 
        x"89", x"87", x"84", x"88", x"89", x"86", x"86", x"88", x"85", x"86", x"86", x"84", x"84", x"85", x"87", 
        x"86", x"85", x"87", x"8b", x"8a", x"88", x"86", x"85", x"85", x"85", x"84", x"85", x"87", x"87", x"84", 
        x"80", x"7e", x"82", x"85", x"89", x"94", x"a2", x"ae", x"b8", x"c1", x"cc", x"d4", x"d9", x"da", x"d9", 
        x"d7", x"d7", x"d8", x"d8", x"d7", x"d5", x"d4", x"d4", x"d5", x"d6", x"d5", x"d3", x"d4", x"d5", x"d5", 
        x"d5", x"d5", x"d4", x"d7", x"d7", x"d5", x"d6", x"d5", x"d3", x"d5", x"d7", x"d6", x"d5", x"d6", x"d5", 
        x"d7", x"d6", x"d6", x"d5", x"d9", x"db", x"d5", x"c8", x"ba", x"ad", x"9f", x"97", x"95", x"9a", x"9b", 
        x"84", x"82", x"82", x"84", x"82", x"81", x"81", x"80", x"7f", x"80", x"81", x"81", x"80", x"7f", x"80", 
        x"80", x"82", x"81", x"80", x"80", x"81", x"81", x"80", x"81", x"83", x"81", x"81", x"81", x"80", x"80", 
        x"7f", x"7f", x"80", x"80", x"80", x"7f", x"81", x"81", x"7f", x"7e", x"80", x"81", x"7f", x"82", x"82", 
        x"83", x"84", x"84", x"84", x"84", x"83", x"82", x"82", x"82", x"82", x"81", x"80", x"81", x"82", x"81", 
        x"81", x"83", x"83", x"83", x"81", x"82", x"83", x"84", x"83", x"82", x"83", x"84", x"82", x"82", x"82", 
        x"82", x"82", x"83", x"83", x"83", x"83", x"84", x"85", x"84", x"83", x"82", x"82", x"83", x"84", x"81", 
        x"81", x"83", x"83", x"83", x"89", x"8b", x"74", x"6f", x"98", x"ca", x"da", x"d9", x"cd", x"ce", x"d1", 
        x"cf", x"d3", x"d5", x"da", x"c5", x"88", x"41", x"1f", x"1d", x"1e", x"1f", x"22", x"22", x"24", x"24", 
        x"1e", x"1f", x"1e", x"20", x"20", x"1a", x"11", x"0b", x"07", x"03", x"01", x"02", x"04", x"07", x"08", 
        x"07", x"06", x"07", x"08", x"09", x"08", x"08", x"09", x"0d", x"16", x"24", x"2f", x"31", x"34", x"32", 
        x"3a", x"a3", x"dc", x"d4", x"d6", x"d7", x"d6", x"d9", x"cf", x"d1", x"d2", x"d1", x"d1", x"d1", x"cf", 
        x"ce", x"d1", x"d3", x"d1", x"ce", x"cd", x"d0", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", 
        x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d2", x"d0", x"d2", x"d1", x"cf", x"d3", x"d2", 
        x"d1", x"d2", x"d2", x"d0", x"d2", x"d0", x"d0", x"ce", x"de", x"d6", x"d6", x"d6", x"d4", x"d3", x"d5", 
        x"d6", x"ee", x"ef", x"f0", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ea", x"ed", x"f2", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f0", x"f1", x"f0", x"ef", x"ed", 
        x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"e3", x"d1", x"c1", x"bb", x"ba", x"c7", x"da", x"e7", x"ef", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", x"ee", x"f1", x"f2", x"f3", x"f2", x"f1", x"f2", x"f1", 
        x"eb", x"d9", x"c8", x"c0", x"bf", x"c8", x"dd", x"ed", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", 
        x"f3", x"f2", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"ed", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"ed", 
        x"f2", x"f3", x"eb", x"e2", x"da", x"d5", x"d7", x"d5", x"c4", x"a2", x"86", x"7b", x"82", x"8b", x"8b", 
        x"89", x"8a", x"8e", x"8e", x"8b", x"8a", x"8b", x"8b", x"8a", x"89", x"8a", x"8b", x"8c", x"8a", x"89", 
        x"89", x"89", x"89", x"8a", x"8a", x"89", x"88", x"87", x"88", x"89", x"88", x"87", x"88", x"88", x"87", 
        x"86", x"87", x"87", x"88", x"89", x"8a", x"89", x"88", x"86", x"87", x"88", x"88", x"87", x"87", x"87", 
        x"87", x"88", x"88", x"87", x"89", x"89", x"88", x"8a", x"88", x"86", x"88", x"88", x"88", x"88", x"88", 
        x"87", x"85", x"86", x"87", x"85", x"87", x"86", x"86", x"88", x"86", x"84", x"87", x"87", x"86", x"88", 
        x"88", x"85", x"87", x"89", x"88", x"86", x"87", x"88", x"87", x"87", x"87", x"85", x"85", x"86", x"87", 
        x"86", x"86", x"85", x"85", x"85", x"86", x"86", x"87", x"88", x"88", x"86", x"87", x"84", x"7f", x"80", 
        x"85", x"8b", x"94", x"a1", x"ad", x"b9", x"c5", x"d0", x"d5", x"d8", x"db", x"d9", x"d6", x"d3", x"d4", 
        x"d6", x"d7", x"d8", x"d8", x"d8", x"d8", x"d6", x"d6", x"d6", x"d6", x"d5", x"d4", x"d3", x"d5", x"d6", 
        x"d6", x"d5", x"d3", x"d6", x"d7", x"d5", x"d6", x"d6", x"d3", x"d5", x"d6", x"d5", x"d5", x"d6", x"d5", 
        x"d7", x"db", x"db", x"d4", x"c5", x"b8", x"a8", x"9b", x"94", x"96", x"9b", x"9d", x"9f", x"a0", x"a4", 
        x"85", x"81", x"80", x"83", x"84", x"82", x"81", x"80", x"7f", x"7f", x"7f", x"80", x"80", x"81", x"82", 
        x"81", x"82", x"82", x"81", x"80", x"81", x"81", x"7f", x"80", x"83", x"81", x"81", x"81", x"7f", x"80", 
        x"7e", x"7d", x"7f", x"81", x"83", x"83", x"7f", x"7f", x"7e", x"80", x"83", x"83", x"81", x"81", x"81", 
        x"82", x"83", x"82", x"83", x"83", x"83", x"83", x"82", x"82", x"82", x"81", x"81", x"81", x"82", x"80", 
        x"80", x"83", x"85", x"85", x"82", x"82", x"83", x"83", x"83", x"83", x"84", x"85", x"83", x"84", x"84", 
        x"84", x"83", x"83", x"84", x"84", x"83", x"83", x"83", x"83", x"84", x"85", x"84", x"84", x"87", x"88", 
        x"85", x"85", x"87", x"8f", x"7e", x"61", x"7d", x"b7", x"d6", x"d5", x"d0", x"d6", x"d0", x"cf", x"d0", 
        x"d2", x"de", x"d9", x"ac", x"51", x"26", x"1a", x"1f", x"24", x"20", x"1f", x"20", x"1e", x"1e", x"1e", 
        x"19", x"1b", x"1f", x"1d", x"18", x"10", x"08", x"03", x"01", x"03", x"04", x"05", x"05", x"06", x"07", 
        x"08", x"08", x"08", x"0a", x"09", x"08", x"0c", x"16", x"22", x"2f", x"31", x"33", x"32", x"36", x"33", 
        x"39", x"a5", x"dc", x"d4", x"d5", x"d6", x"d6", x"da", x"ce", x"d0", x"d1", x"d1", x"d2", x"d3", x"d2", 
        x"d0", x"d0", x"d1", x"d1", x"ce", x"cd", x"d0", x"d2", x"d3", x"d2", x"d1", x"d1", x"d2", x"d3", x"d2", 
        x"d2", x"d2", x"d3", x"d3", x"d3", x"d3", x"d3", x"d2", x"d1", x"d0", x"d2", x"d1", x"d0", x"d3", x"d2", 
        x"d1", x"d3", x"d3", x"d1", x"d1", x"d0", x"d0", x"cd", x"db", x"d3", x"d4", x"d5", x"d5", x"d3", x"d6", 
        x"d7", x"ee", x"ef", x"f1", x"f0", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f2", x"f1", x"f0", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ea", x"ed", x"f2", x"f0", x"f0", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"f2", x"f0", x"ee", x"f0", 
        x"f3", x"f2", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"e9", x"e7", x"de", x"ce", x"b8", x"b7", x"c4", 
        x"d9", x"e9", x"f2", x"f4", x"f1", x"ee", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ed", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", 
        x"ef", x"ed", x"ee", x"ea", x"da", x"c8", x"bc", x"bb", x"ce", x"e7", x"f1", x"f2", x"f5", x"f2", x"f1", 
        x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"ed", 
        x"ee", x"f0", x"ee", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"f0", x"ee", x"e7", x"e1", x"db", x"d7", x"db", x"d6", x"b5", x"88", x"73", x"7e", 
        x"8a", x"8b", x"8a", x"8b", x"8a", x"8c", x"8d", x"8d", x"8b", x"89", x"89", x"8a", x"8b", x"8a", x"8a", 
        x"89", x"89", x"8a", x"8a", x"89", x"89", x"88", x"88", x"89", x"89", x"88", x"88", x"88", x"88", x"86", 
        x"85", x"87", x"88", x"88", x"89", x"89", x"88", x"88", x"87", x"87", x"89", x"8a", x"88", x"87", x"87", 
        x"87", x"87", x"88", x"86", x"87", x"88", x"89", x"8c", x"8b", x"89", x"88", x"86", x"86", x"87", x"87", 
        x"88", x"87", x"87", x"85", x"86", x"89", x"88", x"87", x"89", x"87", x"85", x"86", x"85", x"84", x"86", 
        x"87", x"87", x"89", x"89", x"88", x"86", x"87", x"87", x"87", x"88", x"88", x"87", x"86", x"88", x"88", 
        x"88", x"87", x"85", x"84", x"86", x"87", x"86", x"85", x"83", x"80", x"7e", x"83", x"8a", x"90", x"99", 
        x"a5", x"ad", x"ba", x"ca", x"d6", x"d7", x"d7", x"d8", x"d7", x"d6", x"d4", x"d5", x"d7", x"d7", x"d7", 
        x"d7", x"d7", x"d8", x"d8", x"d7", x"d5", x"d4", x"d5", x"d7", x"d6", x"d5", x"d5", x"d4", x"d4", x"d5", 
        x"d7", x"d5", x"d2", x"d5", x"d6", x"d6", x"d7", x"d4", x"d3", x"d5", x"d6", x"d6", x"d8", x"dc", x"dd", 
        x"d2", x"bf", x"a9", x"9a", x"95", x"97", x"9a", x"9b", x"9d", x"9e", x"a2", x"a6", x"a9", x"af", x"b2", 
        x"84", x"82", x"82", x"84", x"83", x"81", x"82", x"81", x"80", x"7f", x"7f", x"80", x"81", x"82", x"82", 
        x"81", x"82", x"83", x"82", x"80", x"82", x"83", x"80", x"81", x"84", x"82", x"83", x"84", x"81", x"80", 
        x"7e", x"7e", x"7f", x"80", x"81", x"81", x"81", x"7e", x"7d", x"7f", x"81", x"7f", x"7e", x"7f", x"81", 
        x"82", x"83", x"82", x"82", x"84", x"82", x"82", x"83", x"84", x"84", x"83", x"82", x"81", x"84", x"82", 
        x"81", x"82", x"84", x"86", x"83", x"84", x"83", x"82", x"83", x"83", x"84", x"84", x"83", x"85", x"85", 
        x"84", x"83", x"82", x"83", x"86", x"85", x"85", x"84", x"85", x"86", x"87", x"83", x"82", x"84", x"83", 
        x"86", x"8a", x"86", x"6e", x"72", x"9c", x"cd", x"d4", x"cd", x"cc", x"cf", x"d6", x"ce", x"cd", x"d4", 
        x"d7", x"be", x"78", x"34", x"1d", x"1d", x"23", x"20", x"1e", x"22", x"22", x"20", x"1e", x"1e", x"1c", 
        x"19", x"1b", x"19", x"11", x"08", x"04", x"02", x"02", x"03", x"02", x"03", x"06", x"08", x"0a", x"09", 
        x"08", x"08", x"09", x"08", x"0c", x"13", x"20", x"2b", x"34", x"35", x"32", x"33", x"32", x"38", x"36", 
        x"3b", x"a6", x"dd", x"d4", x"d4", x"d6", x"d6", x"da", x"cf", x"d0", x"d1", x"d1", x"d2", x"d4", x"d3", 
        x"d2", x"d1", x"d2", x"d2", x"d0", x"ce", x"d0", x"d2", x"d1", x"d2", x"d1", x"d1", x"d2", x"d1", x"d2", 
        x"d4", x"d3", x"d2", x"d3", x"d3", x"d4", x"d4", x"d2", x"d1", x"d0", x"d2", x"d1", x"d0", x"d3", x"d2", 
        x"d1", x"d3", x"d2", x"d0", x"d2", x"d0", x"d2", x"cf", x"dd", x"d4", x"d4", x"d5", x"d5", x"d3", x"d6", 
        x"d8", x"ed", x"ee", x"f0", x"f0", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f2", x"f1", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"eb", x"ed", x"f2", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"ee", x"f2", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"ef", x"ee", x"f0", x"f1", x"ef", x"ed", x"eb", x"ee", x"ef", x"ee", x"e9", x"de", x"d0", 
        x"be", x"be", x"c9", x"d7", x"e5", x"ed", x"f1", x"f2", x"f3", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f2", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"f0", x"ee", x"f0", x"ee", x"ee", x"f2", x"f3", x"f1", x"f0", 
        x"f0", x"f2", x"f2", x"f1", x"ef", x"ed", x"e6", x"d7", x"c5", x"ba", x"c2", x"d6", x"e6", x"ef", x"ef", 
        x"ef", x"f1", x"f1", x"ef", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"ed", 
        x"ed", x"ef", x"ee", x"f0", x"f2", x"f0", x"f0", x"ef", x"f1", x"f3", x"f4", x"f3", x"f1", x"ef", x"ed", 
        x"ee", x"ef", x"f1", x"ef", x"ef", x"f0", x"ee", x"eb", x"e5", x"e1", x"df", x"db", x"d4", x"bb", x"97", 
        x"7b", x"7d", x"86", x"89", x"8a", x"8b", x"8b", x"8b", x"8a", x"87", x"87", x"88", x"89", x"8a", x"8a", 
        x"89", x"89", x"8a", x"8a", x"88", x"89", x"89", x"8a", x"88", x"8a", x"88", x"88", x"86", x"89", x"89", 
        x"88", x"89", x"87", x"85", x"89", x"87", x"88", x"89", x"88", x"88", x"8a", x"8a", x"89", x"88", x"88", 
        x"87", x"87", x"86", x"86", x"88", x"87", x"87", x"89", x"88", x"87", x"88", x"85", x"86", x"87", x"88", 
        x"88", x"87", x"88", x"86", x"88", x"8a", x"88", x"87", x"89", x"88", x"88", x"86", x"86", x"86", x"87", 
        x"87", x"88", x"89", x"89", x"88", x"88", x"88", x"87", x"85", x"86", x"87", x"87", x"87", x"87", x"88", 
        x"89", x"8a", x"88", x"88", x"88", x"85", x"7f", x"7f", x"82", x"88", x"94", x"a2", x"ac", x"b2", x"bc", 
        x"c9", x"d6", x"d8", x"d9", x"d8", x"d6", x"d5", x"d6", x"d4", x"d6", x"d7", x"d6", x"d4", x"d5", x"d9", 
        x"d9", x"d8", x"d7", x"d6", x"d6", x"d8", x"d9", x"d8", x"d6", x"d5", x"d5", x"d6", x"d5", x"d3", x"d2", 
        x"d6", x"d6", x"d4", x"d6", x"d6", x"d5", x"d9", x"d9", x"d6", x"d9", x"da", x"d4", x"c8", x"bc", x"a2", 
        x"97", x"95", x"96", x"9d", x"a0", x"a1", x"a4", x"a5", x"a6", x"a9", x"ad", x"a9", x"9d", x"85", x"60", 
        x"83", x"83", x"84", x"85", x"82", x"80", x"83", x"80", x"7f", x"80", x"81", x"81", x"81", x"81", x"81", 
        x"81", x"82", x"83", x"82", x"81", x"82", x"82", x"7f", x"7f", x"81", x"80", x"81", x"83", x"82", x"82", 
        x"81", x"80", x"7f", x"7f", x"7e", x"7e", x"82", x"7f", x"7e", x"81", x"82", x"81", x"82", x"81", x"83", 
        x"85", x"84", x"83", x"83", x"85", x"82", x"82", x"84", x"85", x"85", x"84", x"83", x"82", x"85", x"83", 
        x"81", x"81", x"83", x"86", x"84", x"85", x"83", x"82", x"83", x"84", x"83", x"83", x"83", x"84", x"85", 
        x"85", x"84", x"82", x"82", x"83", x"84", x"84", x"84", x"84", x"83", x"82", x"81", x"82", x"83", x"86", 
        x"8a", x"7f", x"69", x"86", x"bc", x"d8", x"d3", x"d0", x"d2", x"d0", x"cf", x"d8", x"d4", x"d5", x"d5", 
        x"9c", x"47", x"22", x"20", x"22", x"22", x"1f", x"1f", x"22", x"1e", x"1c", x"1d", x"1c", x"1d", x"1e", 
        x"1c", x"16", x"0e", x"06", x"02", x"03", x"03", x"03", x"03", x"03", x"03", x"05", x"08", x"0b", x"0d", 
        x"0a", x"0a", x"0a", x"0d", x"1a", x"2a", x"34", x"35", x"34", x"33", x"35", x"37", x"36", x"3b", x"3d", 
        x"42", x"a6", x"de", x"d4", x"d5", x"d5", x"d5", x"d9", x"d0", x"d1", x"d2", x"d0", x"d1", x"d3", x"d3", 
        x"d3", x"d2", x"d2", x"d3", x"d1", x"d0", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", 
        x"d5", x"d3", x"d1", x"d1", x"d3", x"d5", x"d5", x"d2", x"d1", x"d0", x"d2", x"d1", x"d0", x"d3", x"d4", 
        x"d2", x"d2", x"d1", x"d0", x"d2", x"d2", x"d1", x"ce", x"dc", x"d2", x"d2", x"d2", x"d2", x"d2", x"d5", 
        x"d7", x"ec", x"ee", x"f0", x"f0", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"ed", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f2", x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", 
        x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"eb", x"ed", x"f2", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ee", x"f2", x"f0", x"ef", x"f1", 
        x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"ee", x"ed", x"ef", 
        x"ec", x"e1", x"d0", x"be", x"b8", x"c5", x"d9", x"e8", x"ee", x"f1", x"f1", x"f0", x"ef", x"f0", x"f2", 
        x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ed", x"f1", x"f2", x"f2", x"ef", x"ef", x"f0", x"f2", 
        x"f3", x"f2", x"f1", x"f0", x"f3", x"f3", x"f1", x"f1", x"ee", x"e3", x"cb", x"bc", x"bb", x"c9", x"e1", 
        x"ed", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f2", x"f2", x"f2", x"f3", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"ec", 
        x"ed", x"ef", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"f0", x"f1", x"f2", x"f1", x"f0", x"ef", x"ed", x"e7", x"dd", x"d7", x"dc", x"d9", 
        x"c1", x"9b", x"7e", x"7b", x"86", x"89", x"8b", x"8c", x"8b", x"8a", x"8b", x"8c", x"8a", x"89", x"8a", 
        x"89", x"89", x"8a", x"89", x"88", x"8a", x"8a", x"8b", x"88", x"8a", x"89", x"89", x"88", x"89", x"88", 
        x"87", x"89", x"88", x"86", x"88", x"87", x"87", x"8a", x"8a", x"8a", x"8a", x"89", x"89", x"89", x"89", 
        x"88", x"87", x"86", x"85", x"87", x"86", x"84", x"87", x"87", x"88", x"8a", x"88", x"88", x"88", x"88", 
        x"88", x"87", x"88", x"89", x"89", x"89", x"86", x"86", x"88", x"89", x"88", x"87", x"89", x"8a", x"88", 
        x"87", x"88", x"89", x"88", x"88", x"89", x"89", x"87", x"84", x"84", x"86", x"87", x"88", x"87", x"87", 
        x"88", x"89", x"87", x"82", x"81", x"81", x"88", x"97", x"a4", x"a9", x"af", x"ba", x"c9", x"d4", x"d8", 
        x"d7", x"d6", x"d9", x"d8", x"d6", x"d6", x"d7", x"d6", x"d7", x"d8", x"d8", x"d7", x"d7", x"d7", x"d8", 
        x"d8", x"d7", x"d7", x"d7", x"d7", x"d7", x"d7", x"d7", x"d6", x"d5", x"d5", x"d6", x"d5", x"d3", x"d2", 
        x"d5", x"d6", x"d5", x"d8", x"d8", x"d7", x"d8", x"d6", x"d4", x"cb", x"b7", x"9f", x"93", x"93", x"9c", 
        x"9d", x"a0", x"a1", x"a4", x"a5", x"a7", x"a9", x"ab", x"a6", x"99", x"7f", x"56", x"2d", x"1d", x"1c", 
        x"84", x"82", x"83", x"86", x"84", x"81", x"81", x"81", x"81", x"82", x"82", x"82", x"82", x"82", x"7e", 
        x"80", x"83", x"81", x"82", x"85", x"83", x"81", x"82", x"83", x"81", x"81", x"83", x"83", x"82", x"82", 
        x"82", x"82", x"82", x"82", x"82", x"81", x"81", x"81", x"82", x"83", x"83", x"81", x"81", x"81", x"82", 
        x"82", x"83", x"83", x"83", x"83", x"82", x"82", x"82", x"82", x"82", x"82", x"82", x"82", x"83", x"83", 
        x"83", x"83", x"84", x"85", x"84", x"81", x"82", x"82", x"83", x"84", x"84", x"84", x"82", x"81", x"82", 
        x"84", x"85", x"86", x"87", x"84", x"85", x"85", x"84", x"85", x"85", x"83", x"82", x"81", x"84", x"86", 
        x"70", x"70", x"9f", x"d2", x"d5", x"d0", x"d3", x"d4", x"d3", x"d1", x"d3", x"dc", x"db", x"b3", x"6c", 
        x"2d", x"1b", x"23", x"23", x"1f", x"1e", x"1f", x"21", x"21", x"1e", x"1c", x"1f", x"21", x"21", x"1b", 
        x"11", x"08", x"05", x"03", x"06", x"06", x"02", x"03", x"03", x"02", x"02", x"05", x"09", x"0b", x"0b", 
        x"0c", x"10", x"18", x"28", x"33", x"34", x"30", x"33", x"35", x"35", x"34", x"36", x"45", x"47", x"3d", 
        x"3a", x"a4", x"de", x"d4", x"d6", x"d3", x"d5", x"d9", x"d0", x"d1", x"d3", x"d0", x"d0", x"d1", x"d1", 
        x"d0", x"d2", x"d2", x"d0", x"d0", x"d2", x"d2", x"d2", x"d0", x"d1", x"d4", x"d2", x"d1", x"d2", x"d3", 
        x"d4", x"d3", x"d3", x"d3", x"d3", x"d3", x"d2", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d6", 
        x"d3", x"d3", x"d3", x"d2", x"d2", x"d4", x"cf", x"cf", x"dd", x"d3", x"d5", x"d5", x"d2", x"d2", x"d3", 
        x"d5", x"ed", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ed", x"ee", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", 
        x"ed", x"ee", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f1", x"f0", x"ef", x"ee", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ea", x"ee", x"f0", x"f0", x"ef", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", 
        x"f1", x"f0", x"ef", x"ec", x"e3", x"d3", x"c0", x"bb", x"c5", x"d5", x"e5", x"eb", x"ed", x"ef", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f2", x"f1", x"ee", x"ef", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ed", x"f0", x"f4", x"f2", x"f1", x"f2", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"ec", x"dd", x"c6", x"b7", 
        x"c1", x"d4", x"e5", x"ed", x"f0", x"f1", x"f1", x"f2", x"f1", x"ee", x"ee", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f3", x"f3", x"f1", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"ee", 
        x"ed", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"e9", x"dd", x"da", 
        x"dd", x"dc", x"ca", x"a4", x"8a", x"83", x"86", x"89", x"8a", x"8b", x"8d", x"8c", x"8b", x"8a", x"89", 
        x"8a", x"8a", x"8a", x"8b", x"8c", x"8b", x"8d", x"8b", x"89", x"8a", x"8b", x"89", x"8b", x"87", x"87", 
        x"88", x"89", x"88", x"88", x"86", x"88", x"88", x"88", x"8a", x"8b", x"8a", x"88", x"88", x"89", x"8a", 
        x"8a", x"89", x"89", x"87", x"89", x"8a", x"87", x"86", x"87", x"89", x"88", x"87", x"87", x"89", x"89", 
        x"8a", x"89", x"88", x"87", x"8a", x"89", x"87", x"89", x"88", x"87", x"89", x"86", x"88", x"88", x"87", 
        x"89", x"89", x"8a", x"8b", x"89", x"87", x"87", x"89", x"88", x"87", x"88", x"8b", x"8a", x"87", x"84", 
        x"82", x"81", x"83", x"8c", x"98", x"a4", x"a6", x"a9", x"b6", x"ca", x"d7", x"dc", x"d9", x"d6", x"d6", 
        x"d6", x"d7", x"d8", x"d8", x"d7", x"d7", x"d6", x"d5", x"d5", x"d6", x"d7", x"d6", x"d6", x"d6", x"d8", 
        x"d9", x"d7", x"d7", x"d8", x"d7", x"d5", x"d6", x"d7", x"d5", x"d5", x"d7", x"d6", x"d4", x"d4", x"d7", 
        x"d7", x"d7", x"d6", x"d6", x"d5", x"cd", x"c0", x"ae", x"9e", x"95", x"98", x"9c", x"a0", x"a1", x"a4", 
        x"a5", x"ab", x"ad", x"ac", x"aa", x"a3", x"90", x"71", x"49", x"2a", x"1d", x"1f", x"22", x"38", x"50", 
        x"87", x"84", x"83", x"84", x"83", x"81", x"81", x"81", x"81", x"83", x"84", x"83", x"82", x"81", x"7e", 
        x"80", x"82", x"80", x"81", x"84", x"82", x"81", x"82", x"83", x"81", x"81", x"82", x"83", x"82", x"82", 
        x"83", x"83", x"83", x"83", x"83", x"82", x"7f", x"80", x"82", x"83", x"83", x"84", x"83", x"82", x"82", 
        x"82", x"83", x"83", x"83", x"83", x"84", x"84", x"83", x"82", x"82", x"83", x"84", x"84", x"84", x"84", 
        x"84", x"84", x"84", x"84", x"83", x"81", x"82", x"83", x"84", x"84", x"84", x"84", x"85", x"87", x"83", 
        x"7c", x"7a", x"80", x"86", x"84", x"86", x"85", x"84", x"85", x"85", x"84", x"87", x"81", x"87", x"75", 
        x"82", x"c6", x"de", x"d1", x"ce", x"d1", x"d5", x"d2", x"d0", x"d7", x"d8", x"c9", x"8d", x"33", x"16", 
        x"20", x"22", x"21", x"1e", x"1d", x"1e", x"1f", x"20", x"1f", x"1f", x"21", x"22", x"1e", x"16", x"0c", 
        x"05", x"03", x"04", x"05", x"09", x"09", x"04", x"03", x"01", x"04", x"05", x"05", x"09", x"09", x"0a", 
        x"15", x"24", x"31", x"34", x"32", x"33", x"38", x"38", x"35", x"39", x"3f", x"44", x"45", x"3a", x"33", 
        x"3a", x"a7", x"df", x"d3", x"d4", x"d2", x"d5", x"d9", x"cf", x"d1", x"d2", x"d0", x"d0", x"d1", x"d1", 
        x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", x"d2", x"d3", x"d0", x"d1", x"d4", x"d2", x"d1", x"d2", x"d3", 
        x"d5", x"d4", x"d4", x"d4", x"d4", x"d3", x"d2", x"d1", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d5", 
        x"d2", x"d2", x"d2", x"d1", x"d1", x"d2", x"cf", x"cf", x"dd", x"d4", x"d5", x"d5", x"d2", x"d3", x"d3", 
        x"d5", x"ed", x"f0", x"ee", x"f0", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ea", x"ee", x"f0", x"f0", x"ee", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"ee", x"ef", x"f1", x"f2", x"f0", x"e5", x"d1", x"c1", x"ba", x"c4", x"d5", x"e3", x"eb", 
        x"f2", x"f2", x"ef", x"ed", x"ef", x"f1", x"f1", x"ef", x"f1", x"f2", x"f1", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"ed", x"f0", x"f4", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f2", x"f2", x"eb", 
        x"d8", x"bf", x"b3", x"c1", x"d5", x"e7", x"ef", x"f1", x"f3", x"f4", x"f2", x"f3", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f1", x"f4", x"f2", x"ee", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f3", x"f2", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"ef", 
        x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"ed", 
        x"df", x"d8", x"de", x"e3", x"d8", x"b3", x"90", x"7f", x"81", x"88", x"88", x"8a", x"8c", x"8c", x"8c", 
        x"8a", x"8a", x"8b", x"8a", x"8a", x"8d", x"8e", x"8b", x"89", x"8a", x"8a", x"88", x"89", x"89", x"89", 
        x"88", x"88", x"8a", x"8c", x"89", x"8a", x"89", x"87", x"89", x"8a", x"88", x"89", x"89", x"8a", x"8a", 
        x"89", x"88", x"88", x"88", x"89", x"8b", x"8b", x"89", x"8a", x"8a", x"89", x"88", x"89", x"89", x"88", 
        x"88", x"88", x"87", x"85", x"86", x"87", x"88", x"89", x"89", x"88", x"88", x"89", x"8a", x"88", x"89", 
        x"8c", x"8b", x"88", x"87", x"86", x"85", x"88", x"8a", x"8a", x"88", x"84", x"82", x"84", x"83", x"86", 
        x"90", x"9d", x"a7", x"a7", x"aa", x"b8", x"ca", x"d8", x"de", x"d9", x"d8", x"d6", x"d6", x"d6", x"d7", 
        x"d7", x"d8", x"d8", x"d8", x"d7", x"d8", x"d8", x"d8", x"d7", x"d7", x"d9", x"d9", x"d8", x"d8", x"da", 
        x"da", x"d8", x"d7", x"d8", x"d7", x"d7", x"d8", x"d9", x"d7", x"d4", x"d4", x"d9", x"db", x"d8", x"d5", 
        x"d7", x"d7", x"cd", x"b4", x"9d", x"90", x"90", x"9a", x"9e", x"a4", x"a5", x"a5", x"a8", x"ab", x"ac", 
        x"ad", x"b0", x"a5", x"88", x"60", x"3c", x"19", x"17", x"1e", x"2a", x"42", x"5f", x"73", x"70", x"68", 
        x"88", x"85", x"84", x"84", x"83", x"82", x"82", x"80", x"80", x"81", x"83", x"82", x"81", x"80", x"7f", 
        x"81", x"81", x"7f", x"80", x"84", x"83", x"82", x"82", x"82", x"81", x"81", x"82", x"82", x"82", x"82", 
        x"83", x"83", x"83", x"83", x"83", x"82", x"82", x"82", x"82", x"83", x"83", x"83", x"84", x"82", x"82", 
        x"82", x"83", x"83", x"83", x"83", x"84", x"84", x"83", x"83", x"83", x"84", x"84", x"85", x"85", x"85", 
        x"84", x"84", x"84", x"84", x"83", x"82", x"82", x"83", x"84", x"84", x"84", x"84", x"83", x"82", x"85", 
        x"83", x"7b", x"7b", x"83", x"84", x"86", x"85", x"84", x"85", x"85", x"84", x"85", x"87", x"83", x"85", 
        x"c0", x"db", x"d4", x"d5", x"d3", x"d0", x"ce", x"d2", x"db", x"ca", x"90", x"52", x"26", x"1a", x"1d", 
        x"1f", x"1e", x"1e", x"1e", x"1e", x"1e", x"1f", x"20", x"20", x"1f", x"20", x"19", x"0f", x"06", x"03", 
        x"04", x"07", x"09", x"09", x"0c", x"0b", x"06", x"04", x"04", x"03", x"05", x"06", x"08", x"11", x"1f", 
        x"2c", x"33", x"35", x"33", x"35", x"34", x"34", x"39", x"3e", x"41", x"41", x"3d", x"3c", x"38", x"35", 
        x"38", x"a4", x"de", x"d4", x"d5", x"d4", x"d7", x"d9", x"cf", x"d0", x"d2", x"d0", x"d0", x"d2", x"d2", 
        x"d2", x"d1", x"d1", x"d2", x"d2", x"d1", x"d2", x"d3", x"d0", x"d1", x"d3", x"d2", x"d2", x"d2", x"d1", 
        x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d4", 
        x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"cf", x"cf", x"dc", x"d3", x"d5", x"d4", x"d3", x"d3", x"d3", 
        x"d5", x"ed", x"ef", x"ed", x"f0", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"f0", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ea", x"ee", x"f0", x"f0", x"ee", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f1", x"f2", x"f1", x"f1", x"f1", x"eb", x"e1", x"d3", x"ca", x"c4", x"c6", 
        x"d3", x"de", x"e9", x"f0", x"f2", x"f0", x"ee", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"ed", x"ef", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f0", x"f3", 
        x"f2", x"ed", x"dd", x"cb", x"be", x"be", x"c9", x"d7", x"e6", x"ef", x"f1", x"f0", x"ee", x"f0", x"f2", 
        x"f3", x"f2", x"f1", x"ee", x"f1", x"f2", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"ef", 
        x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"ee", x"ef", 
        x"ef", x"eb", x"e5", x"de", x"da", x"dc", x"d4", x"bb", x"9c", x"84", x"81", x"84", x"89", x"8e", x"8e", 
        x"8c", x"8b", x"8d", x"8c", x"8b", x"8b", x"8b", x"89", x"8a", x"8b", x"8b", x"8a", x"89", x"8b", x"8b", 
        x"88", x"88", x"8c", x"8d", x"8a", x"89", x"88", x"87", x"89", x"8b", x"8a", x"8a", x"8a", x"8a", x"8a", 
        x"89", x"88", x"88", x"88", x"87", x"88", x"8a", x"8b", x"89", x"89", x"88", x"87", x"89", x"89", x"88", 
        x"87", x"8a", x"8b", x"88", x"87", x"88", x"88", x"87", x"86", x"87", x"8b", x"8a", x"89", x"86", x"88", 
        x"8b", x"87", x"8a", x"8a", x"88", x"87", x"85", x"83", x"84", x"89", x"87", x"87", x"93", x"9d", x"a3", 
        x"a9", x"b2", x"bf", x"cc", x"d3", x"da", x"dd", x"da", x"d8", x"da", x"d6", x"d5", x"d8", x"d9", x"d8", 
        x"d7", x"d9", x"d8", x"d7", x"d7", x"d8", x"d9", x"d9", x"d5", x"d6", x"d8", x"d8", x"d8", x"d7", x"d7", 
        x"d7", x"d7", x"d7", x"d8", x"d9", x"d6", x"d5", x"d6", x"d8", x"db", x"da", x"da", x"d7", x"ce", x"c2", 
        x"b3", x"a4", x"9a", x"97", x"99", x"9d", x"a1", x"a1", x"a2", x"a7", x"ad", x"af", x"a9", x"a0", x"8d", 
        x"74", x"59", x"3c", x"21", x"22", x"2e", x"38", x"4e", x"63", x"6b", x"6b", x"66", x"5f", x"53", x"4d", 
        x"86", x"85", x"85", x"84", x"84", x"83", x"83", x"82", x"82", x"83", x"83", x"83", x"82", x"82", x"81", 
        x"83", x"83", x"81", x"82", x"84", x"84", x"83", x"83", x"82", x"81", x"81", x"82", x"83", x"83", x"83", 
        x"83", x"83", x"83", x"83", x"83", x"83", x"85", x"84", x"83", x"83", x"83", x"83", x"83", x"82", x"82", 
        x"82", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"84", x"84", x"83", x"83", x"84", x"85", x"85", 
        x"85", x"84", x"84", x"84", x"83", x"82", x"83", x"84", x"85", x"84", x"84", x"84", x"83", x"7f", x"83", 
        x"86", x"83", x"81", x"83", x"84", x"87", x"86", x"84", x"84", x"86", x"86", x"86", x"88", x"83", x"82", 
        x"c3", x"d7", x"d1", x"d6", x"d2", x"ce", x"d1", x"d7", x"bb", x"70", x"2b", x"15", x"1a", x"1b", x"16", 
        x"19", x"1b", x"19", x"1c", x"1b", x"1c", x"1f", x"21", x"1f", x"1b", x"12", x"09", x"03", x"03", x"07", 
        x"0a", x"0b", x"0d", x"0d", x"0c", x"0c", x"08", x"05", x"04", x"05", x"04", x"09", x"16", x"28", x"33", 
        x"33", x"32", x"36", x"38", x"36", x"37", x"3e", x"46", x"46", x"3f", x"3a", x"37", x"3a", x"3a", x"37", 
        x"37", x"9f", x"dd", x"d5", x"d8", x"d7", x"d9", x"d9", x"ce", x"d0", x"d1", x"d0", x"d0", x"d2", x"d2", 
        x"d2", x"d0", x"d0", x"d2", x"d1", x"cf", x"d1", x"d3", x"d0", x"d1", x"d2", x"d1", x"d2", x"d2", x"d1", 
        x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d4", 
        x"d3", x"d2", x"d1", x"d0", x"d0", x"d0", x"d0", x"cf", x"dc", x"d3", x"d4", x"d3", x"d3", x"d3", x"d3", 
        x"d6", x"ec", x"ee", x"ec", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ea", x"ee", x"f0", x"f0", x"ee", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"ee", x"f1", x"f4", x"f0", x"df", x"d1", 
        x"c7", x"c1", x"c5", x"d2", x"e0", x"eb", x"f1", x"f2", x"f1", x"f0", x"ee", x"ee", x"ef", x"f0", x"ef", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"ed", x"ee", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f0", x"f3", x"f1", x"ee", 
        x"ee", x"f1", x"f4", x"f3", x"eb", x"d5", x"bd", x"b6", x"c0", x"cf", x"dd", x"e9", x"ef", x"f1", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"f1", x"f2", x"ef", x"f0", x"f2", x"f3", x"f2", x"f1", x"f0", x"f0", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"ef", 
        x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"ee", x"f1", 
        x"f1", x"ee", x"f0", x"ef", x"e6", x"db", x"dd", x"e0", x"d6", x"bc", x"9c", x"84", x"7d", x"83", x"89", 
        x"8c", x"8d", x"8c", x"8c", x"8c", x"8d", x"8b", x"8a", x"8b", x"8b", x"89", x"8b", x"8a", x"8c", x"8a", 
        x"88", x"8a", x"8b", x"8a", x"8c", x"8b", x"89", x"88", x"88", x"89", x"8a", x"89", x"89", x"8a", x"8b", 
        x"8a", x"89", x"89", x"88", x"86", x"85", x"88", x"89", x"88", x"89", x"89", x"88", x"8a", x"89", x"87", 
        x"86", x"89", x"8b", x"89", x"87", x"89", x"8a", x"89", x"88", x"8a", x"86", x"89", x"8b", x"8a", x"8b", 
        x"8d", x"88", x"88", x"85", x"83", x"84", x"84", x"86", x"8b", x"94", x"9b", x"a3", x"aa", x"b2", x"be", 
        x"cd", x"d9", x"e0", x"dd", x"d7", x"d6", x"d8", x"da", x"d8", x"d7", x"d6", x"d8", x"d9", x"d8", x"d8", 
        x"da", x"da", x"d9", x"d7", x"d6", x"d7", x"d8", x"d9", x"d6", x"d6", x"d8", x"d8", x"d8", x"d7", x"d7", 
        x"d8", x"d9", x"d9", x"d8", x"d7", x"d7", x"d8", x"da", x"da", x"d6", x"ce", x"c0", x"af", x"9f", x"96", 
        x"96", x"99", x"9f", x"a4", x"a6", x"a5", x"a5", x"a9", x"ac", x"ad", x"a6", x"8f", x"6a", x"4d", x"28", 
        x"15", x"1a", x"2b", x"3b", x"54", x"6a", x"70", x"6e", x"68", x"5f", x"55", x"4e", x"48", x"49", x"47", 
        x"82", x"84", x"85", x"84", x"84", x"84", x"83", x"82", x"81", x"81", x"81", x"81", x"81", x"81", x"83", 
        x"84", x"84", x"83", x"83", x"84", x"84", x"84", x"83", x"82", x"83", x"83", x"82", x"83", x"84", x"83", 
        x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"82", x"83", x"83", x"84", x"85", x"82", x"82", 
        x"82", x"83", x"83", x"83", x"82", x"81", x"81", x"83", x"84", x"83", x"82", x"81", x"83", x"85", x"85", 
        x"85", x"84", x"84", x"84", x"84", x"84", x"83", x"84", x"84", x"84", x"84", x"85", x"86", x"83", x"82", 
        x"85", x"86", x"87", x"88", x"85", x"87", x"87", x"84", x"83", x"86", x"86", x"89", x"87", x"85", x"80", 
        x"c0", x"dc", x"ce", x"d3", x"cf", x"d8", x"d0", x"86", x"3b", x"19", x"1a", x"1c", x"19", x"19", x"1d", 
        x"1d", x"19", x"18", x"18", x"17", x"18", x"1a", x"19", x"12", x"0b", x"03", x"02", x"04", x"09", x"0d", 
        x"0d", x"0b", x"0e", x"0d", x"0b", x"0b", x"09", x"03", x"05", x"09", x"12", x"23", x"32", x"35", x"33", 
        x"34", x"33", x"32", x"38", x"42", x"4b", x"4a", x"43", x"3b", x"37", x"37", x"3a", x"3c", x"38", x"37", 
        x"3a", x"a4", x"e0", x"d5", x"d5", x"d5", x"d9", x"d9", x"cf", x"d0", x"d2", x"d0", x"d0", x"d2", x"d1", 
        x"d2", x"d0", x"cf", x"d0", x"d0", x"cf", x"d1", x"d3", x"d1", x"d0", x"d0", x"d0", x"d2", x"d1", x"d0", 
        x"d5", x"d5", x"d5", x"d4", x"d4", x"d4", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d4", x"d5", 
        x"d5", x"d3", x"d2", x"d1", x"d1", x"cf", x"d0", x"ce", x"db", x"d3", x"d4", x"d2", x"d3", x"d3", x"d3", 
        x"d5", x"ec", x"ee", x"ec", x"f0", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"ef", x"ef", 
        x"ee", x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"ef", x"ee", 
        x"ee", x"ef", x"ee", x"ee", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ea", x"ee", x"f0", x"f0", x"ee", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f2", x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", 
        x"ef", x"e4", x"d8", x"cd", x"c0", x"ba", x"c0", x"da", x"ea", x"f4", x"f6", x"f1", x"ef", x"f1", x"ef", 
        x"ee", x"ee", x"ee", x"ed", x"ed", x"ed", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f0", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"ef", x"f1", x"f2", x"ed", x"ed", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f2", x"f0", x"ef", x"f3", x"f3", x"f0", x"e8", x"d5", x"c1", x"b6", x"bc", x"cc", x"e0", x"ef", 
        x"f2", x"f1", x"f0", x"f1", x"ee", x"ef", x"f0", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"ef", 
        x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", 
        x"f1", x"f2", x"f2", x"f0", x"ef", x"ed", x"eb", x"e2", x"d8", x"d6", x"d5", x"ca", x"b4", x"94", x"7a", 
        x"79", x"8a", x"90", x"8f", x"8a", x"89", x"8b", x"89", x"8c", x"8d", x"8b", x"8e", x"8e", x"8c", x"8a", 
        x"8a", x"8d", x"8b", x"88", x"8a", x"88", x"88", x"89", x"8a", x"8b", x"8c", x"89", x"88", x"89", x"8b", 
        x"8b", x"8a", x"8a", x"8a", x"88", x"87", x"89", x"89", x"89", x"8b", x"8b", x"8a", x"8b", x"8a", x"87", 
        x"86", x"87", x"8a", x"89", x"88", x"8a", x"8b", x"8b", x"8b", x"8c", x"89", x"89", x"8c", x"8b", x"89", 
        x"86", x"7f", x"80", x"86", x"8f", x"94", x"94", x"96", x"9f", x"ad", x"bf", x"cd", x"d3", x"d7", x"dd", 
        x"da", x"d7", x"d5", x"d5", x"d7", x"d7", x"d7", x"d8", x"d8", x"d9", x"d8", x"d8", x"d7", x"d6", x"d7", 
        x"da", x"da", x"d9", x"d7", x"d6", x"d6", x"d6", x"d7", x"d6", x"d6", x"d7", x"d8", x"d9", x"da", x"da", 
        x"d9", x"d9", x"da", x"dc", x"de", x"dd", x"d7", x"c8", x"b3", x"a3", x"9c", x"9a", x"99", x"9c", x"a0", 
        x"a2", x"a2", x"a2", x"aa", x"b5", x"b6", x"ad", x"9a", x"7a", x"50", x"34", x"1d", x"11", x"1d", x"37", 
        x"4b", x"61", x"6a", x"66", x"60", x"5a", x"55", x"4e", x"4b", x"4b", x"49", x"43", x"42", x"36", x"2d", 
        x"82", x"85", x"85", x"83", x"83", x"83", x"82", x"83", x"83", x"83", x"82", x"83", x"83", x"83", x"83", 
        x"82", x"83", x"84", x"83", x"83", x"82", x"84", x"84", x"83", x"84", x"84", x"83", x"84", x"85", x"83", 
        x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"82", x"82", x"83", x"83", x"85", x"85", x"83", x"82", 
        x"82", x"83", x"83", x"83", x"82", x"82", x"82", x"82", x"83", x"83", x"82", x"82", x"84", x"85", x"85", 
        x"85", x"85", x"85", x"85", x"85", x"85", x"84", x"84", x"83", x"84", x"85", x"85", x"85", x"83", x"86", 
        x"87", x"85", x"84", x"87", x"85", x"88", x"87", x"84", x"84", x"86", x"87", x"85", x"86", x"84", x"7e", 
        x"c0", x"d6", x"cf", x"d7", x"d1", x"b2", x"69", x"2b", x"19", x"1e", x"1e", x"1c", x"1c", x"1c", x"1f", 
        x"1d", x"1a", x"1b", x"1b", x"18", x"14", x"10", x"0b", x"05", x"03", x"04", x"07", x"08", x"09", x"0a", 
        x"0b", x"0c", x"0c", x"0d", x"0a", x"09", x"06", x"07", x"12", x"20", x"2d", x"37", x"35", x"33", x"35", 
        x"39", x"3e", x"45", x"4b", x"4c", x"46", x"3c", x"37", x"37", x"38", x"38", x"39", x"38", x"39", x"3a", 
        x"3b", x"a7", x"e3", x"d5", x"d3", x"d3", x"d9", x"d9", x"cf", x"d1", x"d2", x"d0", x"d0", x"d1", x"d1", 
        x"d1", x"d2", x"d0", x"d0", x"d0", x"d1", x"d2", x"d2", x"d0", x"d0", x"d0", x"cf", x"d3", x"d2", x"cf", 
        x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d4", 
        x"d5", x"d4", x"d1", x"d1", x"d1", x"cf", x"d0", x"ce", x"db", x"d3", x"d4", x"d2", x"d3", x"d4", x"d2", 
        x"d4", x"ec", x"ef", x"ed", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ea", x"ee", x"f0", x"f0", x"ee", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f2", x"f3", x"f3", x"ee", x"e1", x"d1", x"c7", x"be", x"be", x"c8", x"d9", x"e9", x"ee", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ed", x"ed", x"ec", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"ed", x"ed", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f3", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f0", x"ef", x"f1", x"f2", x"ec", x"dd", x"ce", x"be", x"bc", x"c6", 
        x"da", x"e8", x"ef", x"f4", x"f0", x"ef", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f2", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"ef", 
        x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ed", 
        x"ee", x"f2", x"f2", x"ef", x"ee", x"ed", x"ef", x"ef", x"ea", x"df", x"d6", x"d4", x"d5", x"cb", x"b3", 
        x"95", x"82", x"81", x"89", x"8a", x"88", x"8e", x"8a", x"8c", x"8d", x"8a", x"8e", x"8d", x"8b", x"8b", 
        x"8c", x"8c", x"8b", x"8a", x"8b", x"89", x"89", x"8a", x"8a", x"89", x"8b", x"89", x"89", x"8a", x"8b", 
        x"8b", x"8a", x"8a", x"8a", x"8a", x"8a", x"8a", x"89", x"89", x"8b", x"8b", x"89", x"8a", x"89", x"89", 
        x"88", x"89", x"8a", x"8b", x"8b", x"8a", x"89", x"8a", x"8a", x"8b", x"89", x"85", x"86", x"85", x"82", 
        x"86", x"8d", x"96", x"99", x"9b", x"a4", x"b3", x"c0", x"c9", x"d1", x"db", x"de", x"db", x"d9", x"d9", 
        x"d7", x"d7", x"d6", x"d6", x"da", x"d8", x"d7", x"d7", x"d7", x"d9", x"d9", x"d8", x"d8", x"d8", x"d7", 
        x"d7", x"d9", x"d9", x"d8", x"d7", x"d7", x"d7", x"d8", x"da", x"d8", x"d6", x"d7", x"d7", x"d8", x"d7", 
        x"d9", x"da", x"d5", x"c8", x"b9", x"af", x"a9", x"a2", x"9b", x"9b", x"a0", x"a6", x"a7", x"a7", x"a6", 
        x"a9", x"ac", x"aa", x"a0", x"8e", x"6b", x"48", x"34", x"1f", x"0a", x"04", x"06", x"26", x"54", x"5a", 
        x"5d", x"5e", x"57", x"4e", x"4a", x"44", x"45", x"42", x"3f", x"3d", x"38", x"36", x"3a", x"51", x"6b", 
        x"84", x"87", x"85", x"81", x"80", x"82", x"82", x"81", x"82", x"83", x"84", x"84", x"83", x"82", x"81", 
        x"81", x"82", x"84", x"83", x"81", x"80", x"83", x"85", x"84", x"85", x"85", x"84", x"85", x"86", x"83", 
        x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"83", x"82", x"82", 
        x"82", x"83", x"82", x"83", x"83", x"84", x"84", x"83", x"82", x"82", x"83", x"84", x"84", x"84", x"85", 
        x"85", x"85", x"85", x"86", x"87", x"86", x"84", x"83", x"82", x"83", x"84", x"85", x"84", x"85", x"85", 
        x"85", x"85", x"84", x"84", x"85", x"88", x"87", x"84", x"83", x"86", x"87", x"87", x"85", x"83", x"7e", 
        x"ba", x"d7", x"dc", x"d2", x"8e", x"3c", x"1c", x"1d", x"20", x"20", x"20", x"1e", x"1d", x"1d", x"1c", 
        x"1c", x"1d", x"1b", x"1d", x"17", x"0f", x"06", x"02", x"04", x"07", x"08", x"0a", x"0c", x"0b", x"0a", 
        x"0a", x"0b", x"0b", x"0d", x"0a", x"06", x"06", x"0e", x"25", x"35", x"39", x"37", x"32", x"31", x"37", 
        x"40", x"51", x"58", x"48", x"3e", x"39", x"38", x"37", x"39", x"3b", x"37", x"38", x"3b", x"3a", x"3b", 
        x"3a", x"a4", x"e2", x"d6", x"d4", x"d5", x"d9", x"d9", x"d0", x"d2", x"d2", x"d0", x"d0", x"d1", x"d0", 
        x"d1", x"d4", x"d3", x"d1", x"d1", x"d4", x"d3", x"d2", x"d0", x"cf", x"cf", x"d0", x"d4", x"d2", x"cf", 
        x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", 
        x"d5", x"d3", x"d0", x"d1", x"d0", x"cd", x"d0", x"ce", x"db", x"d3", x"d4", x"d2", x"d3", x"d4", x"d2", 
        x"d4", x"eb", x"ef", x"ee", x"ef", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"f0", x"f1", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f2", x"f1", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"f1", x"ef", x"ef", x"ee", 
        x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ea", x"ee", x"f0", x"f0", x"ee", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f3", x"f4", x"f2", x"f0", 
        x"f0", x"f1", x"ef", x"f0", x"f4", x"f2", x"ea", x"e4", x"dc", x"cc", x"b7", x"ad", x"be", x"d9", x"ed", 
        x"f1", x"f1", x"f1", x"ef", x"ee", x"ed", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f0", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"f0", x"f2", x"f2", x"ed", x"ed", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"f2", 
        x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"eb", x"dc", x"c9", 
        x"b3", x"af", x"c8", x"e7", x"f3", x"f4", x"f2", x"ef", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", 
        x"ef", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"ef", 
        x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"f1", x"f1", x"ee", x"f1", x"f0", x"ec", x"ee", x"ee", x"e3", x"d5", x"cf", x"d0", 
        x"d5", x"c4", x"9e", x"7d", x"75", x"84", x"8e", x"8a", x"8c", x"8d", x"8a", x"8e", x"8b", x"8b", x"8d", 
        x"8d", x"8a", x"8a", x"8e", x"8b", x"88", x"89", x"8c", x"8b", x"8a", x"8c", x"8b", x"8a", x"8b", x"8c", 
        x"8a", x"89", x"89", x"87", x"89", x"8b", x"89", x"87", x"87", x"88", x"89", x"8b", x"8b", x"8a", x"8a", 
        x"89", x"88", x"89", x"8a", x"8b", x"89", x"88", x"8a", x"8b", x"89", x"81", x"7c", x"86", x"97", x"9b", 
        x"98", x"94", x"a2", x"b4", x"c5", x"d1", x"d7", x"db", x"dc", x"dc", x"db", x"d7", x"d7", x"d8", x"d9", 
        x"d9", x"d8", x"d6", x"d8", x"da", x"d8", x"d8", x"d8", x"d7", x"d9", x"da", x"d9", x"d7", x"d8", x"da", 
        x"da", x"d9", x"d9", x"d9", x"d9", x"d9", x"d9", x"d9", x"d8", x"d7", x"d6", x"d8", x"dc", x"de", x"dd", 
        x"cd", x"b6", x"9c", x"8d", x"8f", x"9a", x"9e", x"a1", x"a3", x"a3", x"a1", x"a5", x"af", x"b6", x"b5", 
        x"a8", x"8b", x"5d", x"37", x"21", x"12", x"06", x"03", x"04", x"06", x"07", x"07", x"2f", x"66", x"53", 
        x"43", x"3f", x"3f", x"3d", x"3d", x"3d", x"3a", x"2e", x"26", x"2f", x"50", x"7c", x"a1", x"c5", x"d7", 
        x"85", x"86", x"86", x"86", x"85", x"85", x"84", x"81", x"81", x"83", x"84", x"83", x"82", x"82", x"83", 
        x"83", x"84", x"83", x"83", x"83", x"82", x"83", x"85", x"83", x"83", x"84", x"84", x"84", x"84", x"83", 
        x"83", x"82", x"82", x"82", x"83", x"83", x"82", x"83", x"84", x"85", x"84", x"83", x"82", x"82", x"82", 
        x"84", x"84", x"84", x"84", x"83", x"84", x"86", x"83", x"84", x"84", x"84", x"86", x"86", x"86", x"86", 
        x"87", x"85", x"84", x"85", x"86", x"86", x"87", x"86", x"85", x"84", x"85", x"86", x"84", x"87", x"88", 
        x"87", x"86", x"87", x"87", x"87", x"84", x"86", x"86", x"85", x"87", x"88", x"88", x"89", x"83", x"81", 
        x"bd", x"d4", x"a7", x"53", x"23", x"1a", x"1d", x"1b", x"1c", x"1b", x"19", x"1a", x"1c", x"1c", x"1c", 
        x"1e", x"21", x"19", x"0f", x"06", x"05", x"02", x"02", x"09", x"0c", x"0c", x"0d", x"0d", x"0d", x"0a", 
        x"0a", x"0b", x"0a", x"08", x"0f", x"1c", x"15", x"14", x"2c", x"35", x"35", x"35", x"33", x"3b", x"4b", 
        x"51", x"4e", x"42", x"3a", x"3d", x"3e", x"3c", x"3b", x"38", x"38", x"39", x"3c", x"3a", x"39", x"3a", 
        x"39", x"9e", x"df", x"d3", x"d2", x"d4", x"d8", x"da", x"d0", x"d1", x"d2", x"d1", x"d0", x"d0", x"d0", 
        x"d0", x"d3", x"d3", x"d0", x"d1", x"d5", x"d1", x"cf", x"d0", x"d0", x"d0", x"d1", x"d3", x"d3", x"d2", 
        x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", x"d3", x"d3", x"d3", x"d1", x"d2", 
        x"d5", x"cf", x"cf", x"d3", x"d3", x"d0", x"d0", x"cc", x"d9", x"d3", x"d4", x"d1", x"d1", x"d7", x"d4", 
        x"d2", x"e3", x"ea", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"ee", x"ee", x"ef", x"ee", x"ed", x"ee", x"ef", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", 
        x"ef", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"eb", x"ed", x"f1", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ed", x"f1", x"f1", x"f0", x"f2", x"f1", x"f0", x"f1", x"f2", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f1", x"f0", x"f0", x"f3", x"f2", x"ef", x"e9", x"dc", x"cb", x"bc", x"b4", 
        x"bf", x"d4", x"e7", x"f0", x"f2", x"f0", x"f0", x"f1", x"f0", x"ee", x"ee", x"ef", x"f1", x"f2", x"f3", 
        x"f3", x"f0", x"ee", x"f0", x"f1", x"f1", x"f2", x"f0", x"f0", x"f1", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f1", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"ed", x"ef", x"f1", x"f2", x"f1", x"f3", x"f3", x"f4", 
        x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f0", x"ec", 
        x"e3", x"d9", x"c3", x"b6", x"bc", x"d2", x"e8", x"ee", x"f1", x"f3", x"f2", x"f1", x"f2", x"f3", x"f1", 
        x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f0", 
        x"ec", x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"ee", x"ee", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"e8", x"d9", 
        x"cf", x"d2", x"d8", x"ca", x"a8", x"89", x"7c", x"80", x"87", x"8a", x"8e", x"90", x"8d", x"8c", x"8c", 
        x"8c", x"8a", x"8b", x"8c", x"88", x"8e", x"8d", x"8b", x"8e", x"8e", x"8e", x"8d", x"8b", x"8a", x"8c", 
        x"8b", x"8a", x"89", x"8a", x"8a", x"8a", x"8a", x"8b", x"8b", x"8b", x"8a", x"8a", x"8a", x"8a", x"8a", 
        x"89", x"89", x"89", x"89", x"89", x"8a", x"8a", x"87", x"85", x"8b", x"98", x"9e", x"a0", x"a1", x"ad", 
        x"bb", x"cb", x"d3", x"d6", x"d8", x"d8", x"d7", x"d7", x"d8", x"d7", x"d9", x"d8", x"d8", x"da", x"d9", 
        x"d8", x"d9", x"d8", x"d8", x"d8", x"d9", x"da", x"da", x"da", x"dc", x"dd", x"dd", x"db", x"da", x"da", 
        x"db", x"da", x"db", x"da", x"db", x"d8", x"d8", x"d8", x"db", x"dc", x"dd", x"d3", x"c7", x"b1", x"9f", 
        x"9d", x"9f", x"a0", x"a3", x"a3", x"a1", x"9f", x"a2", x"a8", x"ad", x"b0", x"aa", x"96", x"74", x"49", 
        x"2a", x"1c", x"0f", x"0a", x"0b", x"12", x"20", x"35", x"26", x"08", x"07", x"08", x"2d", x"6b", x"57", 
        x"42", x"38", x"31", x"31", x"34", x"37", x"46", x"6d", x"96", x"b5", x"ce", x"dd", x"e4", x"e4", x"e2", 
        x"86", x"86", x"86", x"85", x"85", x"85", x"86", x"84", x"84", x"84", x"84", x"83", x"81", x"81", x"83", 
        x"84", x"84", x"83", x"83", x"83", x"83", x"83", x"84", x"82", x"82", x"84", x"84", x"83", x"83", x"82", 
        x"83", x"82", x"83", x"83", x"83", x"83", x"81", x"83", x"85", x"86", x"85", x"83", x"82", x"84", x"85", 
        x"86", x"85", x"85", x"84", x"83", x"85", x"87", x"84", x"84", x"84", x"84", x"86", x"85", x"84", x"85", 
        x"86", x"85", x"84", x"85", x"86", x"85", x"86", x"87", x"87", x"86", x"86", x"87", x"86", x"86", x"86", 
        x"88", x"89", x"88", x"86", x"87", x"84", x"87", x"87", x"85", x"87", x"86", x"86", x"88", x"81", x"88", 
        x"a8", x"81", x"37", x"1a", x"17", x"1c", x"1d", x"16", x"1a", x"1b", x"19", x"19", x"1c", x"1d", x"1b", 
        x"1b", x"1a", x"0f", x"03", x"02", x"05", x"05", x"06", x"0c", x"0f", x"0f", x"0a", x"0a", x"0d", x"0b", 
        x"0a", x"0d", x"10", x"17", x"29", x"37", x"22", x"17", x"2c", x"32", x"2f", x"39", x"49", x"51", x"50", 
        x"44", x"3d", x"39", x"3b", x"3f", x"3f", x"3b", x"3d", x"3d", x"3b", x"3e", x"3e", x"3b", x"3b", x"3c", 
        x"3a", x"9b", x"df", x"d6", x"d4", x"d6", x"d8", x"da", x"d0", x"d0", x"d2", x"d1", x"d0", x"d0", x"d0", 
        x"cf", x"d2", x"d2", x"cf", x"d1", x"d5", x"d2", x"d1", x"d2", x"d0", x"ce", x"d1", x"d2", x"d2", x"d2", 
        x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d2", x"d2", x"d1", x"d5", 
        x"d6", x"cf", x"cf", x"cf", x"d1", x"d4", x"d0", x"cc", x"dc", x"d2", x"d1", x"d4", x"d6", x"d9", x"c1", 
        x"9a", x"9f", x"b9", x"cd", x"da", x"e6", x"ec", x"ed", x"ee", x"ed", x"ed", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ed", x"ee", x"ee", x"ef", x"ef", x"ec", x"ea", x"ec", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"eb", x"ec", x"f1", x"ef", x"ee", 
        x"ef", x"f0", x"ee", x"ee", x"f1", x"f0", x"f0", x"f2", x"f0", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f2", x"f2", x"ef", x"eb", x"df", 
        x"cd", x"b9", x"b3", x"c2", x"d7", x"e8", x"ed", x"f0", x"f2", x"f2", x"ef", x"ee", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"f0", x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"ed", x"f0", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f1", x"f0", x"e5", x"ce", x"b8", x"ae", x"c2", x"dd", x"eb", x"f0", x"f2", x"f0", x"ee", x"ef", 
        x"ef", x"f1", x"f0", x"ee", x"ef", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f1", 
        x"ec", x"f0", x"f1", x"ef", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", 
        x"ed", x"da", x"ce", x"d0", x"d9", x"d3", x"b3", x"8e", x"7b", x"7f", x"8b", x"8a", x"8c", x"8e", x"8b", 
        x"8b", x"91", x"91", x"8a", x"88", x"8e", x"8c", x"8b", x"8d", x"8b", x"8c", x"8c", x"8a", x"89", x"8c", 
        x"8c", x"8a", x"8a", x"8c", x"8c", x"8b", x"8b", x"8c", x"8c", x"8b", x"8a", x"8a", x"8b", x"8c", x"8c", 
        x"8b", x"8a", x"8a", x"89", x"8a", x"8c", x"8a", x"89", x"8c", x"9c", x"a5", x"b0", x"bf", x"cf", x"de", 
        x"de", x"db", x"da", x"d9", x"d8", x"d7", x"d7", x"d8", x"d9", x"d7", x"d8", x"d8", x"d7", x"da", x"d8", 
        x"d8", x"d8", x"d8", x"d9", x"d9", x"da", x"d8", x"d7", x"d8", x"db", x"d8", x"d8", x"da", x"db", x"db", 
        x"da", x"dc", x"db", x"da", x"dc", x"db", x"dd", x"dd", x"d8", x"c6", x"ae", x"9e", x"9b", x"9d", x"a0", 
        x"a5", x"a5", x"a4", x"a6", x"aa", x"ae", x"ae", x"ac", x"9f", x"8b", x"6c", x"3e", x"1e", x"0f", x"0b", 
        x"0c", x"0e", x"13", x"29", x"42", x"53", x"59", x"59", x"36", x"07", x"08", x"0a", x"2a", x"65", x"59", 
        x"44", x"37", x"34", x"4c", x"7b", x"a1", x"ca", x"df", x"e4", x"e3", x"e2", x"e2", x"e2", x"e2", x"e4", 
        x"87", x"86", x"85", x"85", x"85", x"85", x"86", x"85", x"84", x"84", x"84", x"84", x"83", x"81", x"83", 
        x"84", x"84", x"84", x"84", x"84", x"84", x"84", x"83", x"83", x"83", x"84", x"83", x"82", x"82", x"82", 
        x"83", x"83", x"83", x"84", x"84", x"84", x"82", x"84", x"87", x"86", x"85", x"83", x"84", x"86", x"87", 
        x"87", x"86", x"85", x"84", x"83", x"85", x"86", x"84", x"84", x"84", x"84", x"86", x"85", x"83", x"84", 
        x"85", x"85", x"84", x"85", x"85", x"83", x"85", x"87", x"87", x"86", x"86", x"87", x"86", x"86", x"86", 
        x"88", x"89", x"88", x"86", x"87", x"86", x"87", x"86", x"85", x"86", x"84", x"85", x"86", x"81", x"80", 
        x"85", x"6f", x"4f", x"36", x"28", x"26", x"20", x"16", x"17", x"17", x"19", x"1c", x"1a", x"1b", x"1a", 
        x"17", x"14", x"0a", x"03", x"04", x"03", x"04", x"07", x"09", x"0b", x"0d", x"0b", x"0e", x"10", x"0e", 
        x"11", x"1b", x"2d", x"31", x"35", x"34", x"2b", x"45", x"46", x"32", x"33", x"4c", x"58", x"4a", x"3f", 
        x"3c", x"3c", x"3c", x"3d", x"3f", x"3f", x"3b", x"3d", x"40", x"3f", x"3f", x"3f", x"3b", x"3c", x"3e", 
        x"3a", x"99", x"de", x"d5", x"d3", x"d3", x"d6", x"d9", x"d0", x"d0", x"d2", x"d1", x"d0", x"d0", x"d0", 
        x"cf", x"d1", x"d1", x"cf", x"d1", x"d5", x"d3", x"d3", x"d3", x"cf", x"cd", x"d1", x"d1", x"d1", x"d2", 
        x"d1", x"d2", x"d3", x"d1", x"d1", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d2", x"d1", x"d0", x"d3", 
        x"d4", x"d3", x"d5", x"d3", x"d3", x"d4", x"cf", x"cd", x"da", x"d7", x"d8", x"ce", x"bf", x"a5", x"9d", 
        x"b4", x"d0", x"c1", x"b2", x"a6", x"ac", x"bb", x"cb", x"dc", x"e7", x"ed", x"f1", x"f2", x"f1", x"ee", 
        x"ee", x"ed", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"eb", x"ec", x"f1", x"ef", x"ee", 
        x"ef", x"f0", x"ef", x"f0", x"f1", x"ef", x"f0", x"f2", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ee", x"ee", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f0", 
        x"f0", x"eb", x"dd", x"cb", x"c0", x"bc", x"c6", x"d2", x"e0", x"eb", x"ef", x"f0", x"f1", x"f0", x"f0", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f2", x"ed", x"ef", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f1", x"ec", x"e0", x"c8", x"b3", x"bb", x"cf", x"e1", x"eb", x"f2", x"f4", 
        x"f2", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f1", 
        x"ec", x"ef", x"f2", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ee", x"eb", x"e2", x"d3", x"cd", x"d7", x"d3", x"b3", x"93", x"87", x"85", x"8a", x"88", x"8c", 
        x"8f", x"8c", x"8c", x"90", x"8e", x"8e", x"8d", x"8c", x"8c", x"8a", x"8c", x"8c", x"8a", x"8a", x"8c", 
        x"8d", x"8c", x"8b", x"8d", x"8d", x"8c", x"8c", x"8c", x"8c", x"8b", x"8a", x"8a", x"8c", x"8d", x"8d", 
        x"8c", x"8a", x"89", x"88", x"8d", x"8f", x"89", x"85", x"84", x"a5", x"d5", x"da", x"df", x"de", x"dc", 
        x"db", x"da", x"d8", x"d8", x"d8", x"d8", x"d8", x"d8", x"d8", x"d8", x"d9", x"d8", x"d6", x"d9", x"d8", 
        x"d8", x"da", x"d9", x"d9", x"d9", x"d8", x"d7", x"d8", x"d8", x"d8", x"da", x"db", x"da", x"d9", x"da", 
        x"db", x"dc", x"db", x"db", x"d9", x"ca", x"b9", x"aa", x"9d", x"9c", x"a0", x"a2", x"a6", x"a7", x"a7", 
        x"aa", x"aa", x"a8", x"a9", x"a6", x"94", x"7c", x"59", x"31", x"1b", x"10", x"0b", x"0d", x"15", x"20", 
        x"33", x"49", x"53", x"55", x"57", x"54", x"4e", x"4b", x"2e", x"0b", x"0b", x"0a", x"26", x"5a", x"58", 
        x"68", x"8d", x"ae", x"cb", x"df", x"e5", x"e5", x"e5", x"e3", x"e1", x"e1", x"e2", x"e3", x"e6", x"e6", 
        x"87", x"87", x"86", x"86", x"86", x"85", x"85", x"84", x"82", x"82", x"83", x"85", x"85", x"83", x"83", 
        x"84", x"84", x"84", x"85", x"85", x"85", x"84", x"83", x"83", x"83", x"84", x"83", x"82", x"82", x"83", 
        x"83", x"83", x"83", x"84", x"86", x"86", x"84", x"85", x"86", x"85", x"84", x"85", x"86", x"86", x"86", 
        x"85", x"85", x"85", x"84", x"84", x"85", x"85", x"85", x"85", x"85", x"85", x"85", x"85", x"84", x"84", 
        x"85", x"85", x"84", x"84", x"85", x"84", x"84", x"86", x"86", x"86", x"86", x"85", x"85", x"87", x"88", 
        x"87", x"86", x"87", x"88", x"87", x"87", x"88", x"86", x"85", x"87", x"83", x"83", x"86", x"85", x"84", 
        x"86", x"91", x"94", x"91", x"85", x"71", x"56", x"3a", x"2a", x"1e", x"18", x"16", x"13", x"15", x"15", 
        x"13", x"12", x"0a", x"05", x"03", x"05", x"03", x"02", x"05", x"06", x"07", x"07", x"08", x"0a", x"15", 
        x"29", x"3e", x"47", x"3b", x"3a", x"39", x"3a", x"85", x"7e", x"3b", x"31", x"43", x"48", x"3c", x"3c", 
        x"40", x"41", x"41", x"3d", x"3d", x"41", x"3e", x"3b", x"3d", x"3f", x"40", x"3f", x"3c", x"3c", x"3d", 
        x"39", x"9a", x"df", x"d6", x"d1", x"d2", x"d6", x"db", x"d0", x"d0", x"d1", x"d1", x"d0", x"d0", x"d0", 
        x"d0", x"d1", x"d1", x"cf", x"d2", x"d4", x"d2", x"d2", x"d2", x"cf", x"ce", x"d2", x"d3", x"d1", x"d1", 
        x"d2", x"d3", x"d3", x"d2", x"d1", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d1", x"d1", x"d4", 
        x"d4", x"d1", x"d0", x"cc", x"cf", x"d2", x"d6", x"d3", x"e1", x"d6", x"be", x"9f", x"91", x"b2", x"cf", 
        x"db", x"f0", x"f3", x"ed", x"e5", x"cf", x"b7", x"a2", x"9c", x"aa", x"c1", x"d5", x"e0", x"e8", x"ef", 
        x"f1", x"ed", x"ea", x"ec", x"ef", x"ec", x"ed", x"ed", x"ee", x"ee", x"ed", x"ee", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ee", x"ef", x"f0", x"f0", 
        x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"eb", x"ec", x"f1", x"ef", x"ee", 
        x"ef", x"f0", x"f0", x"f1", x"f1", x"ee", x"f0", x"f2", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", 
        x"ee", x"ee", x"f2", x"f4", x"ee", x"e3", x"cc", x"bb", x"b4", x"bb", x"ce", x"e0", x"ea", x"ef", x"f3", 
        x"f3", x"f1", x"ef", x"f2", x"f3", x"f2", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ed", x"ef", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f1", x"f3", x"f1", x"f2", x"f5", x"f4", x"ee", x"d1", x"ba", x"b2", x"bd", x"d1", x"e1", 
        x"ee", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"ef", 
        x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", 
        x"eb", x"ef", x"f2", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ed", x"ef", x"f2", 
        x"f1", x"ef", x"ef", x"f1", x"f0", x"e5", x"d0", x"ca", x"d7", x"df", x"c5", x"9d", x"82", x"7f", x"84", 
        x"8c", x"90", x"8f", x"8d", x"8e", x"8d", x"8c", x"8b", x"8c", x"8e", x"8f", x"8d", x"8b", x"8b", x"8c", 
        x"8e", x"8e", x"8d", x"8d", x"8d", x"8c", x"8d", x"8d", x"8d", x"8d", x"8b", x"8a", x"8b", x"8c", x"8c", 
        x"8c", x"8b", x"8b", x"8e", x"91", x"90", x"8a", x"8a", x"88", x"af", x"e0", x"da", x"dd", x"dc", x"d9", 
        x"db", x"da", x"d9", x"d8", x"d9", x"d8", x"d8", x"d7", x"d7", x"d8", x"da", x"d8", x"d7", x"d9", x"d8", 
        x"d9", x"d9", x"d7", x"d7", x"d6", x"d6", x"d6", x"d7", x"d8", x"d9", x"d9", x"db", x"de", x"df", x"db", 
        x"d7", x"d5", x"cd", x"be", x"aa", x"9a", x"97", x"a0", x"a8", x"a7", x"a4", x"a3", x"ab", x"b1", x"af", 
        x"ae", x"a2", x"87", x"65", x"40", x"1e", x"0b", x"05", x"06", x"0f", x"1b", x"25", x"39", x"52", x"5f", 
        x"60", x"5b", x"52", x"4b", x"4a", x"48", x"45", x"40", x"2c", x"17", x"27", x"41", x"6b", x"a3", x"c7", 
        x"db", x"eb", x"eb", x"e4", x"e3", x"e1", x"e2", x"e5", x"e5", x"e5", x"e8", x"e7", x"e4", x"d8", x"c2", 
        x"86", x"87", x"87", x"87", x"86", x"85", x"83", x"84", x"83", x"82", x"82", x"84", x"83", x"82", x"83", 
        x"84", x"84", x"84", x"85", x"86", x"86", x"84", x"83", x"83", x"84", x"84", x"83", x"83", x"83", x"84", 
        x"83", x"83", x"83", x"84", x"86", x"86", x"86", x"85", x"84", x"84", x"84", x"85", x"86", x"85", x"84", 
        x"84", x"84", x"84", x"85", x"85", x"85", x"84", x"86", x"86", x"86", x"85", x"85", x"86", x"85", x"84", 
        x"85", x"85", x"84", x"83", x"85", x"86", x"85", x"85", x"85", x"86", x"86", x"85", x"86", x"87", x"87", 
        x"87", x"86", x"87", x"88", x"88", x"87", x"88", x"86", x"85", x"87", x"85", x"84", x"89", x"85", x"85", 
        x"85", x"82", x"84", x"86", x"89", x"8e", x"91", x"8a", x"7e", x"70", x"5b", x"47", x"36", x"25", x"18", 
        x"0f", x"0d", x"0b", x"0a", x"03", x"09", x"09", x"08", x"0a", x"07", x"04", x"05", x"08", x"17", x"2d", 
        x"3d", x"43", x"41", x"43", x"3e", x"36", x"2e", x"85", x"82", x"3b", x"2f", x"3b", x"43", x"3e", x"3f", 
        x"41", x"41", x"42", x"3d", x"3d", x"41", x"40", x"3d", x"3e", x"3f", x"40", x"40", x"3e", x"3e", x"3e", 
        x"39", x"99", x"de", x"d5", x"d2", x"d3", x"d5", x"d9", x"d0", x"cf", x"d1", x"d0", x"cf", x"cf", x"d0", 
        x"d1", x"d2", x"d1", x"d0", x"d2", x"d3", x"d1", x"d0", x"d0", x"cf", x"d0", x"d4", x"d4", x"d2", x"d2", 
        x"d3", x"d4", x"d4", x"d2", x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", x"d2", x"d3", x"d3", x"d3", x"d2", 
        x"d1", x"d3", x"d6", x"d2", x"d2", x"d2", x"d3", x"d6", x"cb", x"a4", x"93", x"ac", x"cb", x"d8", x"d1", 
        x"d6", x"ee", x"ed", x"ee", x"ee", x"ed", x"ee", x"ea", x"d9", x"c3", x"b2", x"ab", x"ac", x"b3", x"c1", 
        x"d3", x"e2", x"ed", x"f2", x"f3", x"f0", x"f0", x"ef", x"ee", x"ed", x"ed", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ee", x"ee", x"ef", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"eb", x"ec", x"f1", x"ef", x"ee", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"ef", x"f0", x"f2", x"ee", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"f2", x"f1", x"f0", x"ef", x"f0", x"f0", x"ee", x"ef", 
        x"f1", x"f1", x"ef", x"ed", x"ee", x"f2", x"f3", x"ef", x"e2", x"ce", x"be", x"b8", x"be", x"cb", x"db", 
        x"eb", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"ee", x"ee", x"f0", x"f3", x"f3", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"ed", x"ee", x"f2", x"f1", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f0", x"f2", x"f3", x"f1", x"ef", x"f0", x"f2", x"f4", x"f0", x"e3", x"ce", x"bc", x"bb", 
        x"c3", x"d4", x"e2", x"ee", x"f5", x"f4", x"f1", x"f2", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"eb", x"ee", x"f2", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"f0", 
        x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"e6", x"db", x"d6", x"d7", x"d6", x"ca", x"ad", x"91", 
        x"84", x"81", x"88", x"90", x"90", x"8f", x"8e", x"8d", x"8e", x"8f", x"8e", x"8c", x"8c", x"8c", x"8d", 
        x"8e", x"8f", x"8c", x"8c", x"8c", x"8c", x"8d", x"8e", x"8e", x"8e", x"8d", x"8d", x"8d", x"8c", x"8c", 
        x"8c", x"8d", x"8b", x"89", x"8b", x"8d", x"8a", x"8b", x"84", x"a7", x"e5", x"db", x"db", x"dd", x"dc", 
        x"dc", x"d8", x"d8", x"d8", x"d8", x"d8", x"d8", x"d9", x"d9", x"d9", x"da", x"d8", x"d7", x"da", x"d9", 
        x"da", x"db", x"da", x"d9", x"da", x"da", x"da", x"da", x"db", x"de", x"e0", x"e0", x"da", x"cd", x"bf", 
        x"b3", x"a7", x"a3", x"a2", x"a3", x"a5", x"a4", x"a5", x"ab", x"af", x"b2", x"af", x"ab", x"95", x"74", 
        x"59", x"3c", x"1d", x"0b", x"05", x"09", x"13", x"21", x"34", x"4a", x"58", x"5e", x"61", x"59", x"4f", 
        x"4c", x"4a", x"49", x"40", x"36", x"38", x"44", x"52", x"67", x"85", x"ad", x"cd", x"dc", x"e8", x"e5", 
        x"e4", x"e3", x"e1", x"e1", x"e7", x"e5", x"e6", x"e9", x"e5", x"dc", x"c8", x"a4", x"7f", x"59", x"36", 
        x"86", x"87", x"87", x"87", x"86", x"84", x"83", x"85", x"85", x"84", x"83", x"83", x"82", x"82", x"83", 
        x"84", x"85", x"85", x"86", x"86", x"87", x"85", x"83", x"84", x"84", x"84", x"83", x"84", x"84", x"84", 
        x"84", x"84", x"84", x"84", x"85", x"85", x"86", x"85", x"83", x"84", x"85", x"85", x"85", x"86", x"85", 
        x"85", x"84", x"85", x"86", x"86", x"85", x"84", x"86", x"85", x"85", x"85", x"85", x"87", x"86", x"84", 
        x"85", x"85", x"84", x"83", x"85", x"86", x"85", x"85", x"86", x"86", x"86", x"86", x"86", x"87", x"86", 
        x"87", x"87", x"87", x"88", x"88", x"87", x"88", x"87", x"85", x"87", x"86", x"86", x"8a", x"88", x"87", 
        x"89", x"88", x"87", x"85", x"84", x"84", x"87", x"8b", x"8d", x"91", x"90", x"8d", x"80", x"6e", x"5b", 
        x"48", x"38", x"22", x"0e", x"08", x"0a", x"0d", x"0f", x"0d", x"0c", x"11", x"1e", x"28", x"2f", x"35", 
        x"38", x"37", x"37", x"3f", x"3f", x"44", x"36", x"80", x"7f", x"3b", x"31", x"3e", x"45", x"3e", x"3a", 
        x"3e", x"41", x"41", x"3f", x"3f", x"3f", x"40", x"40", x"3f", x"3e", x"3e", x"3e", x"3e", x"3f", x"3f", 
        x"3a", x"99", x"de", x"d6", x"d4", x"d5", x"d7", x"d9", x"cf", x"cf", x"d1", x"d0", x"cf", x"cf", x"d0", 
        x"d1", x"d2", x"d0", x"d1", x"d2", x"d2", x"d1", x"cf", x"d0", x"d0", x"d1", x"d4", x"d3", x"d1", x"d2", 
        x"d3", x"d4", x"d4", x"d2", x"d1", x"d1", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", x"d3", x"d3", 
        x"d2", x"d2", x"d3", x"d1", x"d5", x"d5", x"c9", x"ae", x"a1", x"a6", x"c6", x"d6", x"d5", x"d3", x"d2", 
        x"d4", x"ee", x"f1", x"ec", x"ec", x"ed", x"ec", x"ed", x"f1", x"f2", x"ec", x"e0", x"ce", x"bc", x"b7", 
        x"b4", x"b6", x"c1", x"d0", x"db", x"e7", x"ef", x"f2", x"f0", x"eb", x"ec", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"eb", x"ec", x"f1", x"ef", x"ee", 
        x"ef", x"f0", x"ef", x"ef", x"f1", x"f0", x"f0", x"f2", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"f2", x"f2", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"ed", x"df", x"c9", x"c0", x"bf", 
        x"c3", x"ce", x"dd", x"eb", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"ee", x"ee", x"f3", x"f2", x"f3", x"f4", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", 
        x"f2", x"f4", x"f5", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f4", x"f3", x"f3", x"ec", x"da", 
        x"c5", x"bc", x"c0", x"cb", x"dd", x"ec", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"eb", x"ee", x"f2", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"ee", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"ea", x"db", x"d5", x"db", x"dc", x"cb", 
        x"ae", x"93", x"83", x"7f", x"8a", x"8c", x"8f", x"90", x"8f", x"8e", x"8b", x"8c", x"8e", x"8d", x"8d", 
        x"8f", x"8f", x"8c", x"8c", x"8c", x"8c", x"8c", x"8e", x"8e", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", 
        x"8d", x"8d", x"8d", x"8c", x"8a", x"8c", x"8a", x"8d", x"85", x"a2", x"e2", x"dc", x"dc", x"db", x"da", 
        x"d9", x"d6", x"d8", x"d8", x"d8", x"d9", x"d9", x"da", x"db", x"da", x"db", x"da", x"d9", x"dc", x"da", 
        x"db", x"dc", x"da", x"d7", x"d7", x"da", x"dd", x"dd", x"db", x"d4", x"c9", x"bd", x"b1", x"a7", x"a0", 
        x"9c", x"9f", x"a5", x"a9", x"a6", x"a9", x"aa", x"ad", x"b0", x"a4", x"8d", x"6f", x"54", x"33", x"15", 
        x"07", x"06", x"0e", x"1b", x"2a", x"3a", x"48", x"54", x"5e", x"63", x"5e", x"52", x"4d", x"49", x"45", 
        x"41", x"3b", x"3c", x"45", x"58", x"76", x"98", x"b8", x"d3", x"e5", x"ea", x"e9", x"e3", x"e2", x"e1", 
        x"e3", x"e3", x"e4", x"e5", x"e7", x"df", x"d2", x"bc", x"99", x"73", x"4d", x"2b", x"10", x"08", x"0b", 
        x"88", x"88", x"86", x"86", x"85", x"84", x"84", x"84", x"85", x"85", x"84", x"83", x"83", x"85", x"85", 
        x"84", x"85", x"85", x"86", x"87", x"87", x"86", x"85", x"85", x"85", x"83", x"83", x"84", x"85", x"82", 
        x"84", x"86", x"86", x"85", x"82", x"82", x"85", x"84", x"83", x"85", x"87", x"86", x"83", x"87", x"88", 
        x"87", x"85", x"85", x"85", x"86", x"87", x"85", x"86", x"83", x"83", x"85", x"85", x"88", x"85", x"83", 
        x"85", x"86", x"86", x"85", x"86", x"84", x"84", x"86", x"88", x"88", x"87", x"86", x"85", x"88", x"89", 
        x"86", x"83", x"87", x"8b", x"8a", x"86", x"88", x"88", x"86", x"88", x"88", x"88", x"85", x"89", x"8a", 
        x"89", x"87", x"85", x"87", x"8a", x"87", x"89", x"89", x"88", x"8b", x"89", x"8c", x"8d", x"8f", x"90", 
        x"8f", x"8a", x"5e", x"25", x"3d", x"35", x"24", x"12", x"09", x"15", x"30", x"3f", x"48", x"48", x"43", 
        x"3e", x"3b", x"36", x"39", x"4e", x"5a", x"3a", x"7b", x"7d", x"3f", x"35", x"3b", x"40", x"3e", x"3c", 
        x"3e", x"43", x"43", x"41", x"40", x"3d", x"3f", x"40", x"3d", x"3d", x"3b", x"3a", x"39", x"3c", x"3e", 
        x"3a", x"9c", x"df", x"d5", x"d3", x"d5", x"d8", x"da", x"d0", x"cf", x"d1", x"d0", x"cf", x"cf", x"cf", 
        x"d0", x"cf", x"cf", x"d1", x"d3", x"d2", x"d1", x"d1", x"d2", x"d1", x"d0", x"d2", x"d1", x"d1", x"d2", 
        x"d4", x"d5", x"d4", x"d2", x"d1", x"d1", x"d2", x"d4", x"d2", x"d1", x"d0", x"d1", x"d2", x"d3", x"d3", 
        x"d3", x"d1", x"d5", x"dc", x"ce", x"a9", x"8e", x"99", x"be", x"d6", x"d5", x"cf", x"d1", x"d3", x"d2", 
        x"d5", x"ec", x"f0", x"ea", x"ea", x"ef", x"ed", x"ee", x"ed", x"ec", x"ed", x"f1", x"f3", x"f1", x"e9", 
        x"de", x"d2", x"c5", x"b6", x"ac", x"ab", x"b8", x"cd", x"e2", x"f1", x"f5", x"f3", x"f0", x"ef", x"ee", 
        x"ee", x"ee", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ee", x"ee", x"ef", 
        x"f1", x"f0", x"ef", x"ee", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"eb", x"ec", x"f1", x"ef", x"ee", 
        x"ef", x"f0", x"ee", x"ed", x"f1", x"f1", x"f0", x"f2", x"f1", x"f1", x"ef", x"ef", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f0", x"ee", x"ee", x"f0", x"f0", 
        x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"ef", x"e3", 
        x"d2", x"c7", x"be", x"bb", x"c4", x"d6", x"ec", x"f3", x"f6", x"f3", x"f0", x"f0", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", 
        x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"ef", x"ee", x"f3", x"f2", x"f3", x"f4", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f4", x"f4", x"f3", x"f2", 
        x"f3", x"f4", x"f3", x"f3", x"f0", x"f0", x"f2", x"f4", x"f2", x"f5", x"f3", x"f2", x"f2", x"f3", x"f2", 
        x"f1", x"e4", x"d8", x"c9", x"ba", x"ba", x"cc", x"e5", x"f4", x"f7", x"f3", x"f0", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"ea", x"ed", x"f2", x"f0", x"ee", x"ef", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"f1", x"f0", 
        x"ee", x"f0", x"ef", x"ee", x"f0", x"f1", x"f2", x"ee", x"ef", x"f2", x"f1", x"ed", x"e4", x"db", x"d5", 
        x"d8", x"d8", x"bb", x"98", x"7e", x"78", x"85", x"8e", x"8e", x"8d", x"8b", x"8d", x"8f", x"8f", x"8d", 
        x"8e", x"8f", x"8c", x"8d", x"8e", x"8d", x"8d", x"8e", x"8e", x"8d", x"8c", x"8b", x"8c", x"8d", x"8d", 
        x"8d", x"8c", x"8d", x"8e", x"8b", x"8b", x"88", x"8a", x"85", x"9c", x"df", x"dd", x"dd", x"dc", x"db", 
        x"da", x"d8", x"da", x"db", x"db", x"da", x"d9", x"d9", x"d8", x"d9", x"db", x"db", x"db", x"dd", x"db", 
        x"db", x"da", x"da", x"dd", x"e1", x"df", x"d2", x"c0", x"b3", x"a9", x"a2", x"9f", x"a1", x"a6", x"aa", 
        x"aa", x"aa", x"ac", x"b1", x"b6", x"b4", x"9b", x"78", x"58", x"3e", x"21", x"0c", x"04", x"04", x"0a", 
        x"1d", x"34", x"4b", x"59", x"5f", x"60", x"5e", x"59", x"4f", x"4b", x"4b", x"42", x"38", x"32", x"33", 
        x"48", x"66", x"8c", x"af", x"cd", x"dd", x"e7", x"eb", x"e8", x"e3", x"e1", x"e3", x"e2", x"e2", x"e6", 
        x"ec", x"ed", x"e5", x"cd", x"a6", x"7c", x"52", x"35", x"1a", x"07", x"03", x"0c", x"1d", x"2f", x"3e", 
        x"8a", x"89", x"88", x"88", x"87", x"86", x"84", x"84", x"84", x"85", x"85", x"85", x"84", x"84", x"85", 
        x"85", x"84", x"83", x"83", x"84", x"86", x"86", x"85", x"84", x"83", x"83", x"84", x"83", x"83", x"85", 
        x"83", x"84", x"86", x"86", x"84", x"82", x"82", x"84", x"86", x"85", x"84", x"83", x"85", x"86", x"87", 
        x"85", x"86", x"87", x"85", x"85", x"87", x"86", x"86", x"85", x"86", x"86", x"84", x"87", x"87", x"87", 
        x"86", x"86", x"87", x"85", x"86", x"86", x"86", x"87", x"88", x"87", x"86", x"85", x"88", x"89", x"89", 
        x"87", x"86", x"86", x"88", x"89", x"87", x"87", x"87", x"86", x"88", x"88", x"88", x"87", x"88", x"88", 
        x"87", x"87", x"87", x"87", x"88", x"87", x"87", x"88", x"89", x"89", x"89", x"89", x"86", x"87", x"89", 
        x"8b", x"93", x"6c", x"34", x"6b", x"73", x"6c", x"5e", x"4f", x"4b", x"4a", x"43", x"41", x"45", x"45", 
        x"44", x"44", x"41", x"44", x"49", x"43", x"34", x"7d", x"7d", x"40", x"3b", x"3c", x"41", x"3f", x"3c", 
        x"40", x"41", x"40", x"41", x"41", x"40", x"41", x"3f", x"3c", x"3b", x"38", x"38", x"38", x"36", x"36", 
        x"38", x"9d", x"e0", x"d4", x"d2", x"d3", x"d6", x"da", x"d1", x"d0", x"d1", x"cf", x"cf", x"d0", x"d0", 
        x"d0", x"d0", x"d0", x"cf", x"d1", x"d3", x"d2", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", 
        x"d4", x"d4", x"d1", x"d2", x"d1", x"d0", x"d2", x"d3", x"d2", x"d0", x"cf", x"d2", x"d4", x"d1", x"ce", 
        x"d1", x"d6", x"ce", x"ad", x"92", x"9d", x"b5", x"ca", x"dc", x"d4", x"ce", x"d0", x"d2", x"d2", x"d3", 
        x"d6", x"ec", x"ef", x"ed", x"ed", x"ee", x"ee", x"ee", x"ed", x"ed", x"ed", x"ee", x"ef", x"ed", x"eb", 
        x"ee", x"ef", x"ec", x"e3", x"db", x"cd", x"be", x"af", x"a7", x"b0", x"c5", x"d8", x"e8", x"ef", x"f1", 
        x"f0", x"f0", x"ed", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"f0", x"ee", 
        x"ed", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f0", x"ef", x"ef", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"ed", x"ec", x"f0", x"ef", x"ee", 
        x"ef", x"f1", x"ef", x"ef", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"ee", x"e5", x"d6", x"c9", x"c1", x"bb", x"bf", x"d3", x"e7", x"ef", x"f1", x"f1", x"f5", x"f2", 
        x"f0", x"ef", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f3", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"ee", x"ec", x"f2", x"f3", x"f3", x"f4", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f1", x"f2", x"f2", x"f0", x"ef", 
        x"f1", x"f4", x"f4", x"ef", x"e3", x"d3", x"c5", x"b9", x"c4", x"d6", x"e6", x"f0", x"f0", x"ee", x"f0", 
        x"f1", x"f0", x"f0", x"f2", x"f2", x"f0", x"ef", x"f1", x"f0", x"f0", x"f1", x"f3", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"eb", x"ef", x"f1", x"f1", x"f0", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"ef", x"f0", x"f2", x"f1", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ed", x"e5", 
        x"de", x"db", x"d9", x"d4", x"c4", x"a7", x"8b", x"7c", x"80", x"8a", x"8d", x"8c", x"8e", x"8e", x"8d", 
        x"8e", x"8e", x"8c", x"8d", x"8e", x"8c", x"8b", x"8d", x"90", x"8f", x"8d", x"8c", x"8c", x"8c", x"8c", 
        x"8c", x"8c", x"8d", x"8c", x"8b", x"8c", x"89", x"8b", x"85", x"96", x"df", x"de", x"dd", x"db", x"da", 
        x"d8", x"d7", x"d9", x"da", x"da", x"db", x"da", x"da", x"d9", x"da", x"d9", x"da", x"db", x"da", x"dc", 
        x"e0", x"df", x"d9", x"c8", x"b9", x"af", x"a5", x"a0", x"a0", x"a4", x"a5", x"a5", x"a7", x"aa", x"ae", 
        x"b5", x"b1", x"9c", x"89", x"7b", x"60", x"35", x"1e", x"0e", x"08", x"0a", x"17", x"2a", x"3e", x"4c", 
        x"57", x"5c", x"5c", x"57", x"52", x"4d", x"49", x"47", x"3f", x"33", x"31", x"42", x"5f", x"7f", x"9f", 
        x"bb", x"d1", x"e1", x"e7", x"e9", x"e4", x"e0", x"e6", x"e5", x"e1", x"e5", x"ea", x"e8", x"e0", x"d0", 
        x"b1", x"88", x"63", x"41", x"28", x"15", x"0a", x"0c", x"15", x"23", x"34", x"41", x"4b", x"4c", x"48", 
        x"8a", x"89", x"88", x"88", x"87", x"86", x"84", x"85", x"85", x"85", x"84", x"84", x"84", x"84", x"85", 
        x"86", x"86", x"85", x"81", x"81", x"84", x"86", x"85", x"84", x"84", x"84", x"84", x"83", x"84", x"86", 
        x"83", x"82", x"84", x"85", x"85", x"84", x"83", x"85", x"86", x"85", x"84", x"85", x"85", x"85", x"87", 
        x"85", x"86", x"88", x"85", x"85", x"85", x"84", x"85", x"86", x"88", x"86", x"84", x"86", x"86", x"87", 
        x"86", x"86", x"88", x"86", x"87", x"85", x"86", x"87", x"87", x"87", x"87", x"87", x"87", x"86", x"86", 
        x"87", x"88", x"88", x"88", x"88", x"88", x"88", x"87", x"87", x"87", x"88", x"87", x"88", x"88", x"86", 
        x"87", x"89", x"88", x"88", x"88", x"87", x"87", x"88", x"88", x"87", x"87", x"87", x"89", x"89", x"8b", 
        x"89", x"90", x"66", x"2f", x"68", x"77", x"7e", x"7f", x"7b", x"77", x"73", x"66", x"58", x"4d", x"43", 
        x"40", x"42", x"40", x"46", x"47", x"3a", x"32", x"7c", x"80", x"41", x"3c", x"3d", x"40", x"3f", x"3c", 
        x"41", x"42", x"41", x"40", x"40", x"44", x"46", x"43", x"42", x"43", x"40", x"40", x"3f", x"3b", x"35", 
        x"35", x"98", x"de", x"d3", x"d2", x"d4", x"d7", x"dc", x"d0", x"d1", x"d2", x"cf", x"cf", x"d0", x"cf", 
        x"cf", x"d1", x"d0", x"cf", x"d0", x"d3", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d0", 
        x"d0", x"d4", x"d1", x"d1", x"d0", x"cf", x"d2", x"d3", x"d2", x"cd", x"d4", x"d4", x"ce", x"d4", x"d2", 
        x"cf", x"b2", x"92", x"95", x"b9", x"cc", x"d3", x"cf", x"d7", x"d3", x"d0", x"d1", x"d2", x"d3", x"d3", 
        x"d4", x"ed", x"f0", x"ee", x"ef", x"ef", x"f0", x"ef", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ec", 
        x"ed", x"ed", x"ec", x"ef", x"f2", x"f1", x"eb", x"e2", x"d7", x"c9", x"ba", x"af", x"ab", x"bc", x"ce", 
        x"e0", x"ec", x"ef", x"f4", x"ef", x"ee", x"f0", x"f1", x"f1", x"ef", x"ed", x"ef", x"f0", x"ee", x"ec", 
        x"ef", x"f2", x"ef", x"ed", x"ef", x"ef", x"ef", x"f1", x"f2", x"f3", x"f2", x"f1", x"f0", x"ef", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"ec", x"eb", x"f0", x"f0", x"ef", 
        x"ef", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", 
        x"ef", x"ef", x"f2", x"f3", x"ee", x"e6", x"d8", x"c3", x"b7", x"b2", x"bd", x"d5", x"e9", x"f2", x"f2", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"ef", x"ef", x"f0", x"f1", x"f2", x"f2", x"ef", x"f0", x"f0", x"f0", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"ef", 
        x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"ee", x"eb", x"f2", x"f4", x"f3", x"f4", x"f4", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f3", x"f3", x"ec", x"df", x"cd", x"be", x"b9", x"c6", x"dd", x"ee", x"f1", 
        x"ef", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"f0", x"f3", x"f0", x"ef", x"f0", x"f0", x"f2", x"f3", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"f1", 
        x"ec", x"ef", x"f2", x"f0", x"f1", x"ee", x"ef", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"f1", 
        x"f1", x"e9", x"e1", x"df", x"d9", x"db", x"ce", x"ad", x"88", x"7d", x"83", x"8a", x"8f", x"90", x"8d", 
        x"8e", x"90", x"8c", x"8a", x"8b", x"8b", x"8c", x"8d", x"8d", x"8d", x"8e", x"8d", x"8c", x"8c", x"8b", 
        x"8c", x"8d", x"8d", x"8c", x"8c", x"8b", x"8a", x"8c", x"86", x"93", x"de", x"de", x"dd", x"dc", x"dc", 
        x"dc", x"db", x"d9", x"db", x"de", x"dc", x"da", x"d9", x"dc", x"dc", x"da", x"dc", x"e0", x"e0", x"dd", 
        x"ce", x"be", x"b1", x"a7", x"a0", x"a2", x"a4", x"a4", x"a7", x"a9", x"aa", x"ad", x"b6", x"b1", x"9d", 
        x"84", x"5a", x"38", x"27", x"24", x"17", x"0c", x"0c", x"16", x"2e", x"42", x"4e", x"58", x"5c", x"56", 
        x"52", x"4f", x"49", x"46", x"44", x"3f", x"35", x"32", x"48", x"67", x"8a", x"b1", x"c9", x"d9", x"e4", 
        x"e5", x"e5", x"e4", x"e2", x"e4", x"e4", x"e3", x"e5", x"ea", x"e8", x"e1", x"cd", x"a6", x"7a", x"4c", 
        x"30", x"1a", x"0e", x"08", x"0e", x"18", x"2c", x"39", x"45", x"4f", x"51", x"47", x"3c", x"32", x"2a", 
        x"8a", x"88", x"87", x"87", x"87", x"86", x"85", x"87", x"87", x"85", x"84", x"84", x"85", x"86", x"84", 
        x"84", x"86", x"86", x"83", x"83", x"84", x"85", x"85", x"86", x"85", x"85", x"85", x"85", x"85", x"85", 
        x"84", x"83", x"83", x"84", x"85", x"86", x"87", x"85", x"84", x"85", x"87", x"87", x"85", x"86", x"87", 
        x"85", x"86", x"89", x"85", x"85", x"85", x"85", x"86", x"87", x"88", x"87", x"86", x"86", x"85", x"87", 
        x"87", x"87", x"87", x"86", x"87", x"86", x"86", x"86", x"87", x"87", x"88", x"89", x"87", x"87", x"87", 
        x"87", x"87", x"87", x"87", x"88", x"88", x"88", x"89", x"89", x"88", x"88", x"87", x"88", x"88", x"86", 
        x"87", x"89", x"88", x"88", x"88", x"88", x"88", x"88", x"89", x"88", x"87", x"88", x"8a", x"88", x"88", 
        x"8b", x"92", x"68", x"2f", x"65", x"72", x"75", x"75", x"76", x"77", x"79", x"77", x"75", x"75", x"73", 
        x"6b", x"61", x"4c", x"45", x"43", x"3c", x"32", x"7b", x"7d", x"42", x"40", x"40", x"3f", x"40", x"40", 
        x"43", x"43", x"41", x"40", x"42", x"44", x"46", x"44", x"43", x"43", x"42", x"43", x"45", x"45", x"40", 
        x"39", x"94", x"db", x"d2", x"d3", x"d5", x"d8", x"dc", x"d0", x"d1", x"d2", x"d0", x"d0", x"d1", x"cf", 
        x"cf", x"d1", x"d1", x"cf", x"d0", x"d3", x"d2", x"d1", x"d1", x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", 
        x"d5", x"d3", x"d3", x"d4", x"d1", x"d1", x"d5", x"d3", x"d3", x"cf", x"d2", x"d6", x"d6", x"d1", x"b3", 
        x"8c", x"95", x"b7", x"cb", x"d3", x"d2", x"ce", x"cc", x"d7", x"d4", x"d1", x"d2", x"d1", x"d2", x"d2", 
        x"d4", x"ed", x"f0", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ec", 
        x"ee", x"ee", x"ec", x"eb", x"ee", x"f0", x"ef", x"ef", x"f2", x"f1", x"ea", x"e1", x"d3", x"c5", x"b3", 
        x"a7", x"b1", x"c3", x"d9", x"e8", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", x"ed", 
        x"ee", x"f0", x"ee", x"ed", x"ed", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"eb", x"eb", x"f1", x"f1", x"ef", 
        x"ef", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f2", x"f0", x"f0", x"ef", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f0", 
        x"f2", x"f1", x"ef", x"f1", x"f3", x"f1", x"eb", x"ec", x"e9", x"da", x"c2", x"b2", x"ae", x"c0", x"d4", 
        x"e7", x"f1", x"f2", x"f2", x"f2", x"f0", x"f2", x"f2", x"f1", x"f2", x"f4", x"f1", x"f1", x"ef", x"ed", 
        x"f1", x"f1", x"f0", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"ef", x"ec", x"f2", x"f3", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f5", x"f0", x"e9", x"dc", x"c4", x"b1", x"b6", x"d2", 
        x"e7", x"f1", x"f3", x"ef", x"ef", x"f1", x"f1", x"f0", x"f2", x"f2", x"f1", x"f2", x"f3", x"f4", x"f4", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"ee", x"f2", 
        x"ee", x"ef", x"f2", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"f1", x"ef", 
        x"f1", x"f3", x"f2", x"ed", x"e6", x"d9", x"d3", x"d6", x"d3", x"b3", x"8b", x"7c", x"7f", x"87", x"8e", 
        x"8f", x"8d", x"92", x"92", x"8f", x"8d", x"8e", x"8d", x"8c", x"90", x"91", x"8e", x"8e", x"8d", x"8d", 
        x"8d", x"8e", x"8e", x"8d", x"8d", x"8c", x"8c", x"8e", x"86", x"8f", x"dd", x"e1", x"de", x"db", x"da", 
        x"db", x"df", x"d9", x"d9", x"db", x"db", x"da", x"da", x"dc", x"df", x"de", x"d8", x"cb", x"bb", x"af", 
        x"a7", x"a5", x"a6", x"a4", x"a7", x"a9", x"ac", x"ac", x"af", x"b7", x"ad", x"9c", x"7d", x"50", x"2e", 
        x"22", x"1b", x"1d", x"26", x"3c", x"26", x"0f", x"12", x"4d", x"64", x"5a", x"4c", x"4a", x"4a", x"48", 
        x"45", x"41", x"39", x"2e", x"2e", x"4b", x"75", x"a2", x"c5", x"d7", x"e4", x"ea", x"e7", x"e4", x"e4", 
        x"e2", x"e3", x"e5", x"e3", x"e5", x"e7", x"e2", x"d6", x"bd", x"94", x"66", x"3b", x"21", x"13", x"09", 
        x"08", x"10", x"1c", x"2b", x"3b", x"47", x"4b", x"49", x"43", x"3b", x"32", x"2b", x"28", x"25", x"25", 
        x"8a", x"88", x"86", x"86", x"87", x"87", x"86", x"88", x"88", x"86", x"85", x"85", x"86", x"87", x"85", 
        x"83", x"82", x"84", x"86", x"87", x"86", x"83", x"84", x"85", x"85", x"85", x"84", x"85", x"86", x"86", 
        x"85", x"84", x"83", x"84", x"85", x"87", x"88", x"86", x"85", x"85", x"86", x"87", x"87", x"86", x"87", 
        x"85", x"86", x"89", x"86", x"86", x"86", x"87", x"89", x"88", x"87", x"86", x"86", x"86", x"85", x"87", 
        x"87", x"88", x"87", x"86", x"87", x"89", x"88", x"87", x"86", x"86", x"87", x"87", x"86", x"87", x"88", 
        x"87", x"86", x"87", x"88", x"87", x"87", x"88", x"89", x"89", x"88", x"88", x"88", x"89", x"88", x"86", 
        x"87", x"89", x"89", x"88", x"89", x"89", x"89", x"89", x"89", x"89", x"89", x"8a", x"8b", x"88", x"89", 
        x"8b", x"91", x"67", x"2f", x"66", x"75", x"77", x"76", x"75", x"74", x"79", x"77", x"75", x"73", x"75", 
        x"7a", x"7d", x"7c", x"70", x"6e", x"63", x"40", x"78", x"7c", x"3f", x"3c", x"3f", x"3c", x"3e", x"40", 
        x"41", x"40", x"3e", x"40", x"40", x"3f", x"41", x"44", x"46", x"44", x"45", x"43", x"43", x"44", x"42", 
        x"3b", x"96", x"dd", x"d4", x"d3", x"d5", x"d7", x"db", x"cf", x"d1", x"d3", x"d1", x"d1", x"d1", x"cf", 
        x"cf", x"d1", x"d1", x"d0", x"d1", x"d3", x"d2", x"d0", x"d0", x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", 
        x"d3", x"d4", x"d6", x"d4", x"cf", x"cd", x"d1", x"d1", x"d0", x"d3", x"d5", x"ce", x"b0", x"91", x"99", 
        x"be", x"d4", x"d1", x"d0", x"d0", x"cf", x"d1", x"cf", x"da", x"d5", x"d0", x"d0", x"d1", x"d2", x"d1", 
        x"d4", x"ed", x"f0", x"ee", x"ef", x"ed", x"ed", x"ee", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ec", 
        x"ef", x"f0", x"ed", x"eb", x"eb", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"f1", x"ef", x"f0", x"ed", 
        x"e4", x"d2", x"bf", x"ae", x"ac", x"b6", x"c8", x"dc", x"e7", x"ed", x"ee", x"f1", x"f2", x"f0", x"ef", 
        x"f0", x"f1", x"f1", x"ef", x"ed", x"f1", x"f0", x"ef", x"ef", x"f1", x"f2", x"f0", x"f1", x"f1", x"ef", 
        x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"eb", x"eb", x"f1", x"f1", x"ef", 
        x"ee", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f2", x"f0", x"f0", x"ee", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"f0", x"f3", x"f4", x"f4", x"f1", x"f3", x"f5", x"f2", x"ec", x"e0", x"c8", x"b7", 
        x"af", x"bb", x"d3", x"e4", x"ec", x"f2", x"f4", x"f3", x"f1", x"f2", x"f3", x"ef", x"f2", x"f1", x"f1", 
        x"f2", x"f0", x"ef", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"ef", x"ed", x"f2", x"f2", x"f0", x"f2", x"f3", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"f0", x"f2", x"f2", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"ea", x"d6", x"bb", 
        x"b2", x"bf", x"d9", x"e7", x"ef", x"ef", x"ee", x"ee", x"f0", x"f4", x"f4", x"f1", x"f1", x"f2", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f2", 
        x"ef", x"ef", x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", 
        x"f1", x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ed", x"ee", x"f3", x"f1", 
        x"ef", x"ef", x"f2", x"f2", x"ed", x"f0", x"e9", x"da", x"d0", x"d4", x"da", x"be", x"9b", x"84", x"82", 
        x"88", x"8a", x"8e", x"8e", x"8d", x"8c", x"8f", x"8f", x"8d", x"8b", x"8c", x"8e", x"8e", x"8e", x"8e", 
        x"8e", x"8e", x"8e", x"8c", x"8d", x"8e", x"8f", x"8f", x"86", x"88", x"d9", x"e0", x"dd", x"de", x"dd", 
        x"db", x"db", x"dd", x"dc", x"dd", x"df", x"de", x"da", x"d2", x"c0", x"ae", x"a8", x"a9", x"a7", x"a7", 
        x"ac", x"ad", x"ab", x"ac", x"b1", x"b1", x"ad", x"a0", x"8a", x"64", x"39", x"20", x"1e", x"20", x"2f", 
        x"4d", x"64", x"6c", x"59", x"6d", x"41", x"0b", x"17", x"5c", x"6a", x"54", x"46", x"3f", x"34", x"35", 
        x"33", x"3c", x"5b", x"88", x"b2", x"d1", x"e1", x"e6", x"e5", x"e6", x"e5", x"e3", x"e2", x"e3", x"e6", 
        x"e5", x"e5", x"e7", x"e2", x"d3", x"b1", x"7e", x"49", x"27", x"13", x"0b", x"07", x"0a", x"12", x"21", 
        x"2c", x"38", x"41", x"46", x"46", x"45", x"43", x"3e", x"38", x"32", x"2e", x"2d", x"2c", x"2b", x"29", 
        x"8a", x"88", x"86", x"86", x"87", x"87", x"87", x"87", x"87", x"87", x"87", x"86", x"86", x"86", x"86", 
        x"86", x"84", x"85", x"85", x"86", x"85", x"84", x"83", x"85", x"85", x"84", x"84", x"85", x"86", x"85", 
        x"86", x"86", x"84", x"84", x"85", x"87", x"87", x"87", x"87", x"85", x"85", x"86", x"88", x"86", x"88", 
        x"85", x"87", x"89", x"86", x"86", x"87", x"88", x"88", x"88", x"87", x"87", x"87", x"85", x"85", x"86", 
        x"87", x"88", x"88", x"88", x"88", x"89", x"88", x"87", x"87", x"87", x"87", x"87", x"85", x"86", x"87", 
        x"87", x"87", x"89", x"89", x"86", x"87", x"88", x"89", x"89", x"88", x"88", x"88", x"89", x"89", x"87", 
        x"87", x"89", x"89", x"89", x"8a", x"8a", x"8a", x"89", x"89", x"89", x"8a", x"89", x"8a", x"8a", x"8b", 
        x"8b", x"90", x"67", x"31", x"63", x"72", x"75", x"78", x"7a", x"76", x"78", x"76", x"76", x"77", x"76", 
        x"75", x"76", x"78", x"70", x"7a", x"78", x"47", x"73", x"7f", x"43", x"3d", x"45", x"40", x"3d", x"3f", 
        x"3e", x"3e", x"3c", x"41", x"43", x"42", x"40", x"3c", x"3d", x"43", x"46", x"46", x"42", x"41", x"3f", 
        x"3b", x"98", x"de", x"d4", x"d4", x"d5", x"d7", x"dc", x"d0", x"d1", x"d3", x"d1", x"d1", x"d2", x"d0", 
        x"cf", x"d1", x"d2", x"d1", x"d2", x"d3", x"d2", x"d0", x"d0", x"d3", x"d3", x"d3", x"d2", x"d2", x"d3", 
        x"d5", x"d5", x"d4", x"d3", x"d2", x"d1", x"d0", x"d4", x"d4", x"cb", x"b7", x"9a", x"99", x"bb", x"d0", 
        x"d5", x"cd", x"cd", x"d1", x"ce", x"d1", x"d1", x"ce", x"d9", x"d4", x"d0", x"d1", x"d2", x"d2", x"d1", 
        x"d3", x"ec", x"f0", x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ed", x"ef", x"f0", x"ed", 
        x"ef", x"f0", x"ee", x"ed", x"ee", x"f0", x"ee", x"ee", x"ee", x"f0", x"ef", x"ef", x"ec", x"ec", x"ef", 
        x"f1", x"ee", x"ec", x"e8", x"dc", x"cc", x"b9", x"af", x"b5", x"c3", x"d3", x"de", x"e5", x"ea", x"ef", 
        x"f1", x"ef", x"ed", x"ed", x"ef", x"ee", x"ed", x"ee", x"ee", x"ed", x"ed", x"f0", x"f1", x"f1", x"ef", 
        x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"eb", x"eb", x"f1", x"f1", x"ef", 
        x"ee", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f2", x"f0", x"f0", x"ee", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ef", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"f3", x"f3", x"f0", x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"eb", 
        x"dc", x"c4", x"b6", x"b8", x"c3", x"d4", x"e2", x"ee", x"f3", x"f3", x"f4", x"f3", x"f2", x"f0", x"f0", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"ed", x"f2", x"f1", x"f0", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f2", x"f2", x"f4", x"f5", x"f4", x"f1", x"ed", 
        x"e2", x"cc", x"b6", x"b4", x"c7", x"dd", x"e9", x"ee", x"f1", x"f2", x"f0", x"f0", x"f3", x"f3", x"f0", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", 
        x"ef", x"ed", x"f2", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", 
        x"f1", x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f3", x"ef", x"ef", x"f0", x"e9", x"da", x"d0", x"d5", x"d5", x"c2", x"9f", 
        x"86", x"83", x"85", x"8a", x"8f", x"8f", x"8d", x"8f", x"90", x"91", x"8f", x"8e", x"8f", x"8f", x"8f", 
        x"8f", x"8e", x"8e", x"8d", x"8c", x"8d", x"8d", x"8e", x"87", x"86", x"d1", x"e1", x"dc", x"da", x"da", 
        x"da", x"dd", x"de", x"d9", x"d3", x"ca", x"bf", x"b1", x"a3", x"a5", x"a5", x"a9", x"b0", x"b0", x"b1", 
        x"b5", x"b5", x"b0", x"a7", x"98", x"7d", x"5a", x"33", x"1e", x"24", x"2b", x"3c", x"56", x"65", x"6e", 
        x"75", x"70", x"68", x"4d", x"6e", x"48", x"10", x"17", x"5a", x"65", x"4b", x"41", x"43", x"4e", x"6a", 
        x"92", x"b7", x"d4", x"e2", x"e6", x"e7", x"e5", x"e5", x"e3", x"e2", x"e4", x"e6", x"ea", x"eb", x"e7", 
        x"db", x"c5", x"a8", x"7e", x"58", x"33", x"10", x"0a", x"06", x"03", x"08", x"15", x"27", x"34", x"3d", 
        x"3f", x"42", x"43", x"46", x"46", x"45", x"41", x"3d", x"39", x"37", x"36", x"33", x"2d", x"2a", x"27", 
        x"89", x"88", x"87", x"87", x"88", x"87", x"86", x"86", x"87", x"88", x"88", x"87", x"86", x"85", x"84", 
        x"85", x"88", x"87", x"84", x"84", x"87", x"87", x"84", x"85", x"85", x"85", x"86", x"86", x"86", x"85", 
        x"86", x"86", x"86", x"85", x"85", x"86", x"86", x"87", x"87", x"86", x"85", x"86", x"87", x"87", x"88", 
        x"86", x"87", x"89", x"86", x"86", x"86", x"86", x"86", x"87", x"88", x"88", x"89", x"88", x"88", x"87", 
        x"88", x"88", x"87", x"88", x"87", x"87", x"88", x"88", x"88", x"89", x"89", x"89", x"88", x"88", x"88", 
        x"88", x"88", x"88", x"88", x"86", x"87", x"87", x"88", x"89", x"89", x"89", x"89", x"8a", x"89", x"87", 
        x"88", x"8a", x"8a", x"89", x"8a", x"8b", x"8a", x"89", x"89", x"8a", x"8b", x"8a", x"89", x"86", x"89", 
        x"8b", x"91", x"67", x"2d", x"5f", x"72", x"76", x"77", x"7a", x"77", x"79", x"77", x"76", x"77", x"76", 
        x"73", x"71", x"77", x"6e", x"77", x"7b", x"46", x"6c", x"7b", x"3e", x"3d", x"5f", x"69", x"5f", x"54", 
        x"45", x"3e", x"3c", x"3e", x"3c", x"3d", x"3d", x"34", x"31", x"38", x"3c", x"40", x"42", x"42", x"42", 
        x"3e", x"97", x"dd", x"d4", x"d4", x"d6", x"d8", x"dd", x"d1", x"d1", x"d3", x"d1", x"d1", x"d2", x"d0", 
        x"cf", x"d1", x"d2", x"d1", x"d2", x"d3", x"d2", x"d1", x"d1", x"d3", x"d3", x"d2", x"d2", x"d2", x"d4", 
        x"d2", x"d2", x"d3", x"cf", x"cd", x"d0", x"d3", x"d0", x"bc", x"98", x"97", x"b5", x"d1", x"d5", x"cf", 
        x"cf", x"ce", x"ce", x"cf", x"cf", x"ce", x"cf", x"cd", x"d7", x"d4", x"d0", x"d1", x"d1", x"d0", x"d0", 
        x"d3", x"eb", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", 
        x"ef", x"f0", x"ed", x"ee", x"ef", x"ed", x"ee", x"f0", x"f1", x"f1", x"ef", x"ed", x"ee", x"ed", x"ee", 
        x"ed", x"ed", x"ef", x"ef", x"ee", x"f0", x"ef", x"e6", x"d4", x"c0", x"af", x"b1", x"ba", x"c9", x"d9", 
        x"e3", x"e9", x"f0", x"f2", x"ef", x"ec", x"ec", x"ef", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"eb", x"eb", x"f1", x"f0", x"ef", 
        x"ef", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f2", x"f0", x"f0", x"ef", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f2", x"f4", x"f3", x"ef", x"f0", x"f1", x"f2", x"f4", x"f2", x"f2", x"f0", x"f0", x"f2", x"f3", x"f2", 
        x"f3", x"f3", x"ea", x"da", x"c6", x"b6", x"ba", x"c6", x"d5", x"e1", x"eb", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f1", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ee", x"f2", x"f1", x"f1", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f0", x"f0", x"f1", x"f2", x"f3", x"f4", x"f4", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"ea", x"d6", x"bf", x"b2", x"be", x"d3", x"e4", x"ee", x"f3", x"f2", x"ef", x"ef", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"ee", x"ed", x"f2", x"f1", x"f0", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f1", x"ef", x"ef", x"f0", x"f3", x"f1", x"ee", x"ed", x"db", x"cc", x"cd", x"d4", 
        x"c6", x"a3", x"89", x"81", x"85", x"8d", x"8e", x"8e", x"8f", x"8e", x"8e", x"8e", x"8f", x"8f", x"8f", 
        x"8f", x"8e", x"8e", x"8e", x"8c", x"8c", x"8b", x"8d", x"8a", x"86", x"c9", x"df", x"da", x"dc", x"de", 
        x"db", x"d5", x"c8", x"ba", x"ab", x"a2", x"a3", x"a6", x"a9", x"ab", x"ac", x"b3", x"b6", x"b4", x"b1", 
        x"a4", x"8f", x"76", x"50", x"2a", x"1a", x"23", x"30", x"3e", x"5c", x"70", x"78", x"73", x"6a", x"62", 
        x"61", x"60", x"5c", x"4b", x"69", x"42", x"0f", x"15", x"4f", x"63", x"62", x"7c", x"a0", x"c7", x"df", 
        x"eb", x"eb", x"e6", x"e3", x"e4", x"e6", x"e5", x"e5", x"e6", x"e9", x"ec", x"e3", x"d2", x"bd", x"9d", 
        x"70", x"48", x"26", x"0f", x"0c", x"0f", x"08", x"0a", x"09", x"03", x"0c", x"1a", x"27", x"31", x"3d", 
        x"3e", x"3f", x"40", x"45", x"46", x"44", x"45", x"41", x"3a", x"37", x"37", x"35", x"32", x"2e", x"2a", 
        x"88", x"87", x"87", x"88", x"89", x"88", x"86", x"86", x"86", x"87", x"87", x"87", x"86", x"84", x"84", 
        x"86", x"89", x"89", x"87", x"85", x"86", x"87", x"88", x"87", x"86", x"87", x"87", x"87", x"86", x"84", 
        x"85", x"87", x"87", x"86", x"85", x"85", x"86", x"85", x"85", x"87", x"88", x"87", x"85", x"86", x"88", 
        x"86", x"87", x"8a", x"86", x"86", x"87", x"86", x"86", x"86", x"87", x"88", x"88", x"88", x"8b", x"88", 
        x"88", x"88", x"86", x"88", x"87", x"88", x"89", x"89", x"89", x"89", x"89", x"89", x"8a", x"89", x"89", 
        x"89", x"89", x"88", x"87", x"87", x"87", x"87", x"87", x"88", x"8a", x"8a", x"89", x"8a", x"89", x"87", 
        x"88", x"8a", x"8a", x"89", x"8a", x"8b", x"8b", x"89", x"89", x"8a", x"89", x"8a", x"8c", x"88", x"89", 
        x"8c", x"8e", x"6c", x"41", x"60", x"6f", x"78", x"7a", x"7b", x"79", x"7a", x"7d", x"7b", x"75", x"75", 
        x"77", x"77", x"7a", x"72", x"79", x"79", x"42", x"67", x"7b", x"3e", x"3c", x"6d", x"84", x"7e", x"7f", 
        x"7b", x"70", x"64", x"5b", x"4b", x"42", x"40", x"36", x"31", x"33", x"32", x"39", x"43", x"48", x"48", 
        x"44", x"95", x"dc", x"d4", x"d5", x"d6", x"d7", x"dc", x"d1", x"d2", x"d3", x"d0", x"d0", x"d2", x"d1", 
        x"cf", x"d1", x"d2", x"d2", x"d3", x"d4", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d3", x"d4", 
        x"d4", x"d3", x"d1", x"d4", x"da", x"ce", x"af", x"96", x"96", x"b7", x"d7", x"dc", x"d4", x"d2", x"cf", 
        x"cf", x"d0", x"cf", x"ce", x"d1", x"d1", x"d2", x"ce", x"d7", x"d4", x"d2", x"d2", x"d1", x"d0", x"d0", 
        x"d2", x"eb", x"ef", x"ee", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", 
        x"ef", x"ef", x"ec", x"ec", x"ee", x"ef", x"ee", x"ed", x"ed", x"ed", x"ed", x"ed", x"ef", x"ee", x"f2", 
        x"f2", x"ef", x"f0", x"ef", x"ef", x"ed", x"ec", x"f0", x"f3", x"f1", x"ea", x"df", x"d0", x"bb", x"b2", 
        x"b4", x"be", x"cb", x"d8", x"e3", x"ee", x"f3", x"f3", x"f0", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"ec", x"eb", x"f0", x"f0", x"ef", 
        x"f0", x"f2", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"f0", x"f0", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", 
        x"ee", x"f0", x"f0", x"ee", x"f1", x"f3", x"f1", x"f1", x"f0", x"f4", x"f3", x"f1", x"f2", x"f1", x"f2", 
        x"f2", x"f1", x"f2", x"f4", x"f6", x"f2", x"e0", x"c9", x"bb", x"b9", x"bf", x"cb", x"da", x"ea", x"f6", 
        x"f5", x"f1", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"ef", x"f1", x"f0", x"ee", x"f2", x"f0", x"f2", x"f4", x"f4", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f4", x"f4", x"f3", x"f1", x"f0", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f4", x"f3", x"f4", x"f3", x"e6", x"ce", x"bc", x"b8", x"c1", x"d1", x"e6", x"f2", x"f4", x"f3", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", 
        x"ed", x"ec", x"f2", x"f1", x"f0", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f3", x"f2", 
        x"f0", x"f0", x"f1", x"f0", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"f0", x"f0", x"ef", x"e0", x"ca", 
        x"cb", x"d6", x"d1", x"b4", x"99", x"82", x"7c", x"86", x"8f", x"90", x"8d", x"8e", x"8e", x"8f", x"8f", 
        x"8f", x"8e", x"8c", x"8d", x"8e", x"90", x"8e", x"90", x"8d", x"87", x"c5", x"e0", x"d5", x"cb", x"c0", 
        x"b4", x"a6", x"a0", x"a2", x"a6", x"a9", x"ab", x"af", x"b4", x"ba", x"b9", x"b1", x"a0", x"81", x"5e", 
        x"38", x"17", x"12", x"27", x"39", x"53", x"6e", x"79", x"7d", x"7a", x"6f", x"63", x"60", x"60", x"5d", 
        x"57", x"4e", x"47", x"39", x"53", x"4a", x"43", x"65", x"95", x"bb", x"d7", x"ea", x"ec", x"ea", x"e3", 
        x"e2", x"e2", x"e3", x"e5", x"e7", x"e7", x"ea", x"ea", x"db", x"c7", x"ab", x"7d", x"53", x"30", x"15", 
        x"08", x"09", x"11", x"1d", x"31", x"37", x"21", x"1d", x"19", x"08", x"0c", x"1b", x"1f", x"27", x"35", 
        x"38", x"38", x"3b", x"43", x"45", x"41", x"40", x"3f", x"3d", x"3a", x"37", x"34", x"31", x"2e", x"2c", 
        x"89", x"89", x"88", x"88", x"88", x"87", x"86", x"87", x"87", x"87", x"86", x"86", x"85", x"85", x"86", 
        x"88", x"89", x"88", x"87", x"86", x"86", x"87", x"88", x"87", x"87", x"88", x"88", x"87", x"85", x"84", 
        x"85", x"87", x"87", x"87", x"86", x"85", x"87", x"85", x"85", x"86", x"88", x"88", x"87", x"88", x"89", 
        x"88", x"88", x"88", x"85", x"85", x"88", x"88", x"86", x"86", x"89", x"89", x"86", x"87", x"89", x"87", 
        x"88", x"88", x"89", x"89", x"88", x"88", x"89", x"89", x"89", x"89", x"88", x"87", x"89", x"89", x"89", 
        x"89", x"89", x"89", x"88", x"89", x"89", x"89", x"89", x"89", x"8a", x"8a", x"88", x"89", x"89", x"88", 
        x"89", x"89", x"89", x"89", x"89", x"89", x"89", x"8a", x"8a", x"89", x"88", x"89", x"8d", x"8b", x"8a", 
        x"8d", x"8a", x"79", x"83", x"71", x"70", x"77", x"7a", x"7b", x"77", x"79", x"7a", x"77", x"78", x"79", 
        x"7a", x"77", x"79", x"70", x"76", x"7a", x"46", x"6b", x"7d", x"3f", x"39", x"67", x"7d", x"76", x"7a", 
        x"7a", x"7c", x"7c", x"7b", x"74", x"6e", x"6c", x"4f", x"32", x"34", x"32", x"37", x"41", x"4e", x"54", 
        x"4d", x"92", x"de", x"d5", x"d5", x"d5", x"d5", x"db", x"d2", x"d1", x"d3", x"d1", x"d1", x"d1", x"d1", 
        x"d1", x"d0", x"d1", x"d1", x"d2", x"d4", x"d3", x"d2", x"d2", x"d3", x"d4", x"d4", x"d3", x"d3", x"d3", 
        x"d3", x"d7", x"d8", x"cb", x"ae", x"97", x"9c", x"b2", x"cd", x"d5", x"d1", x"d0", x"d0", x"d1", x"cf", 
        x"cf", x"d0", x"d1", x"cf", x"cf", x"d2", x"d1", x"ce", x"d9", x"d4", x"d1", x"d2", x"d2", x"d0", x"d0", 
        x"d0", x"ea", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ee", x"ed", x"ec", x"ee", x"ee", x"ed", x"ed", x"ee", x"ef", x"ed", x"eb", x"ed", x"ed", x"ef", 
        x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"ef", x"eb", x"e3", 
        x"d8", x"cc", x"c5", x"c0", x"bb", x"be", x"cc", x"dd", x"e9", x"ee", x"f1", x"f2", x"f0", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"f1", x"f2", x"f1", x"ef", x"ee", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f2", x"f1", x"f0", x"f1", x"ed", x"ed", x"ef", x"ef", x"f1", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", x"f0", x"f2", x"f2", x"f1", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f2", x"f2", x"f0", x"f3", x"f2", x"e9", x"dd", x"cf", x"c2", x"c0", x"c1", x"ca", 
        x"dc", x"ed", x"f4", x"f5", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f1", x"f0", x"f1", x"f0", x"f1", x"f2", x"f0", x"ee", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f4", x"f3", x"f1", x"f1", x"f2", x"f3", x"f1", 
        x"f1", x"f3", x"f2", x"f1", x"f2", x"f4", x"f2", x"eb", x"db", x"cd", x"c1", x"bd", x"c8", x"da", x"ea", 
        x"f2", x"f4", x"f1", x"ee", x"f1", x"f3", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", 
        x"ee", x"ed", x"f1", x"f0", x"ee", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f1", x"f0", x"ed", x"ef", x"ee", x"ef", x"f0", x"ed", x"ed", x"f0", x"f1", x"f0", x"f0", x"ea", 
        x"dd", x"d5", x"d5", x"d4", x"cb", x"ba", x"9e", x"87", x"81", x"89", x"90", x"8f", x"8e", x"8e", x"8f", 
        x"8e", x"8e", x"8e", x"8e", x"91", x"91", x"8f", x"8f", x"8d", x"87", x"aa", x"ba", x"b1", x"a6", x"a1", 
        x"a4", x"ab", x"af", x"b0", x"b4", x"b7", x"b8", x"b2", x"a7", x"90", x"70", x"54", x"39", x"22", x"22", 
        x"38", x"48", x"57", x"6a", x"74", x"79", x"76", x"6d", x"65", x"63", x"60", x"5b", x"59", x"52", x"4a", 
        x"42", x"3f", x"4c", x"5e", x"8a", x"a7", x"bf", x"d8", x"e7", x"e8", x"e8", x"e8", x"e3", x"e5", x"e5", 
        x"e5", x"e7", x"eb", x"e9", x"e2", x"cf", x"b4", x"96", x"6d", x"4a", x"2d", x"14", x"0d", x"13", x"1e", 
        x"2b", x"36", x"42", x"47", x"4b", x"41", x"24", x"22", x"1d", x"09", x"10", x"23", x"22", x"2e", x"3a", 
        x"37", x"35", x"37", x"3e", x"40", x"40", x"3e", x"3e", x"3c", x"39", x"36", x"35", x"35", x"34", x"30", 
        x"89", x"89", x"89", x"88", x"87", x"87", x"87", x"88", x"87", x"87", x"87", x"87", x"87", x"85", x"86", 
        x"87", x"88", x"87", x"86", x"86", x"87", x"88", x"87", x"86", x"86", x"87", x"87", x"86", x"85", x"84", 
        x"85", x"87", x"87", x"87", x"86", x"86", x"86", x"86", x"86", x"87", x"87", x"88", x"89", x"88", x"88", 
        x"88", x"87", x"87", x"86", x"86", x"88", x"87", x"87", x"87", x"89", x"89", x"85", x"87", x"88", x"87", 
        x"87", x"88", x"89", x"89", x"88", x"88", x"8a", x"88", x"87", x"89", x"89", x"87", x"89", x"8a", x"8a", 
        x"89", x"8a", x"8a", x"8a", x"8a", x"89", x"88", x"88", x"88", x"89", x"8a", x"88", x"87", x"88", x"89", 
        x"8a", x"8a", x"8a", x"8a", x"89", x"88", x"89", x"8c", x"8b", x"89", x"89", x"8a", x"8c", x"8b", x"87", 
        x"8d", x"89", x"7f", x"a5", x"7a", x"75", x"78", x"79", x"7c", x"7a", x"7a", x"79", x"77", x"7b", x"79", 
        x"7a", x"79", x"7b", x"71", x"79", x"7e", x"47", x"6a", x"79", x"3f", x"3a", x"67", x"7d", x"76", x"78", 
        x"74", x"76", x"76", x"79", x"7d", x"80", x"86", x"63", x"36", x"38", x"36", x"45", x"57", x"5b", x"55", 
        x"40", x"8d", x"dd", x"d5", x"d4", x"d4", x"d6", x"dc", x"d3", x"d2", x"d4", x"d3", x"d2", x"d2", x"d3", 
        x"d4", x"d0", x"d3", x"d2", x"d2", x"d3", x"d1", x"d3", x"d2", x"d2", x"d3", x"d1", x"d2", x"d4", x"d5", 
        x"d8", x"d2", x"b1", x"95", x"9a", x"b1", x"d0", x"d9", x"d3", x"cd", x"cd", x"d0", x"d2", x"d2", x"d2", 
        x"d1", x"d2", x"d1", x"cf", x"cf", x"d1", x"cf", x"ce", x"d9", x"d4", x"ce", x"d1", x"d1", x"d1", x"d1", 
        x"cf", x"e9", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ee", x"ed", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ec", x"ef", 
        x"f3", x"f2", x"ec", x"e1", x"d2", x"c5", x"bc", x"b7", x"ba", x"c6", x"d7", x"e9", x"f0", x"f2", x"f0", 
        x"ed", x"ee", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", 
        x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"f2", x"f1", x"f0", x"ef", x"eb", x"ed", x"ee", x"f0", x"f3", 
        x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f3", x"f2", x"f0", x"f5", x"f7", x"ec", x"dd", x"cc", x"bc", 
        x"b9", x"be", x"ca", x"df", x"ef", x"f5", x"f5", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"ef", x"f0", x"f3", x"f2", x"f2", x"f0", x"f1", x"ee", x"f1", x"f4", x"f3", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"e9", x"d4", x"c3", x"bc", x"c0", 
        x"d1", x"e5", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"ef", x"ee", x"ef", x"f0", x"ef", x"f1", x"f3", 
        x"ef", x"ed", x"ef", x"ef", x"ed", x"ee", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"f1", x"f1", x"ef", x"ef", x"f1", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ed", x"ee", 
        x"f2", x"ef", x"e5", x"d5", x"d1", x"d5", x"d3", x"c3", x"a6", x"8a", x"7e", x"83", x"8e", x"90", x"8e", 
        x"8f", x"92", x"91", x"90", x"8f", x"90", x"8f", x"8f", x"8f", x"8a", x"89", x"91", x"9d", x"aa", x"b0", 
        x"b0", x"af", x"b1", x"b4", x"b9", x"a7", x"91", x"65", x"44", x"2b", x"15", x"1f", x"38", x"4d", x"65", 
        x"75", x"79", x"77", x"73", x"6a", x"64", x"61", x"5e", x"5a", x"59", x"50", x"43", x"38", x"3c", x"52", 
        x"6a", x"89", x"aa", x"cc", x"e2", x"ea", x"eb", x"e9", x"e9", x"e5", x"e6", x"e5", x"e4", x"ea", x"ed", 
        x"ee", x"e1", x"ca", x"af", x"8a", x"5b", x"3a", x"21", x"0c", x"07", x"0e", x"1f", x"31", x"40", x"4b", 
        x"4f", x"49", x"43", x"36", x"2f", x"36", x"2e", x"20", x"1d", x"0e", x"1a", x"2a", x"21", x"32", x"3d", 
        x"36", x"32", x"33", x"38", x"3a", x"3d", x"3c", x"3b", x"3b", x"3a", x"38", x"36", x"35", x"36", x"33", 
        x"88", x"88", x"89", x"89", x"88", x"88", x"89", x"86", x"86", x"87", x"88", x"88", x"87", x"86", x"86", 
        x"86", x"88", x"87", x"86", x"86", x"87", x"89", x"89", x"86", x"86", x"87", x"87", x"87", x"86", x"84", 
        x"86", x"88", x"87", x"86", x"86", x"87", x"86", x"86", x"88", x"88", x"88", x"87", x"86", x"86", x"87", 
        x"87", x"87", x"88", x"8a", x"8b", x"88", x"86", x"87", x"87", x"88", x"88", x"85", x"88", x"89", x"87", 
        x"87", x"88", x"8a", x"8a", x"89", x"89", x"8b", x"89", x"86", x"86", x"89", x"8a", x"88", x"88", x"89", 
        x"89", x"8a", x"8a", x"8b", x"8b", x"89", x"88", x"87", x"87", x"8a", x"8c", x"88", x"87", x"88", x"89", 
        x"8a", x"8b", x"8c", x"8c", x"8b", x"8a", x"8a", x"8c", x"8d", x"8a", x"8a", x"8b", x"8c", x"8a", x"88", 
        x"8d", x"89", x"7d", x"a0", x"7c", x"78", x"7a", x"79", x"7c", x"7c", x"78", x"78", x"77", x"7a", x"79", 
        x"79", x"77", x"7c", x"73", x"79", x"7b", x"44", x"65", x"77", x"3f", x"3a", x"68", x"7d", x"77", x"7a", 
        x"78", x"78", x"77", x"77", x"77", x"79", x"81", x"5f", x"34", x"36", x"3a", x"69", x"7e", x"4a", x"2c", 
        x"24", x"8b", x"dc", x"d5", x"d3", x"d4", x"d5", x"da", x"d3", x"d3", x"d5", x"d4", x"d3", x"d3", x"d3", 
        x"d1", x"d1", x"d4", x"d1", x"d1", x"d1", x"d2", x"d1", x"d3", x"d4", x"d2", x"d1", x"d1", x"d6", x"d5", 
        x"ab", x"8e", x"9c", x"ba", x"d1", x"d8", x"d3", x"d3", x"d0", x"ce", x"cf", x"d0", x"d0", x"cf", x"d0", 
        x"cf", x"cf", x"cf", x"d0", x"d1", x"d1", x"d2", x"d0", x"d9", x"d5", x"d0", x"d1", x"d2", x"d2", x"d1", 
        x"cf", x"e9", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ed", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"f1", x"f3", x"f4", x"f3", x"ee", x"e9", x"e1", x"d7", x"c9", x"be", x"b7", x"be", x"ca", x"db", 
        x"e8", x"ef", x"f0", x"ee", x"f0", x"f1", x"ef", x"ed", x"ee", x"f1", x"f0", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f2", x"f0", x"ef", x"ee", x"ea", x"ec", x"ee", x"ef", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f4", x"f3", x"f0", x"f2", x"f5", x"f3", x"f2", x"f2", x"ea", 
        x"df", x"d4", x"c7", x"bb", x"b9", x"c8", x"e1", x"f1", x"f3", x"f1", x"f1", x"f3", x"f4", x"f2", x"f1", 
        x"f3", x"f4", x"f2", x"ef", x"ef", x"f0", x"f1", x"f3", x"ee", x"ef", x"f1", x"f2", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f5", x"f5", x"ef", x"e4", x"d8", 
        x"c6", x"bc", x"be", x"d4", x"eb", x"f3", x"f1", x"ef", x"f0", x"f0", x"ee", x"ee", x"f0", x"f4", x"f2", 
        x"f0", x"ef", x"ef", x"f0", x"f2", x"f0", x"ef", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"ee", x"ef", x"f0", x"ef", x"f1", x"f1", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"ee", 
        x"ee", x"f1", x"f2", x"f0", x"e9", x"df", x"d8", x"d9", x"d7", x"cd", x"af", x"8d", x"7d", x"83", x"8e", 
        x"8f", x"8f", x"92", x"8f", x"8e", x"93", x"93", x"8f", x"90", x"90", x"8c", x"8b", x"8c", x"93", x"9f", 
        x"ac", x"ba", x"b7", x"b5", x"88", x"32", x"20", x"0d", x"1d", x"39", x"48", x"64", x"73", x"72", x"72", 
        x"6f", x"69", x"61", x"5c", x"5b", x"5b", x"55", x"49", x"3e", x"3a", x"47", x"60", x"84", x"a9", x"c8", 
        x"d8", x"e5", x"e8", x"ea", x"e8", x"e3", x"e3", x"e4", x"e4", x"e8", x"ea", x"ec", x"e8", x"d4", x"b8", 
        x"95", x"68", x"3d", x"28", x"18", x"0b", x"0f", x"1c", x"2f", x"40", x"4d", x"50", x"4b", x"45", x"3e", 
        x"32", x"2b", x"36", x"4a", x"5b", x"5e", x"41", x"20", x"1f", x"12", x"1c", x"2c", x"21", x"2e", x"40", 
        x"38", x"32", x"32", x"35", x"37", x"3b", x"3a", x"3a", x"3a", x"3a", x"38", x"36", x"34", x"35", x"32", 
        x"89", x"89", x"89", x"89", x"89", x"89", x"88", x"86", x"87", x"89", x"89", x"88", x"87", x"87", x"87", 
        x"87", x"88", x"87", x"86", x"86", x"88", x"89", x"89", x"87", x"87", x"87", x"88", x"87", x"86", x"85", 
        x"87", x"88", x"87", x"86", x"87", x"88", x"86", x"87", x"88", x"88", x"87", x"86", x"86", x"88", x"88", 
        x"87", x"87", x"88", x"8a", x"8a", x"87", x"87", x"8a", x"89", x"89", x"89", x"88", x"8a", x"89", x"87", 
        x"87", x"88", x"89", x"89", x"89", x"8a", x"8b", x"8a", x"88", x"88", x"8a", x"8a", x"88", x"88", x"88", 
        x"89", x"89", x"8a", x"8a", x"8b", x"8a", x"8a", x"8a", x"8b", x"8c", x"8e", x"8c", x"8a", x"89", x"89", 
        x"89", x"8a", x"8b", x"8b", x"8a", x"8a", x"8a", x"8c", x"8c", x"8a", x"8a", x"8b", x"8c", x"8a", x"88", 
        x"8d", x"89", x"7d", x"a3", x"7b", x"75", x"7a", x"7b", x"7a", x"79", x"78", x"7b", x"79", x"7a", x"79", 
        x"7b", x"78", x"7d", x"75", x"79", x"79", x"42", x"63", x"79", x"41", x"3a", x"68", x"7e", x"79", x"7c", 
        x"7b", x"7c", x"7a", x"78", x"78", x"7b", x"7f", x"5d", x"36", x"38", x"3a", x"4a", x"43", x"25", x"15", 
        x"1a", x"8b", x"dd", x"d6", x"d4", x"d4", x"d4", x"da", x"d2", x"d2", x"d3", x"d2", x"d1", x"d1", x"d2", 
        x"d2", x"d4", x"d4", x"d1", x"d0", x"d1", x"d2", x"d2", x"d4", x"d5", x"d6", x"d7", x"d2", x"b7", x"97", 
        x"98", x"b3", x"cc", x"d2", x"d6", x"d5", x"d0", x"cf", x"cf", x"d0", x"d0", x"d0", x"cf", x"cf", x"d1", 
        x"d2", x"d1", x"d1", x"d2", x"cf", x"cb", x"d1", x"d0", x"da", x"d7", x"d0", x"d0", x"d0", x"d1", x"d1", 
        x"cf", x"e9", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ed", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ed", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ee", x"ef", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"ed", x"ec", x"f1", x"f1", x"ef", x"f0", x"ed", x"e7", x"df", x"d5", x"c5", x"b5", 
        x"b5", x"c3", x"d3", x"e3", x"e8", x"ed", x"f1", x"f1", x"f1", x"f0", x"ee", x"ee", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"ef", x"f0", x"ed", x"ee", x"f1", x"ef", x"f1", 
        x"f2", x"f0", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"ef", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f1", x"f1", x"f3", x"f4", x"f0", x"f1", x"f3", 
        x"f1", x"f1", x"ee", x"e1", x"d7", x"cc", x"bf", x"be", x"cd", x"e1", x"ec", x"ef", x"f1", x"f4", x"f3", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f2", x"f3", x"ee", x"f1", x"f5", x"f3", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f0", x"f0", x"f0", x"f1", x"f3", x"f4", 
        x"eb", x"e0", x"d1", x"c1", x"bd", x"c9", x"e2", x"ec", x"ef", x"ef", x"ef", x"f1", x"f4", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"ee", x"ee", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ed", x"ef", x"f0", x"ee", x"ea", x"e2", x"d9", x"d6", x"d8", x"d1", x"b6", x"94", x"82", 
        x"84", x"8f", x"93", x"92", x"8f", x"90", x"90", x"91", x"92", x"8f", x"8d", x"91", x"8f", x"8d", x"8c", 
        x"8f", x"9d", x"8b", x"92", x"65", x"0a", x"0d", x"0c", x"3e", x"69", x"65", x"62", x"63", x"5f", x"5c", 
        x"59", x"55", x"50", x"4d", x"48", x"40", x"40", x"55", x"71", x"95", x"b3", x"cf", x"dc", x"e1", x"e7", 
        x"e7", x"e5", x"e6", x"e8", x"e5", x"e4", x"e7", x"e9", x"e6", x"e0", x"c6", x"a7", x"85", x"56", x"33", 
        x"20", x"16", x"0f", x"16", x"29", x"3c", x"45", x"4c", x"4e", x"48", x"40", x"38", x"2e", x"30", x"3e", 
        x"49", x"55", x"5d", x"52", x"47", x"3a", x"25", x"24", x"26", x"12", x"18", x"2b", x"22", x"2d", x"47", 
        x"40", x"37", x"34", x"36", x"37", x"3a", x"3a", x"39", x"39", x"39", x"37", x"36", x"34", x"33", x"31", 
        x"8a", x"8a", x"8a", x"89", x"88", x"88", x"88", x"87", x"88", x"8a", x"8a", x"88", x"86", x"86", x"88", 
        x"89", x"87", x"86", x"85", x"86", x"89", x"8a", x"89", x"88", x"88", x"89", x"89", x"87", x"86", x"86", 
        x"88", x"89", x"87", x"86", x"87", x"89", x"87", x"87", x"88", x"87", x"87", x"86", x"86", x"87", x"88", 
        x"88", x"88", x"88", x"88", x"87", x"86", x"87", x"8b", x"8a", x"89", x"89", x"89", x"8a", x"88", x"87", 
        x"87", x"88", x"89", x"88", x"88", x"89", x"88", x"89", x"8b", x"8b", x"8a", x"89", x"8a", x"8b", x"8b", 
        x"8b", x"8b", x"8b", x"8b", x"8a", x"8a", x"8a", x"8a", x"8b", x"8c", x"8d", x"8c", x"8b", x"8a", x"89", 
        x"89", x"89", x"89", x"8a", x"8a", x"8a", x"8a", x"8b", x"8b", x"89", x"8a", x"8b", x"8c", x"8a", x"88", 
        x"8e", x"89", x"7d", x"a4", x"79", x"72", x"79", x"7b", x"79", x"78", x"7b", x"7e", x"7b", x"7b", x"7a", 
        x"7e", x"7c", x"7b", x"75", x"7b", x"7d", x"45", x"64", x"78", x"41", x"3a", x"68", x"7f", x"7a", x"7d", 
        x"7c", x"7b", x"7d", x"7c", x"77", x"7a", x"80", x"5f", x"38", x"31", x"27", x"20", x"16", x"12", x"09", 
        x"18", x"8a", x"dd", x"d6", x"d5", x"d6", x"d7", x"dc", x"d2", x"d1", x"d3", x"d2", x"d1", x"d1", x"d1", 
        x"d1", x"cf", x"d0", x"d5", x"d4", x"d0", x"d0", x"d2", x"d2", x"d6", x"d7", x"bc", x"94", x"90", x"b1", 
        x"cf", x"d6", x"d3", x"d1", x"d0", x"d0", x"d1", x"d1", x"d1", x"d2", x"d1", x"d1", x"d1", x"d1", x"d3", 
        x"d3", x"d2", x"d2", x"d3", x"cf", x"ca", x"d0", x"cf", x"da", x"d8", x"d2", x"d0", x"ce", x"d0", x"d1", 
        x"cf", x"e9", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", x"ee", x"ef", x"f2", x"f1", x"f0", x"f0", x"ed", x"ea", x"e5", 
        x"d8", x"c8", x"b9", x"b0", x"bb", x"cd", x"df", x"ea", x"f0", x"f2", x"f3", x"f2", x"f2", x"f0", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f2", x"f2", x"f0", x"f1", x"eb", x"ec", x"f2", x"ef", x"f0", 
        x"f1", x"f0", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"ef", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f0", x"f1", x"f1", 
        x"f0", x"f1", x"f4", x"f4", x"f0", x"ee", x"e8", x"d7", x"c2", x"b9", x"c0", x"d0", x"e6", x"ef", x"f3", 
        x"f3", x"f3", x"f5", x"f4", x"f1", x"f1", x"f1", x"f2", x"ee", x"f1", x"f4", x"f3", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f1", x"f2", x"f2", x"ec", x"dc", x"c9", x"bd", x"c4", x"d8", x"ee", x"f1", x"eb", x"eb", x"f2", x"f3", 
        x"ee", x"ed", x"f1", x"f0", x"ed", x"ed", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ee", x"ef", 
        x"f0", x"f1", x"ef", x"ef", x"f0", x"ef", x"ee", x"f0", x"ef", x"e9", x"db", x"d2", x"d9", x"d9", x"c1", 
        x"95", x"7c", x"7f", x"88", x"8d", x"92", x"90", x"8d", x"8e", x"8c", x"8c", x"90", x"92", x"93", x"8e", 
        x"88", x"89", x"9a", x"aa", x"75", x"0c", x"10", x"0d", x"46", x"75", x"67", x"55", x"50", x"4f", x"4a", 
        x"46", x"44", x"3c", x"3e", x"56", x"7d", x"ab", x"c9", x"db", x"e4", x"e9", x"eb", x"e6", x"e4", x"e5", 
        x"e3", x"e8", x"e6", x"e9", x"ec", x"e9", x"dd", x"bf", x"9e", x"7a", x"44", x"23", x"18", x"10", x"10", 
        x"18", x"2d", x"41", x"4f", x"58", x"51", x"43", x"38", x"34", x"2f", x"2f", x"3c", x"49", x"54", x"5a", 
        x"4b", x"3a", x"32", x"2e", x"31", x"2e", x"24", x"29", x"2e", x"15", x"19", x"2e", x"26", x"2d", x"4d", 
        x"46", x"3c", x"38", x"38", x"37", x"39", x"39", x"38", x"38", x"37", x"36", x"35", x"34", x"33", x"32", 
        x"8c", x"8b", x"8a", x"89", x"88", x"88", x"88", x"88", x"89", x"8a", x"8a", x"88", x"86", x"86", x"87", 
        x"89", x"88", x"86", x"85", x"86", x"89", x"8a", x"88", x"88", x"88", x"89", x"89", x"87", x"86", x"87", 
        x"88", x"88", x"87", x"87", x"89", x"8a", x"88", x"88", x"87", x"87", x"87", x"88", x"88", x"87", x"87", 
        x"88", x"89", x"88", x"88", x"87", x"85", x"85", x"89", x"89", x"88", x"88", x"88", x"89", x"87", x"87", 
        x"88", x"89", x"89", x"88", x"8a", x"8a", x"88", x"8a", x"8d", x"8d", x"8a", x"88", x"8a", x"8a", x"8a", 
        x"8a", x"8a", x"8a", x"8a", x"89", x"89", x"88", x"88", x"88", x"8a", x"8b", x"8b", x"8a", x"8a", x"8a", 
        x"8a", x"8b", x"8b", x"8a", x"8a", x"8a", x"8b", x"8b", x"8a", x"8a", x"8b", x"8b", x"8b", x"8a", x"89", 
        x"8e", x"89", x"7c", x"a2", x"7a", x"71", x"78", x"7a", x"79", x"7c", x"7d", x"7e", x"7c", x"7d", x"7b", 
        x"7e", x"7e", x"7b", x"75", x"7b", x"7d", x"46", x"64", x"79", x"42", x"3b", x"69", x"80", x"7a", x"7d", 
        x"7c", x"7d", x"7d", x"78", x"77", x"81", x"83", x"59", x"2d", x"22", x"16", x"0e", x"08", x"05", x"03", 
        x"18", x"8a", x"dd", x"d6", x"d5", x"d6", x"d7", x"dd", x"d4", x"d3", x"d4", x"d4", x"d3", x"d3", x"d3", 
        x"d3", x"d0", x"d2", x"d5", x"ce", x"cd", x"d7", x"da", x"d3", x"b9", x"94", x"8d", x"b2", x"d0", x"d5", 
        x"d3", x"d5", x"d6", x"d3", x"d0", x"d3", x"d4", x"d3", x"d3", x"d3", x"d2", x"d2", x"d3", x"d3", x"d2", 
        x"d0", x"cf", x"d1", x"d4", x"d3", x"d1", x"d0", x"ce", x"da", x"d8", x"d2", x"d1", x"ce", x"d0", x"d1", 
        x"cf", x"e9", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", 
        x"f1", x"f1", x"ef", x"ef", x"ef", x"ec", x"ec", x"ee", x"ef", x"ed", x"ec", x"ed", x"f0", x"f0", x"f1", 
        x"ef", x"ee", x"ec", x"e2", x"d2", x"be", x"ad", x"af", x"be", x"d1", x"de", x"e6", x"ee", x"ef", x"ed", 
        x"ed", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"e6", x"e8", x"ef", x"ed", x"ee", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f4", x"f3", x"f2", x"f2", x"f3", x"f3", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f0", x"ef", x"f0", x"f3", x"f4", x"f2", x"f4", x"f1", x"e9", x"d9", x"c6", x"b7", x"bc", x"c6", 
        x"d9", x"e8", x"ef", x"f2", x"f4", x"f3", x"ef", x"ef", x"ee", x"f1", x"f1", x"f2", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f5", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f2", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f3", x"f3", x"f0", x"f2", x"f5", x"f0", x"e6", x"d5", x"c9", x"c3", x"cc", x"de", x"ec", x"f1", x"f3", 
        x"ef", x"ed", x"f2", x"f4", x"f0", x"f0", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f2", 
        x"f0", x"ee", x"ef", x"f0", x"ef", x"ed", x"f0", x"f0", x"ef", x"f0", x"ef", x"eb", x"e0", x"d9", x"de", 
        x"dc", x"c2", x"a0", x"86", x"81", x"88", x"8f", x"92", x"92", x"8f", x"8f", x"8d", x"8d", x"91", x"93", 
        x"91", x"8b", x"a6", x"b6", x"81", x"13", x"16", x"13", x"40", x"73", x"68", x"54", x"48", x"3e", x"39", 
        x"47", x"6b", x"94", x"bc", x"d7", x"e4", x"e9", x"e8", x"e7", x"e9", x"e4", x"e3", x"e2", x"e8", x"ec", 
        x"e5", x"e8", x"df", x"d0", x"ac", x"85", x"5b", x"2f", x"19", x"15", x"13", x"1a", x"29", x"3e", x"4e", 
        x"54", x"53", x"4a", x"44", x"3b", x"2d", x"32", x"3c", x"40", x"41", x"42", x"45", x"40", x"34", x"2d", 
        x"2d", x"2e", x"2d", x"29", x"2a", x"29", x"26", x"29", x"31", x"17", x"16", x"2d", x"29", x"2d", x"50", 
        x"4b", x"41", x"3c", x"39", x"35", x"35", x"38", x"38", x"37", x"36", x"34", x"34", x"35", x"34", x"33", 
        x"8a", x"8a", x"8a", x"89", x"89", x"89", x"89", x"89", x"89", x"88", x"88", x"89", x"88", x"87", x"87", 
        x"88", x"89", x"88", x"87", x"87", x"88", x"89", x"88", x"87", x"87", x"88", x"88", x"87", x"87", x"89", 
        x"88", x"88", x"87", x"88", x"89", x"8a", x"88", x"88", x"88", x"88", x"88", x"89", x"8a", x"89", x"89", 
        x"89", x"89", x"89", x"88", x"88", x"86", x"86", x"89", x"89", x"89", x"8a", x"88", x"8a", x"89", x"88", 
        x"88", x"8a", x"8b", x"8b", x"8c", x"8b", x"89", x"8b", x"8c", x"8b", x"8a", x"8a", x"88", x"88", x"88", 
        x"89", x"89", x"8a", x"8a", x"8a", x"8a", x"8b", x"8b", x"8b", x"8a", x"8a", x"8a", x"8a", x"8a", x"8b", 
        x"8a", x"8a", x"8a", x"8b", x"8b", x"8b", x"8c", x"8b", x"8b", x"8b", x"8c", x"8b", x"8b", x"8a", x"89", 
        x"8e", x"89", x"7c", x"a4", x"7d", x"74", x"79", x"7a", x"78", x"7b", x"7b", x"7b", x"7b", x"7d", x"79", 
        x"7a", x"7c", x"7a", x"75", x"7a", x"7b", x"45", x"63", x"77", x"41", x"3b", x"6a", x"81", x"7b", x"7d", 
        x"7a", x"7a", x"7a", x"7f", x"83", x"76", x"54", x"31", x"19", x"13", x"0b", x"04", x"01", x"03", x"04", 
        x"17", x"8a", x"dd", x"d5", x"d3", x"d5", x"d6", x"dc", x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d3", 
        x"d2", x"d1", x"d1", x"d1", x"d2", x"dd", x"d3", x"b7", x"94", x"88", x"a7", x"d4", x"d9", x"d1", x"cf", 
        x"d2", x"d2", x"d4", x"d3", x"d0", x"d2", x"d0", x"d1", x"d0", x"d1", x"d3", x"d4", x"d6", x"d5", x"d4", 
        x"d1", x"d0", x"d2", x"d2", x"d0", x"d0", x"d0", x"cf", x"da", x"d7", x"d3", x"d4", x"d0", x"d0", x"d1", 
        x"cf", x"e9", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ed", x"ed", x"ef", x"f1", 
        x"f1", x"f0", x"ee", x"ed", x"ef", x"f0", x"ee", x"ed", x"ef", x"ef", x"ef", x"ee", x"f0", x"ef", x"ee", 
        x"ed", x"ef", x"f0", x"ed", x"f0", x"f2", x"ea", x"da", x"c6", x"b7", x"b1", x"b8", x"c7", x"d6", x"e2", 
        x"eb", x"f1", x"f5", x"f4", x"f2", x"f1", x"f0", x"f1", x"f0", x"f1", x"e7", x"e8", x"f2", x"ee", x"ef", 
        x"f1", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f1", x"f1", x"f1", 
        x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f3", x"f2", x"f1", x"f2", x"f3", x"f1", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f2", x"f3", x"f5", x"f4", x"f3", x"ea", x"d3", x"bd", 
        x"b4", x"ba", x"c8", x"d7", x"e5", x"f0", x"f4", x"f0", x"ed", x"f1", x"f2", x"f3", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f3", x"f4", x"f5", x"f5", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f4", x"f5", x"f4", x"f1", 
        x"f1", x"f1", x"ee", x"ef", x"f2", x"f3", x"f2", x"f4", x"f0", x"e1", x"cd", x"c2", x"c5", x"d7", x"e4", 
        x"ea", x"f0", x"f4", x"f1", x"ee", x"f1", x"f4", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", x"f0", 
        x"ee", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"ec", x"eb", x"ee", x"f0", 
        x"ef", x"ed", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", x"f1", x"ed", x"ec", x"f0", x"f2", x"ee", x"e4", 
        x"db", x"dd", x"df", x"cf", x"a7", x"8b", x"82", x"89", x"8e", x"8b", x"90", x"91", x"92", x"8e", x"8e", 
        x"91", x"8c", x"ad", x"b9", x"8a", x"1d", x"16", x"13", x"3d", x"6d", x"63", x"53", x"5d", x"7f", x"a6", 
        x"cc", x"e4", x"ec", x"ed", x"e9", x"e6", x"e7", x"e7", x"e6", x"e8", x"ea", x"ed", x"e9", x"e4", x"da", 
        x"bf", x"97", x"6e", x"41", x"18", x"10", x"19", x"1d", x"26", x"33", x"47", x"55", x"5e", x"5e", x"4d", 
        x"37", x"30", x"29", x"2a", x"31", x"3a", x"51", x"50", x"37", x"2c", x"2a", x"2b", x"2d", x"2f", x"2b", 
        x"27", x"2a", x"26", x"28", x"2d", x"27", x"24", x"28", x"36", x"1b", x"13", x"27", x"28", x"2c", x"54", 
        x"50", x"48", x"42", x"3e", x"37", x"35", x"36", x"37", x"37", x"36", x"35", x"34", x"33", x"33", x"32", 
        x"8a", x"8a", x"8b", x"8a", x"8a", x"8a", x"8a", x"8a", x"89", x"89", x"89", x"89", x"89", x"88", x"87", 
        x"88", x"89", x"89", x"89", x"88", x"87", x"87", x"88", x"88", x"87", x"88", x"88", x"86", x"87", x"8a", 
        x"89", x"88", x"87", x"88", x"89", x"89", x"88", x"89", x"8a", x"89", x"89", x"8a", x"8a", x"8a", x"89", 
        x"89", x"88", x"88", x"89", x"8a", x"88", x"87", x"89", x"8a", x"8a", x"8b", x"8b", x"8b", x"8b", x"8a", 
        x"89", x"8a", x"8b", x"8b", x"8b", x"8a", x"8a", x"8b", x"8b", x"89", x"8b", x"8d", x"8a", x"8a", x"8b", 
        x"8b", x"8b", x"8b", x"8c", x"8b", x"8d", x"8e", x"8e", x"8d", x"8b", x"8a", x"8b", x"8b", x"8b", x"8b", 
        x"8b", x"8b", x"8a", x"8a", x"8b", x"8b", x"8b", x"8b", x"8c", x"8c", x"8c", x"8c", x"8c", x"8b", x"8b", 
        x"8f", x"89", x"7e", x"a6", x"7d", x"73", x"7b", x"7c", x"79", x"7b", x"7a", x"79", x"79", x"7a", x"78", 
        x"79", x"7a", x"79", x"73", x"79", x"7d", x"47", x"63", x"75", x"40", x"3b", x"67", x"80", x"7c", x"7d", 
        x"7c", x"80", x"85", x"78", x"58", x"35", x"1a", x"11", x"0d", x"06", x"05", x"04", x"03", x"05", x"06", 
        x"18", x"87", x"db", x"d4", x"d2", x"d4", x"d5", x"dd", x"d1", x"d2", x"d4", x"d2", x"d1", x"d1", x"d2", 
        x"d1", x"d4", x"d6", x"d8", x"d3", x"b9", x"9d", x"8f", x"a7", x"c8", x"d5", x"d3", x"d2", x"d1", x"d0", 
        x"d4", x"d3", x"d4", x"d7", x"d3", x"d1", x"d2", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", 
        x"d0", x"d0", x"d2", x"d2", x"d0", x"d1", x"d1", x"d1", x"da", x"d8", x"d3", x"d5", x"d2", x"d0", x"d1", 
        x"cf", x"e8", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ee", x"ef", x"f0", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f1", x"f0", x"ef", x"f0", x"ee", x"ed", x"ee", 
        x"ef", x"ef", x"ee", x"f0", x"ef", x"ef", x"f0", x"f1", x"ef", x"eb", x"df", x"d0", x"c0", x"ba", x"be", 
        x"c7", x"ce", x"d9", x"e3", x"eb", x"f1", x"f2", x"f1", x"ef", x"f1", x"ea", x"eb", x"f4", x"ee", x"f1", 
        x"f2", x"ef", x"ef", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f1", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f1", 
        x"ef", x"f1", x"f2", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", 
        x"e7", x"d5", x"c1", x"b6", x"bc", x"c8", x"d5", x"e2", x"ef", x"f5", x"f5", x"f3", x"f4", x"f3", x"f4", 
        x"f4", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f5", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f3", x"f2", x"f3", x"f4", x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"ef", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"e9", x"da", x"cd", x"ca", 
        x"d1", x"de", x"e7", x"ed", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f0", 
        x"ee", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"ef", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f0", 
        x"ee", x"ed", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f1", x"ef", x"ef", 
        x"f0", x"e9", x"de", x"dd", x"e0", x"d1", x"b1", x"93", x"88", x"84", x"88", x"90", x"95", x"90", x"8e", 
        x"91", x"8c", x"b0", x"ba", x"87", x"19", x"1f", x"31", x"56", x"83", x"9e", x"b8", x"cd", x"df", x"e8", 
        x"e8", x"e9", x"e7", x"e6", x"e8", x"ea", x"ea", x"eb", x"ec", x"e8", x"da", x"cb", x"aa", x"84", x"62", 
        x"3a", x"1f", x"17", x"0a", x"20", x"3b", x"54", x"65", x"6a", x"5d", x"56", x"4d", x"49", x"4b", x"3e", 
        x"2d", x"2e", x"2e", x"2e", x"30", x"2f", x"2e", x"2d", x"2a", x"2d", x"30", x"2c", x"28", x"2a", x"2b", 
        x"2a", x"2a", x"27", x"29", x"2a", x"27", x"27", x"28", x"38", x"1f", x"13", x"27", x"29", x"2c", x"55", 
        x"56", x"4d", x"47", x"42", x"3b", x"39", x"38", x"37", x"37", x"37", x"36", x"34", x"33", x"32", x"32", 
        x"8c", x"89", x"8c", x"8b", x"89", x"8b", x"8a", x"8a", x"8a", x"8a", x"8a", x"8a", x"89", x"88", x"8a", 
        x"8a", x"88", x"88", x"89", x"89", x"88", x"85", x"87", x"8a", x"89", x"8b", x"8a", x"86", x"87", x"8b", 
        x"8b", x"89", x"85", x"89", x"89", x"89", x"88", x"8a", x"8a", x"89", x"88", x"89", x"89", x"86", x"87", 
        x"88", x"88", x"88", x"8a", x"8b", x"8b", x"88", x"88", x"89", x"87", x"89", x"8a", x"89", x"8a", x"8a", 
        x"8a", x"8a", x"8a", x"8a", x"89", x"89", x"8a", x"8b", x"8a", x"8a", x"8c", x"8c", x"8a", x"8b", x"8c", 
        x"8a", x"88", x"88", x"89", x"8c", x"8c", x"8b", x"8a", x"8a", x"89", x"88", x"8a", x"8b", x"8b", x"8c", 
        x"8c", x"8d", x"8d", x"8a", x"89", x"89", x"89", x"8a", x"8c", x"8d", x"8c", x"8d", x"8e", x"8c", x"8c", 
        x"90", x"89", x"80", x"a7", x"7b", x"71", x"7b", x"7e", x"7a", x"7c", x"7d", x"7b", x"78", x"78", x"7a", 
        x"7b", x"7a", x"7c", x"73", x"78", x"7e", x"46", x"63", x"76", x"44", x"3b", x"63", x"7f", x"7e", x"82", 
        x"86", x"80", x"67", x"3b", x"1c", x"12", x"0c", x"04", x"03", x"05", x"06", x"05", x"07", x"14", x"2a", 
        x"35", x"7e", x"db", x"d6", x"d1", x"d3", x"d4", x"df", x"d4", x"d2", x"d3", x"d2", x"d1", x"d2", x"d0", 
        x"d0", x"db", x"d5", x"bb", x"a0", x"86", x"9f", x"cd", x"da", x"d4", x"d0", x"d0", x"d1", x"d1", x"d2", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d3", x"d3", x"d2", x"d1", x"d1", x"d0", x"cf", x"d0", x"d1", 
        x"d0", x"d0", x"d0", x"d0", x"d1", x"d2", x"d0", x"d2", x"d9", x"da", x"d2", x"d4", x"d2", x"cf", x"d0", 
        x"d0", x"e6", x"f0", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f4", x"f3", x"ed", x"df", 
        x"cc", x"bd", x"b8", x"ba", x"c3", x"cf", x"dc", x"e9", x"ef", x"f3", x"ed", x"e8", x"f0", x"ee", x"f2", 
        x"f1", x"ef", x"ef", x"f1", x"ee", x"f2", x"f3", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f2", 
        x"f4", x"f5", x"f3", x"eb", x"d4", x"be", x"b3", x"bb", x"d2", x"dc", x"e6", x"f1", x"f4", x"f5", x"f4", 
        x"f3", x"f2", x"f2", x"f3", x"f3", x"f0", x"f2", x"f5", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", 
        x"f4", x"f5", x"f5", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"e7", 
        x"d7", x"cb", x"c9", x"d3", x"e3", x"ed", x"f3", x"f4", x"f1", x"ee", x"ef", x"f2", x"f2", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f4", x"f3", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f3", 
        x"f0", x"ee", x"ef", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f0", x"ef", x"ef", x"ef", 
        x"f1", x"f3", x"f2", x"e9", x"e0", x"e1", x"e6", x"db", x"bc", x"9d", x"85", x"80", x"85", x"8e", x"93", 
        x"8f", x"81", x"a2", x"b2", x"93", x"54", x"79", x"a6", x"ce", x"e2", x"ed", x"ee", x"e9", x"e6", x"e3", 
        x"e6", x"e8", x"ea", x"ea", x"ec", x"ef", x"e7", x"d9", x"c0", x"99", x"72", x"4e", x"24", x"13", x"1d", 
        x"2a", x"40", x"35", x"13", x"57", x"83", x"82", x"80", x"70", x"47", x"3a", x"3d", x"3e", x"45", x"3d", 
        x"2e", x"2a", x"2d", x"2b", x"28", x"2a", x"2a", x"2b", x"2c", x"2b", x"2b", x"2a", x"28", x"28", x"2a", 
        x"2a", x"2b", x"2a", x"2a", x"2a", x"2b", x"28", x"24", x"31", x"1c", x"10", x"29", x"30", x"2c", x"56", 
        x"5b", x"51", x"48", x"45", x"40", x"3e", x"3b", x"38", x"36", x"37", x"37", x"35", x"34", x"31", x"32", 
        x"8c", x"8a", x"8c", x"8b", x"89", x"8a", x"89", x"8b", x"8b", x"89", x"88", x"88", x"89", x"8a", x"8b", 
        x"8a", x"89", x"88", x"87", x"88", x"8a", x"89", x"88", x"8a", x"8b", x"8b", x"8a", x"89", x"8a", x"89", 
        x"89", x"89", x"88", x"89", x"89", x"8a", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"89", x"8a", 
        x"8a", x"89", x"89", x"8a", x"8b", x"8c", x"89", x"89", x"89", x"87", x"88", x"88", x"88", x"8a", x"89", 
        x"88", x"88", x"89", x"8a", x"8a", x"8a", x"8b", x"8b", x"8a", x"8a", x"8b", x"8b", x"8a", x"8b", x"8b", 
        x"8b", x"8a", x"8a", x"8b", x"8b", x"8a", x"8a", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8c", 
        x"8c", x"8c", x"8c", x"8a", x"8a", x"8b", x"8b", x"8c", x"8c", x"8c", x"8c", x"8d", x"8e", x"8b", x"8b", 
        x"8e", x"89", x"80", x"a6", x"7f", x"72", x"7a", x"7e", x"7b", x"79", x"78", x"7b", x"7b", x"79", x"7a", 
        x"7d", x"7e", x"7c", x"77", x"7c", x"7d", x"45", x"60", x"74", x"43", x"3d", x"67", x"86", x"87", x"7f", 
        x"62", x"44", x"2d", x"1e", x"12", x"07", x"04", x"05", x"04", x"05", x"08", x"1e", x"40", x"59", x"6c", 
        x"5b", x"76", x"d7", x"d5", x"d2", x"d6", x"d5", x"dd", x"d1", x"cf", x"d1", x"d5", x"d3", x"cf", x"d8", 
        x"d6", x"b3", x"95", x"93", x"a8", x"c9", x"d4", x"d3", x"cf", x"cf", x"d0", x"d3", x"d3", x"d0", x"d0", 
        x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d3", x"d2", x"d1", x"d1", x"d0", x"cf", x"cf", x"d0", x"d1", 
        x"d1", x"d0", x"d0", x"d0", x"d1", x"d1", x"d1", x"d2", x"d8", x"d9", x"d0", x"d3", x"d2", x"d0", x"d1", 
        x"d0", x"e5", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", 
        x"ee", x"eb", x"e4", x"d9", x"cd", x"c1", x"ba", x"ba", x"bd", x"c6", x"de", x"e7", x"f1", x"f4", x"f2", 
        x"f0", x"f4", x"f2", x"f1", x"f1", x"f2", x"ee", x"ee", x"f3", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"ef", x"ea", x"dc", x"d2", x"cb", x"cb", x"c8", x"cf", x"df", x"eb", 
        x"f3", x"f3", x"f2", x"f1", x"f3", x"f2", x"f0", x"f4", x"f3", x"f1", x"f1", x"f3", x"f4", x"f4", x"f4", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f4", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"ef", x"f3", 
        x"f4", x"ed", x"e3", x"d7", x"cd", x"cb", x"d2", x"e0", x"ec", x"f2", x"f3", x"f0", x"ef", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f2", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f3", 
        x"f0", x"ee", x"ef", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f3", x"f2", x"f1", x"f0", x"ed", x"e8", x"e4", x"e1", x"dd", x"c7", x"a9", x"90", x"7c", x"7b", 
        x"88", x"8e", x"b2", x"cc", x"d6", x"d1", x"e5", x"ea", x"eb", x"ea", x"e4", x"e5", x"e8", x"e7", x"e9", 
        x"ec", x"ed", x"e9", x"d6", x"c1", x"a1", x"73", x"52", x"36", x"1e", x"1f", x"31", x"42", x"55", x"67", 
        x"6d", x"6f", x"48", x"12", x"47", x"78", x"7a", x"7b", x"73", x"4b", x"3c", x"3f", x"3f", x"42", x"37", 
        x"2e", x"29", x"2a", x"2b", x"2c", x"2d", x"2a", x"28", x"29", x"29", x"29", x"2a", x"2a", x"2a", x"2b", 
        x"2d", x"2c", x"2b", x"29", x"28", x"2b", x"27", x"21", x"2d", x"1c", x"12", x"2a", x"32", x"2c", x"56", 
        x"60", x"55", x"4e", x"4b", x"46", x"43", x"3d", x"39", x"38", x"38", x"38", x"36", x"34", x"31", x"2e", 
        x"8c", x"8b", x"8b", x"8a", x"89", x"89", x"88", x"8b", x"8b", x"89", x"88", x"88", x"89", x"8b", x"8b", 
        x"8b", x"8a", x"88", x"87", x"88", x"8b", x"8c", x"89", x"88", x"8c", x"8b", x"8a", x"8c", x"8b", x"88", 
        x"87", x"8a", x"8a", x"8a", x"88", x"8b", x"8a", x"89", x"88", x"89", x"8a", x"8a", x"88", x"8a", x"8a", 
        x"8a", x"89", x"89", x"8a", x"8b", x"8b", x"88", x"89", x"89", x"87", x"8a", x"8a", x"8a", x"8b", x"89", 
        x"88", x"88", x"89", x"8b", x"8b", x"8b", x"8c", x"8b", x"8a", x"8a", x"8b", x"8b", x"8b", x"8b", x"8b", 
        x"8b", x"8b", x"8c", x"8d", x"8b", x"8a", x"8a", x"8b", x"8b", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", 
        x"8c", x"8c", x"8c", x"8b", x"8b", x"8c", x"8d", x"8d", x"8c", x"8c", x"8b", x"8c", x"8e", x"8d", x"8d", 
        x"8f", x"89", x"7f", x"a6", x"7e", x"71", x"7a", x"7c", x"7b", x"7b", x"78", x"7c", x"7d", x"7a", x"7b", 
        x"7d", x"7d", x"7c", x"84", x"7d", x"7a", x"43", x"5c", x"72", x"41", x"40", x"6f", x"81", x"65", x"4a", 
        x"2e", x"1c", x"15", x"0e", x"07", x"03", x"04", x"06", x"05", x"08", x"16", x"4b", x"7b", x"76", x"74", 
        x"59", x"78", x"d8", x"d4", x"d4", x"d6", x"d5", x"de", x"d5", x"d0", x"d1", x"d5", x"d8", x"d4", x"bd", 
        x"9a", x"8e", x"a4", x"c2", x"d3", x"d5", x"cf", x"cc", x"cd", x"ce", x"d0", x"d2", x"d2", x"cf", x"d1", 
        x"d5", x"d5", x"d5", x"d5", x"d5", x"d5", x"d4", x"d3", x"d3", x"d2", x"d2", x"d1", x"d1", x"d1", x"d2", 
        x"d2", x"d1", x"d1", x"d1", x"d0", x"d0", x"d1", x"d2", x"d8", x"d8", x"d0", x"d3", x"d2", x"d1", x"d2", 
        x"cf", x"e5", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f2", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"eb", x"de", x"cf", x"c4", x"bc", x"c9", x"c5", x"c0", x"ce", x"df", 
        x"e9", x"f1", x"f4", x"f3", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"f1", x"f2", x"f1", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f4", x"ef", x"e9", x"e1", x"d2", x"ca", x"c5", x"c7", 
        x"d1", x"e0", x"ea", x"f1", x"f6", x"f4", x"f2", x"f3", x"f3", x"f2", x"f3", x"f4", x"f3", x"f3", x"f3", 
        x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f4", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", 
        x"f1", x"f2", x"f4", x"f2", x"e7", x"d9", x"cf", x"c9", x"c9", x"d3", x"e3", x"ee", x"f0", x"f1", x"f3", 
        x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f3", 
        x"f0", x"ee", x"ef", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"ef", x"ea", x"e7", x"e3", x"de", x"d0", x"b2", x"a8", 
        x"be", x"d2", x"e0", x"e9", x"eb", x"ea", x"e8", x"e4", x"e5", x"e9", x"e9", x"ec", x"ee", x"e9", x"df", 
        x"cd", x"b2", x"8b", x"5f", x"45", x"30", x"1b", x"23", x"37", x"48", x"5a", x"6d", x"6e", x"65", x"5c", 
        x"50", x"46", x"31", x"0b", x"36", x"73", x"7f", x"80", x"7e", x"55", x"3d", x"3f", x"3f", x"40", x"37", 
        x"2c", x"27", x"28", x"2a", x"2b", x"2a", x"2a", x"28", x"28", x"29", x"28", x"29", x"2a", x"28", x"28", 
        x"2b", x"2a", x"28", x"26", x"27", x"29", x"26", x"1f", x"2b", x"1d", x"12", x"25", x"31", x"2a", x"54", 
        x"64", x"59", x"53", x"4d", x"46", x"43", x"3f", x"3e", x"3c", x"3a", x"37", x"36", x"34", x"34", x"31", 
        x"8d", x"8c", x"8b", x"8a", x"89", x"88", x"88", x"8a", x"8a", x"89", x"89", x"89", x"89", x"8a", x"8a", 
        x"8b", x"8b", x"8b", x"89", x"8a", x"8b", x"8c", x"89", x"88", x"8b", x"89", x"88", x"8a", x"8a", x"88", 
        x"87", x"8a", x"8c", x"8a", x"88", x"8c", x"8b", x"8a", x"89", x"8a", x"8b", x"8b", x"89", x"89", x"89", 
        x"88", x"89", x"89", x"8a", x"8b", x"8c", x"8a", x"8b", x"8b", x"89", x"8b", x"8b", x"8a", x"8b", x"8a", 
        x"8a", x"8a", x"8a", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8c", x"8b", x"8b", 
        x"8b", x"8c", x"8d", x"8d", x"8c", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8c", x"8d", x"8d", x"8d", 
        x"8c", x"8c", x"8c", x"8d", x"8d", x"8d", x"8c", x"8c", x"8c", x"8c", x"8b", x"8b", x"8e", x"8e", x"8e", 
        x"8f", x"89", x"7e", x"9f", x"78", x"71", x"7d", x"7e", x"7f", x"80", x"7a", x"7b", x"7c", x"7c", x"7e", 
        x"7e", x"7a", x"7c", x"91", x"7d", x"78", x"3e", x"5b", x"75", x"46", x"47", x"51", x"42", x"32", x"25", 
        x"14", x"0a", x"07", x"04", x"03", x"05", x"04", x"09", x"11", x"23", x"35", x"65", x"7e", x"68", x"70", 
        x"5e", x"78", x"da", x"d6", x"d4", x"d6", x"d6", x"dd", x"d2", x"d3", x"d7", x"df", x"c6", x"91", x"87", 
        x"a2", x"c5", x"d5", x"d1", x"d0", x"cd", x"ce", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d1", x"d2", 
        x"d5", x"d5", x"d5", x"d5", x"d5", x"d5", x"d4", x"d2", x"d1", x"d1", x"d0", x"d0", x"cf", x"d0", x"d2", 
        x"d3", x"d2", x"d2", x"d1", x"d0", x"d0", x"d1", x"d3", x"d8", x"d8", x"d0", x"d4", x"d3", x"d2", x"d2", 
        x"cf", x"e4", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ee", x"f0", x"f0", x"ef", x"f0", x"f2", x"f2", x"ef", x"e7", x"e6", x"d8", x"c8", x"b3", x"a4", 
        x"a6", x"b7", x"d6", x"eb", x"f6", x"f4", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f4", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f1", 
        x"f0", x"f0", x"f2", x"f3", x"f0", x"f1", x"f2", x"f2", x"ed", x"f0", x"f2", x"f1", x"ee", x"e5", x"d9", 
        x"cb", x"c0", x"bd", x"cf", x"e1", x"f1", x"f6", x"f3", x"ef", x"f0", x"f2", x"f3", x"f2", x"f2", x"f1", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", 
        x"ee", x"f2", x"f3", x"f3", x"f1", x"f1", x"ef", x"e9", x"db", x"ca", x"bd", x"c3", x"db", x"f1", x"f5", 
        x"f3", x"f1", x"f4", x"f5", x"f3", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f3", x"f2", x"f0", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f3", 
        x"f0", x"ee", x"ef", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f3", x"ef", x"ee", x"ef", x"f1", x"f1", x"ef", x"ed", x"e2", x"e7", x"ed", x"ed", 
        x"ec", x"e8", x"eb", x"eb", x"e6", x"e7", x"e7", x"ec", x"ef", x"f3", x"f2", x"e1", x"c7", x"a1", x"6d", 
        x"42", x"2a", x"19", x"16", x"27", x"45", x"5f", x"6d", x"74", x"6f", x"62", x"50", x"39", x"2c", x"29", 
        x"29", x"31", x"31", x"1a", x"37", x"7a", x"89", x"81", x"89", x"61", x"40", x"3f", x"3e", x"40", x"39", 
        x"2c", x"27", x"26", x"27", x"27", x"26", x"29", x"28", x"27", x"28", x"27", x"27", x"29", x"27", x"25", 
        x"27", x"26", x"24", x"24", x"26", x"2a", x"28", x"20", x"2a", x"20", x"11", x"21", x"33", x"2b", x"53", 
        x"6b", x"5d", x"55", x"4d", x"48", x"47", x"41", x"3e", x"3d", x"3d", x"3d", x"3b", x"38", x"35", x"2c", 
        x"8c", x"8c", x"8b", x"8a", x"8a", x"88", x"89", x"88", x"89", x"8a", x"8b", x"8b", x"8a", x"89", x"89", 
        x"89", x"8a", x"8a", x"8a", x"8a", x"8b", x"8b", x"8a", x"89", x"8a", x"88", x"87", x"88", x"89", x"89", 
        x"89", x"8a", x"8a", x"8a", x"89", x"8b", x"89", x"88", x"88", x"88", x"89", x"89", x"88", x"88", x"88", 
        x"88", x"89", x"8a", x"8a", x"8a", x"8b", x"8a", x"8b", x"8c", x"8a", x"8c", x"8d", x"8b", x"8b", x"8b", 
        x"8b", x"8b", x"8b", x"8a", x"8a", x"8b", x"8b", x"8b", x"8c", x"8c", x"8c", x"8c", x"8c", x"8b", x"8b", 
        x"8b", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8b", x"8b", x"8b", x"8b", x"8c", x"8c", x"8c", x"8c", 
        x"8c", x"8c", x"8c", x"8d", x"8e", x"8d", x"8b", x"8b", x"8c", x"8d", x"8d", x"8e", x"8e", x"8d", x"8c", 
        x"8d", x"8b", x"7f", x"9c", x"7e", x"74", x"7c", x"7e", x"7e", x"7a", x"7d", x"7c", x"7b", x"7d", x"7e", 
        x"7c", x"79", x"7c", x"8c", x"7b", x"7a", x"46", x"5f", x"70", x"3e", x"31", x"30", x"23", x"15", x"0b", 
        x"04", x"05", x"05", x"05", x"0a", x"18", x"42", x"4b", x"35", x"3c", x"3c", x"62", x"7f", x"70", x"72", 
        x"58", x"79", x"d6", x"d5", x"d4", x"d4", x"d7", x"e1", x"da", x"d2", x"c2", x"9d", x"8c", x"a8", x"c7", 
        x"d2", x"d3", x"cd", x"cd", x"d0", x"cf", x"cf", x"d0", x"d1", x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", 
        x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d3", x"d2", x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"d2", 
        x"d3", x"d2", x"d2", x"d2", x"d0", x"d0", x"d0", x"d2", x"d8", x"d8", x"d0", x"d3", x"d2", x"d2", x"d2", 
        x"cf", x"e4", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"f0", x"f1", x"f0", x"f1", x"f0", x"e8", x"ed", x"e8", x"de", 
        x"d2", x"c2", x"ad", x"a6", x"ac", x"c3", x"da", x"e8", x"ed", x"f0", x"f1", x"f3", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f0", x"f1", x"f1", 
        x"f0", x"f0", x"f1", x"f3", x"f3", x"f3", x"f2", x"f3", x"ed", x"ef", x"f0", x"f2", x"f2", x"f2", x"f3", 
        x"f0", x"e8", x"e0", x"d2", x"c5", x"c3", x"ce", x"de", x"ec", x"f2", x"f3", x"f4", x"f4", x"f3", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f0", x"ee", x"ee", x"f0", x"f1", x"f0", x"f2", x"f4", x"ef", x"ec", x"e4", x"d5", x"c7", x"c1", x"cc", 
        x"de", x"ed", x"f0", x"ef", x"f1", x"f3", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f3", 
        x"f0", x"ee", x"ef", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f1", x"ef", x"eb", x"eb", x"eb", x"ec", 
        x"ed", x"e9", x"e6", x"e9", x"ee", x"ed", x"e6", x"df", x"c9", x"a9", x"88", x"57", x"34", x"27", x"1f", 
        x"25", x"3c", x"55", x"69", x"71", x"71", x"69", x"54", x"45", x"3e", x"34", x"2e", x"2d", x"2d", x"2b", 
        x"2a", x"30", x"31", x"24", x"39", x"7c", x"91", x"8d", x"8f", x"69", x"45", x"45", x"41", x"40", x"39", 
        x"2d", x"29", x"25", x"25", x"29", x"28", x"28", x"26", x"25", x"26", x"26", x"27", x"28", x"28", x"27", 
        x"26", x"25", x"25", x"25", x"27", x"2a", x"29", x"1f", x"2a", x"24", x"14", x"21", x"3c", x"33", x"4f", 
        x"6b", x"5e", x"5a", x"53", x"4d", x"4b", x"49", x"43", x"3e", x"38", x"2f", x"26", x"23", x"23", x"32", 
        x"8b", x"8d", x"8a", x"8a", x"8b", x"89", x"89", x"88", x"88", x"89", x"8b", x"8b", x"8a", x"89", x"89", 
        x"89", x"89", x"89", x"8a", x"8b", x"8b", x"8a", x"8a", x"8a", x"89", x"8a", x"8a", x"89", x"8a", x"8b", 
        x"8b", x"8a", x"88", x"8a", x"8a", x"8a", x"88", x"89", x"89", x"88", x"88", x"88", x"88", x"89", x"8a", 
        x"8a", x"8b", x"8b", x"8a", x"89", x"8a", x"88", x"89", x"8a", x"89", x"8b", x"8c", x"8b", x"8b", x"8b", 
        x"8b", x"8b", x"8b", x"8b", x"8c", x"8c", x"8b", x"8b", x"8c", x"8c", x"8b", x"8b", x"8c", x"8b", x"8b", 
        x"8c", x"8c", x"8b", x"8a", x"8b", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8b", x"8b", x"8b", x"8c", 
        x"8c", x"8c", x"8c", x"8d", x"8c", x"8c", x"8b", x"8c", x"8c", x"8c", x"8e", x"8f", x"8e", x"8c", x"8b", 
        x"8d", x"8e", x"81", x"98", x"7d", x"72", x"7b", x"7d", x"7f", x"7b", x"7b", x"79", x"7b", x"7e", x"7d", 
        x"7b", x"7c", x"7e", x"8d", x"84", x"7f", x"4f", x"4a", x"4e", x"33", x"23", x"15", x"0b", x"08", x"06", 
        x"03", x"05", x"07", x"14", x"36", x"65", x"8c", x"6f", x"3d", x"3e", x"3b", x"62", x"81", x"75", x"78", 
        x"61", x"7b", x"d7", x"d4", x"d1", x"d5", x"dc", x"d7", x"c7", x"a0", x"81", x"a3", x"c9", x"d0", x"d1", 
        x"d1", x"d3", x"d2", x"d0", x"cb", x"cd", x"d3", x"d1", x"d0", x"d1", x"d2", x"d2", x"d2", x"d1", x"d2", 
        x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d2", x"d2", x"d2", x"d1", x"d1", 
        x"d2", x"d2", x"d3", x"d3", x"d2", x"d1", x"d0", x"d2", x"d8", x"d9", x"d1", x"d3", x"d2", x"d3", x"d3", 
        x"cf", x"e3", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", 
        x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"f2", x"f2", x"ef", x"ee", x"ef", x"ee", x"f0", x"f2", x"f4", x"ed", x"f1", 
        x"f2", x"f0", x"e8", x"dd", x"cc", x"af", x"9f", x"a5", x"b6", x"d2", x"e1", x"ed", x"f0", x"f1", x"f1", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f2", x"f3", x"f1", x"f0", x"ef", x"eb", x"ee", x"f3", x"f1", x"f2", x"f2", x"f0", 
        x"ef", x"f1", x"f4", x"f3", x"eb", x"e0", x"cd", x"be", x"c6", x"d6", x"e4", x"ed", x"f4", x"f6", x"f4", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", 
        x"ef", x"ef", x"f1", x"f4", x"f5", x"f2", x"f0", x"f1", x"f2", x"f2", x"f2", x"ef", x"ea", x"df", x"ca", 
        x"c0", x"c1", x"d6", x"e9", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f3", 
        x"f0", x"ee", x"ef", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"ee", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"eb", x"e7", x"ea", x"ec", 
        x"ea", x"eb", x"ed", x"e7", x"df", x"c1", x"9b", x"70", x"40", x"25", x"1c", x"1a", x"25", x"41", x"5f", 
        x"6f", x"78", x"73", x"64", x"54", x"45", x"39", x"34", x"36", x"34", x"30", x"2e", x"31", x"30", x"2e", 
        x"2e", x"2f", x"2c", x"26", x"39", x"79", x"93", x"96", x"95", x"72", x"4c", x"4c", x"47", x"43", x"3c", 
        x"2c", x"29", x"26", x"25", x"29", x"27", x"26", x"26", x"25", x"25", x"26", x"27", x"27", x"28", x"28", 
        x"27", x"27", x"26", x"25", x"25", x"27", x"25", x"1d", x"29", x"28", x"16", x"1f", x"40", x"3a", x"5a", 
        x"76", x"63", x"61", x"5b", x"50", x"47", x"3a", x"2c", x"21", x"1d", x"25", x"41", x"67", x"93", x"b3", 
        x"8b", x"8d", x"8b", x"8b", x"8c", x"89", x"8a", x"89", x"89", x"8a", x"8a", x"8a", x"8b", x"8a", x"8b", 
        x"8a", x"88", x"88", x"89", x"8b", x"8b", x"8a", x"8a", x"8b", x"8a", x"8c", x"8c", x"8b", x"8c", x"8c", 
        x"8c", x"89", x"87", x"8a", x"8b", x"8a", x"89", x"8a", x"8a", x"89", x"89", x"89", x"8a", x"8c", x"8b", 
        x"8b", x"8c", x"8c", x"8b", x"89", x"8b", x"8a", x"8b", x"8a", x"88", x"89", x"89", x"8a", x"8c", x"8b", 
        x"8b", x"8a", x"8b", x"8c", x"8d", x"8e", x"8c", x"8c", x"8c", x"8c", x"8a", x"8a", x"8c", x"8c", x"8b", 
        x"8c", x"8c", x"8a", x"89", x"8a", x"8a", x"8b", x"8c", x"8d", x"8e", x"8e", x"8c", x"8b", x"8b", x"8c", 
        x"8d", x"8d", x"8e", x"8d", x"8c", x"8c", x"8d", x"8e", x"8d", x"8c", x"8e", x"8f", x"8e", x"8e", x"8d", 
        x"8e", x"8f", x"82", x"9a", x"7c", x"72", x"7b", x"7a", x"7c", x"7d", x"7a", x"79", x"7b", x"7d", x"7a", 
        x"79", x"7d", x"7a", x"92", x"8a", x"71", x"4d", x"30", x"2a", x"1d", x"0c", x"05", x"04", x"03", x"05", 
        x"08", x"11", x"2e", x"5f", x"81", x"88", x"84", x"69", x"3c", x"36", x"38", x"5f", x"7d", x"73", x"72", 
        x"59", x"77", x"d8", x"d5", x"d8", x"d8", x"ba", x"8d", x"7d", x"96", x"be", x"d3", x"d4", x"cf", x"cd", 
        x"cc", x"cd", x"cb", x"cf", x"d1", x"d0", x"d0", x"d0", x"d2", x"d1", x"cf", x"cf", x"cf", x"d0", x"d1", 
        x"d2", x"d2", x"d3", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", 
        x"d0", x"d2", x"d2", x"d3", x"d2", x"d2", x"d1", x"d2", x"d9", x"da", x"d1", x"d4", x"d2", x"d4", x"d4", 
        x"cf", x"e3", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ee", x"ef", x"ee", x"ee", 
        x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ee", x"ed", x"ed", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", x"ec", x"f0", x"ef", x"f0", 
        x"ee", x"f1", x"ee", x"ed", x"ef", x"eb", x"e3", x"d5", x"bd", x"a8", x"a6", x"ae", x"c1", x"d5", x"e4", 
        x"eb", x"f0", x"f2", x"f4", x"f4", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f0", x"f1", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f2", x"f4", x"f4", x"ef", x"ee", x"f2", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f3", x"f2", x"f3", x"f1", x"ea", x"e0", x"d0", x"c3", x"c8", x"d5", x"e2", x"ec", 
        x"f2", x"f5", x"f5", x"f5", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f3", x"f0", x"ef", x"f1", x"f3", x"f2", x"ef", 
        x"e7", x"d9", x"c9", x"c7", x"d3", x"e2", x"e9", x"ed", x"f1", x"ef", x"ef", x"f0", x"f2", x"f2", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f1", x"f2", 
        x"f0", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"f1", x"f0", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f0", x"f0", x"f1", x"ee", x"e7", x"e6", x"e2", 
        x"cc", x"b7", x"a9", x"85", x"5e", x"31", x"22", x"1d", x"1b", x"2a", x"47", x"6c", x"79", x"71", x"6a", 
        x"61", x"59", x"4d", x"45", x"40", x"3d", x"3b", x"37", x"37", x"36", x"33", x"31", x"31", x"2d", x"29", 
        x"2f", x"33", x"2c", x"26", x"3b", x"7f", x"9d", x"9c", x"9c", x"7a", x"52", x"52", x"4c", x"49", x"42", 
        x"2a", x"28", x"28", x"26", x"26", x"24", x"25", x"28", x"26", x"25", x"26", x"26", x"25", x"25", x"27", 
        x"27", x"27", x"24", x"23", x"22", x"23", x"22", x"1b", x"27", x"2a", x"15", x"1c", x"3c", x"3f", x"75", 
        x"82", x"59", x"45", x"33", x"28", x"25", x"29", x"39", x"5b", x"85", x"aa", x"c0", x"d3", x"d6", x"d7", 
        x"8c", x"8e", x"8d", x"8b", x"8b", x"8a", x"88", x"8b", x"8b", x"8a", x"8a", x"8a", x"8a", x"8c", x"8c", 
        x"8b", x"8b", x"8b", x"8a", x"8a", x"8a", x"89", x"89", x"8a", x"8a", x"89", x"88", x"89", x"8a", x"8a", 
        x"88", x"89", x"8c", x"8b", x"8a", x"8b", x"88", x"87", x"87", x"89", x"8a", x"8a", x"89", x"8c", x"8a", 
        x"8c", x"8a", x"88", x"8a", x"8a", x"8b", x"8b", x"8c", x"8c", x"8b", x"8b", x"89", x"8a", x"8b", x"8b", 
        x"8b", x"8b", x"8b", x"8b", x"8c", x"8c", x"8d", x"8d", x"8c", x"8b", x"8b", x"8b", x"8d", x"8d", x"8c", 
        x"8c", x"8c", x"8b", x"8b", x"8a", x"8a", x"8c", x"8e", x"8e", x"8e", x"8d", x"8c", x"8c", x"8c", x"8d", 
        x"8d", x"8d", x"8d", x"8f", x"8e", x"8d", x"8f", x"8e", x"8c", x"8d", x"8d", x"8d", x"8d", x"8e", x"8f", 
        x"8d", x"8e", x"82", x"9a", x"81", x"78", x"7d", x"7b", x"77", x"7a", x"7d", x"7d", x"7d", x"7c", x"7c", 
        x"7d", x"81", x"86", x"84", x"5e", x"26", x"28", x"22", x"0b", x"04", x"05", x"05", x"05", x"08", x"10", 
        x"2d", x"5a", x"84", x"89", x"80", x"7b", x"80", x"6e", x"3d", x"36", x"37", x"5f", x"7b", x"72", x"70", 
        x"5b", x"86", x"de", x"dd", x"c3", x"91", x"5e", x"93", x"cb", x"d9", x"d3", x"cc", x"ce", x"ce", x"cc", 
        x"cc", x"ce", x"ce", x"d0", x"d0", x"d0", x"d0", x"d1", x"d2", x"d0", x"d0", x"d1", x"d2", x"d2", x"d1", 
        x"d1", x"d2", x"d2", x"d0", x"d0", x"d0", x"d2", x"d3", x"d3", x"d3", x"d2", x"d1", x"d0", x"d0", x"d2", 
        x"d1", x"d1", x"d2", x"d1", x"d0", x"d1", x"d2", x"d2", x"d7", x"d9", x"d2", x"d5", x"d4", x"d6", x"d5", 
        x"d0", x"e1", x"f0", x"ee", x"ef", x"ed", x"ed", x"ef", x"f1", x"f0", x"ef", x"ed", x"ed", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f0", x"ef", x"ed", x"ee", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"e9", x"ee", x"f0", x"f1", 
        x"f0", x"f0", x"f1", x"f0", x"ee", x"ee", x"f1", x"f4", x"f6", x"f5", x"e8", x"cc", x"af", x"9c", x"9f", 
        x"b0", x"c8", x"d7", x"e5", x"ee", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f2", x"f3", x"f0", x"f0", x"f2", x"f2", x"f0", x"f0", x"f0", x"ef", x"ed", x"ed", x"ef", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f0", x"ee", x"ef", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f5", x"f4", x"e5", x"ce", x"c1", x"c5", 
        x"d4", x"e2", x"ec", x"f3", x"f4", x"f2", x"f2", x"f3", x"f3", x"f2", x"f3", x"f5", x"f5", x"f3", x"f1", 
        x"f2", x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f3", x"f2", x"e8", x"d4", x"c2", x"c4", x"d5", x"e6", x"ee", x"ef", x"f0", x"f1", x"f4", x"f0", 
        x"ee", x"f1", x"f2", x"f1", x"f2", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"f1", x"ef", x"ef", x"f0", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"ed", x"ed", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"ec", x"c9", x"99", x"85", 
        x"63", x"3b", x"18", x"07", x"06", x"16", x"3a", x"5d", x"7a", x"81", x"78", x"77", x"81", x"7c", x"65", 
        x"52", x"4d", x"4a", x"48", x"49", x"46", x"40", x"3b", x"38", x"39", x"36", x"33", x"32", x"33", x"31", 
        x"30", x"31", x"2e", x"28", x"34", x"7c", x"a2", x"9b", x"9f", x"80", x"55", x"57", x"50", x"4c", x"46", 
        x"2f", x"26", x"25", x"25", x"28", x"26", x"28", x"28", x"25", x"26", x"27", x"26", x"24", x"23", x"24", 
        x"26", x"23", x"21", x"23", x"24", x"26", x"2a", x"20", x"24", x"2f", x"1a", x"20", x"30", x"31", x"36", 
        x"2a", x"20", x"26", x"37", x"5b", x"87", x"ae", x"cc", x"df", x"e1", x"d7", x"d2", x"d2", x"d4", x"d5", 
        x"8c", x"8d", x"8c", x"8a", x"8b", x"8b", x"89", x"8b", x"8b", x"8a", x"89", x"8a", x"8b", x"8c", x"8b", 
        x"8b", x"8b", x"8b", x"8b", x"8b", x"8a", x"8a", x"89", x"8a", x"8a", x"89", x"89", x"8a", x"8b", x"8b", 
        x"89", x"8a", x"8b", x"89", x"89", x"8a", x"89", x"89", x"89", x"8a", x"89", x"89", x"8a", x"8d", x"8e", 
        x"8e", x"8c", x"8b", x"8c", x"8d", x"8c", x"8b", x"8d", x"8c", x"8b", x"8a", x"89", x"8a", x"8a", x"8a", 
        x"8a", x"8a", x"8a", x"8a", x"8b", x"8c", x"8c", x"8d", x"8c", x"8c", x"8c", x"8c", x"8d", x"8d", x"8c", 
        x"8b", x"8b", x"8c", x"8c", x"8c", x"8c", x"8d", x"8d", x"8d", x"8d", x"8c", x"8c", x"8c", x"8c", x"8d", 
        x"8d", x"8d", x"8d", x"8e", x"8d", x"8c", x"8e", x"8e", x"8d", x"8e", x"8f", x"8f", x"8e", x"8d", x"8e", 
        x"8d", x"8f", x"84", x"9b", x"7e", x"74", x"7c", x"7d", x"79", x"78", x"7b", x"7c", x"7b", x"7b", x"81", 
        x"83", x"7c", x"5d", x"3c", x"26", x"19", x"10", x"0a", x"10", x"08", x"04", x"06", x"12", x"2e", x"56", 
        x"7e", x"89", x"87", x"7e", x"7b", x"80", x"83", x"6c", x"3c", x"38", x"38", x"60", x"7e", x"72", x"78", 
        x"79", x"a1", x"c5", x"9f", x"81", x"97", x"bb", x"de", x"d6", x"cf", x"cd", x"cf", x"ce", x"cd", x"cf", 
        x"cd", x"ce", x"cd", x"d0", x"d0", x"d0", x"d0", x"cf", x"cf", x"d0", x"d1", x"d2", x"d1", x"d1", x"d2", 
        x"d3", x"d3", x"d2", x"d0", x"cf", x"cf", x"d1", x"d3", x"d3", x"d3", x"d2", x"d1", x"d0", x"d0", x"d2", 
        x"d1", x"d1", x"d2", x"d1", x"d0", x"d2", x"d0", x"d0", x"d6", x"d9", x"d1", x"d3", x"d1", x"d4", x"d4", 
        x"cf", x"e1", x"f0", x"ed", x"ef", x"ed", x"ee", x"ef", x"f0", x"f0", x"ef", x"ed", x"ed", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"e9", x"ee", x"f0", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"e8", x"d6", 
        x"c6", x"b3", x"ad", x"ad", x"b6", x"c6", x"d9", x"e5", x"f1", x"f4", x"f3", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f0", x"f1", x"f2", x"f2", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f0", x"ee", x"ef", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f1", x"eb", x"e1", 
        x"d6", x"cb", x"cc", x"d5", x"e0", x"ea", x"f0", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f4", x"f5", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f5", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"eb", x"dd", x"d2", x"ca", x"cd", x"d5", x"e1", x"ec", x"f0", x"f3", 
        x"f3", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"ed", x"ed", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ee", x"cf", x"9b", x"78", 
        x"6c", x"70", x"2d", x"14", x"1a", x"46", x"73", x"86", x"93", x"87", x"7b", x"73", x"6e", x"6f", x"73", 
        x"78", x"72", x"5a", x"47", x"48", x"48", x"3d", x"3d", x"40", x"38", x"34", x"34", x"33", x"33", x"35", 
        x"32", x"31", x"2d", x"27", x"2f", x"79", x"a1", x"9a", x"a0", x"86", x"5a", x"59", x"54", x"51", x"49", 
        x"2f", x"26", x"26", x"27", x"27", x"28", x"28", x"26", x"25", x"26", x"27", x"26", x"25", x"23", x"22", 
        x"23", x"25", x"28", x"2a", x"2a", x"2b", x"2e", x"23", x"21", x"2b", x"19", x"18", x"28", x"36", x"49", 
        x"60", x"80", x"a3", x"bf", x"cc", x"d4", x"d4", x"d6", x"d6", x"d4", x"d2", x"d4", x"d4", x"d4", x"d5", 
        x"8c", x"8d", x"8c", x"8a", x"8b", x"8c", x"8b", x"8b", x"8b", x"8b", x"8a", x"8a", x"8b", x"8b", x"8b", 
        x"8a", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8a", x"8b", x"8b", x"8a", x"8a", x"8b", x"8b", x"8b", 
        x"8a", x"8b", x"89", x"88", x"88", x"8a", x"8b", x"8c", x"8c", x"8b", x"8a", x"8a", x"8b", x"8b", x"8d", 
        x"8c", x"8b", x"8b", x"8a", x"8c", x"8b", x"8b", x"8e", x"8d", x"8b", x"8b", x"8a", x"8c", x"8c", x"8c", 
        x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8d", x"8d", x"8d", x"8d", x"8e", x"8e", x"8e", x"8e", x"8d", 
        x"8c", x"8c", x"8c", x"8d", x"8e", x"8e", x"8e", x"8e", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", 
        x"8d", x"8e", x"8e", x"8d", x"8c", x"8c", x"8e", x"8e", x"8e", x"8f", x"8f", x"8f", x"8e", x"8d", x"8d", 
        x"8d", x"8f", x"84", x"97", x"7d", x"73", x"7b", x"7b", x"7d", x"7b", x"77", x"79", x"81", x"89", x"82", 
        x"68", x"44", x"2b", x"20", x"12", x"08", x"05", x"11", x"35", x"17", x"04", x"10", x"45", x"75", x"8b", 
        x"8b", x"85", x"80", x"7e", x"80", x"80", x"7f", x"6c", x"3e", x"37", x"37", x"5c", x"80", x"7e", x"88", 
        x"87", x"86", x"8f", x"92", x"bf", x"df", x"db", x"e0", x"d7", x"cb", x"cb", x"cf", x"ce", x"ce", x"cf", 
        x"cd", x"ce", x"cd", x"cf", x"d0", x"d0", x"d0", x"cf", x"d1", x"d3", x"d2", x"d1", x"d0", x"d0", x"d0", 
        x"d2", x"d2", x"d2", x"d0", x"cf", x"d0", x"d1", x"d3", x"d3", x"d3", x"d2", x"d2", x"d1", x"d1", x"d3", 
        x"d2", x"d2", x"d3", x"d2", x"d1", x"d2", x"d0", x"d0", x"d6", x"d9", x"d1", x"d3", x"d1", x"d3", x"d3", 
        x"cf", x"e0", x"ef", x"ed", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"ef", x"f0", x"ef", x"ee", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"ef", x"e9", x"ee", x"f0", x"f1", 
        x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f2", x"f2", x"f2", x"f4", x"f5", 
        x"f5", x"f0", x"e0", x"c7", x"b4", x"ab", x"af", x"b7", x"c3", x"d0", x"de", x"ec", x"f3", x"f3", x"f1", 
        x"f0", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f0", x"ee", x"f1", x"f5", 
        x"f3", x"ec", x"df", x"d4", x"d0", x"d2", x"d8", x"e1", x"e9", x"f0", x"f3", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f5", x"f6", x"f6", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f2", x"f0", x"ef", x"f1", x"f3", x"f3", x"f2", x"e6", x"d2", x"c3", x"c6", x"d2", x"de", x"eb", 
        x"f4", x"f4", x"f3", x"f3", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"ed", x"ed", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ed", x"f4", x"f5", x"e1", x"b2", 
        x"8b", x"82", x"44", x"26", x"2d", x"61", x"7f", x"80", x"8c", x"87", x"8a", x"89", x"7c", x"71", x"6f", 
        x"70", x"76", x"77", x"60", x"4c", x"43", x"3e", x"3d", x"3d", x"36", x"35", x"37", x"34", x"32", x"32", 
        x"2f", x"30", x"2d", x"27", x"29", x"75", x"a0", x"9c", x"a0", x"8b", x"5f", x"5c", x"56", x"54", x"4c", 
        x"33", x"25", x"24", x"29", x"29", x"25", x"26", x"25", x"23", x"24", x"25", x"26", x"28", x"27", x"25", 
        x"27", x"29", x"29", x"27", x"29", x"2d", x"26", x"19", x"24", x"3d", x"42", x"53", x"76", x"98", x"bb", 
        x"d0", x"d9", x"db", x"db", x"d6", x"d2", x"d6", x"d6", x"d4", x"d4", x"d6", x"d6", x"d3", x"d5", x"d6", 
        x"8c", x"8d", x"8c", x"8a", x"8b", x"8d", x"8b", x"8b", x"8b", x"8b", x"8c", x"8b", x"8b", x"8b", x"8a", 
        x"8a", x"8b", x"8b", x"8c", x"8c", x"8c", x"8b", x"8b", x"8c", x"8c", x"8b", x"8a", x"8b", x"8b", x"89", 
        x"8a", x"8a", x"89", x"89", x"8a", x"8b", x"8b", x"8c", x"8d", x"8b", x"8a", x"8a", x"8b", x"8b", x"8e", 
        x"8c", x"8b", x"8d", x"8a", x"8c", x"8b", x"8b", x"8f", x"8d", x"8b", x"8b", x"8b", x"8c", x"8b", x"8b", 
        x"8b", x"8b", x"8b", x"8b", x"8c", x"8c", x"8c", x"8c", x"8d", x"8d", x"8e", x"8d", x"8d", x"8d", x"8c", 
        x"8c", x"8c", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8e", x"8e", x"8e", x"8e", x"8e", 
        x"8e", x"8e", x"8f", x"8f", x"8f", x"8f", x"8f", x"8f", x"8f", x"8f", x"8e", x"8e", x"8f", x"8f", x"8e", 
        x"8f", x"90", x"83", x"91", x"78", x"6f", x"7b", x"7e", x"81", x"80", x"81", x"8a", x"83", x"66", x"46", 
        x"30", x"1d", x"14", x"0c", x"03", x"03", x"04", x"1e", x"58", x"28", x"05", x"2b", x"81", x"8d", x"80", 
        x"81", x"80", x"7e", x"7f", x"7e", x"80", x"83", x"6a", x"36", x"3d", x"5c", x"78", x"8f", x"8d", x"7d", 
        x"5a", x"6c", x"be", x"dc", x"dd", x"d7", x"d9", x"dd", x"d9", x"ce", x"cf", x"cd", x"cd", x"d0", x"cc", 
        x"cd", x"d0", x"cf", x"d1", x"d1", x"d0", x"d0", x"d1", x"d4", x"d4", x"d3", x"d1", x"cf", x"d0", x"d0", 
        x"d0", x"d0", x"d1", x"d0", x"d1", x"d1", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", x"d1", x"d1", x"d3", 
        x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d7", x"d9", x"d1", x"d4", x"d3", x"d4", x"d3", 
        x"cf", x"e0", x"ef", x"ed", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", 
        x"ef", x"ef", x"f0", x"ee", x"ec", x"ef", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"e9", x"ee", x"f0", x"f1", 
        x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"ed", x"dd", x"ce", x"be", x"b1", x"a6", x"a5", x"b4", x"ce", x"e5", 
        x"f4", x"f6", x"f5", x"f3", x"ef", x"ef", x"f1", x"f2", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"ef", x"f0", x"ef", x"ed", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f2", x"f5", x"f4", x"ed", x"e6", x"dd", x"d5", x"d3", x"d6", x"dd", x"e7", x"f1", x"f5", x"f4", 
        x"f1", x"f0", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f3", x"f4", x"f5", x"f4", x"f3", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"ef", x"f1", x"f2", x"f4", x"f1", x"e5", x"d2", x"c6", x"c4", 
        x"cb", x"dc", x"ed", x"f6", x"f4", x"f2", x"f0", x"f0", x"f2", x"f3", x"f2", x"f0", x"ef", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"ee", x"ed", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f1", x"e6", x"bc", 
        x"9d", x"9b", x"5c", x"25", x"29", x"68", x"83", x"82", x"98", x"89", x"87", x"8b", x"85", x"82", x"82", 
        x"7d", x"6f", x"69", x"6f", x"65", x"4d", x"3e", x"3f", x"3d", x"37", x"38", x"36", x"36", x"36", x"34", 
        x"32", x"32", x"2f", x"2a", x"26", x"71", x"a1", x"9e", x"a2", x"8f", x"64", x"61", x"59", x"53", x"4d", 
        x"31", x"2d", x"2a", x"22", x"24", x"27", x"26", x"25", x"28", x"2b", x"2a", x"27", x"26", x"29", x"2c", 
        x"2c", x"2c", x"26", x"17", x"16", x"2b", x"46", x"62", x"7f", x"a3", x"b8", x"c9", x"d3", x"da", x"da", 
        x"d8", x"d3", x"d0", x"d3", x"d6", x"d4", x"d7", x"d7", x"d6", x"d6", x"d5", x"d4", x"d3", x"d5", x"d7", 
        x"8d", x"8e", x"8d", x"8a", x"8c", x"8d", x"8b", x"8b", x"8c", x"8c", x"8d", x"8c", x"8c", x"8b", x"8a", 
        x"8b", x"8b", x"8b", x"8c", x"8c", x"8c", x"8b", x"8b", x"8c", x"8c", x"8b", x"8a", x"8b", x"8a", x"89", 
        x"8b", x"8a", x"8a", x"8b", x"8c", x"8c", x"8c", x"8d", x"8d", x"8c", x"8b", x"8b", x"8b", x"8a", x"8d", 
        x"8c", x"8b", x"8c", x"8b", x"8d", x"8c", x"8b", x"8e", x"8d", x"8c", x"8b", x"8c", x"8e", x"8d", x"8d", 
        x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8e", x"8d", x"8c", x"8d", x"8d", 
        x"8d", x"8e", x"8e", x"8e", x"8d", x"8d", x"8e", x"8e", x"8f", x"8f", x"8f", x"8e", x"8e", x"8e", x"8e", 
        x"8e", x"8f", x"8f", x"8f", x"90", x"91", x"8f", x"8f", x"90", x"8f", x"8e", x"8d", x"91", x"90", x"8f", 
        x"90", x"90", x"84", x"93", x"7e", x"74", x"7c", x"7e", x"82", x"82", x"83", x"6c", x"4c", x"31", x"22", 
        x"15", x"0a", x"05", x"06", x"07", x"15", x"35", x"50", x"5d", x"3e", x"35", x"66", x"9e", x"84", x"7f", 
        x"83", x"82", x"82", x"7e", x"7a", x"80", x"84", x"70", x"55", x"79", x"89", x"8e", x"80", x"5f", x"43", 
        x"30", x"77", x"de", x"dd", x"db", x"d9", x"d5", x"df", x"db", x"cd", x"d0", x"cf", x"cf", x"d1", x"ce", 
        x"ce", x"d1", x"d0", x"d1", x"d0", x"d0", x"d0", x"d1", x"d3", x"d3", x"d2", x"d1", x"d1", x"d2", x"d3", 
        x"d1", x"d1", x"d2", x"d0", x"d0", x"d0", x"d3", x"d3", x"d3", x"d4", x"d3", x"d3", x"d2", x"d2", x"d2", 
        x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d7", x"d9", x"d2", x"d5", x"d4", x"d4", x"d3", 
        x"cf", x"e0", x"ef", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", 
        x"ef", x"ef", x"ef", x"ed", x"eb", x"ef", x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", x"ee", x"ef", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"e9", x"ee", x"f0", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"ee", x"f0", x"f3", x"f2", x"f2", x"ef", x"e4", x"d4", x"c6", x"bb", x"b3", x"ad", 
        x"b4", x"c3", x"d6", x"e8", x"ef", x"f0", x"f1", x"f2", x"f1", x"ee", x"ee", x"f0", x"f1", x"f0", x"ef", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"ef", x"f0", x"ef", x"ec", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f1", x"ef", x"f0", x"f1", x"f2", x"f4", x"f4", x"ee", x"e8", x"e2", x"db", x"d9", x"dc", x"e3", x"ec", 
        x"f1", x"f1", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f3", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"e8", x"db", 
        x"ce", x"c8", x"c8", x"d6", x"e8", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"f1", x"ef", x"ef", x"f0", 
        x"f2", x"ee", x"ed", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"ee", x"f1", x"ef", x"d8", 
        x"c3", x"b4", x"6e", x"2b", x"37", x"74", x"86", x"82", x"a3", x"91", x"87", x"87", x"84", x"85", x"88", 
        x"8a", x"85", x"79", x"6f", x"77", x"77", x"50", x"36", x"34", x"38", x"38", x"37", x"3a", x"39", x"34", 
        x"32", x"33", x"31", x"2b", x"26", x"6e", x"a3", x"a0", x"a3", x"93", x"6a", x"69", x"5f", x"56", x"52", 
        x"3a", x"3b", x"36", x"24", x"23", x"2a", x"2a", x"2a", x"29", x"28", x"2b", x"2c", x"2a", x"29", x"26", 
        x"22", x"2a", x"40", x"5d", x"78", x"95", x"ae", x"c3", x"cd", x"d4", x"d8", x"d7", x"d5", x"d7", x"d6", 
        x"d5", x"d7", x"d7", x"d6", x"d6", x"d5", x"d5", x"d5", x"d6", x"d7", x"d6", x"d4", x"d4", x"d5", x"d6", 
        x"8d", x"8f", x"8e", x"8b", x"8c", x"8c", x"8a", x"8b", x"8b", x"8c", x"8d", x"8d", x"8c", x"8b", x"8c", 
        x"8c", x"8c", x"8c", x"8c", x"8c", x"8b", x"8b", x"8a", x"8c", x"8b", x"8a", x"8a", x"8b", x"8b", x"8a", 
        x"8b", x"8a", x"8a", x"8c", x"8c", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8b", x"8a", x"8a", 
        x"8b", x"8a", x"8a", x"8b", x"8d", x"8c", x"8b", x"8e", x"8d", x"8d", x"8d", x"8d", x"8d", x"8c", x"8c", 
        x"8c", x"8c", x"8c", x"8c", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8c", x"8b", x"8c", x"8e", 
        x"8e", x"8e", x"8e", x"8d", x"8d", x"8e", x"8e", x"8f", x"8f", x"8e", x"8d", x"8d", x"8d", x"8d", x"8e", 
        x"8e", x"8e", x"8f", x"8e", x"8f", x"90", x"8d", x"8d", x"8f", x"8e", x"8e", x"8e", x"91", x"90", x"8e", 
        x"90", x"91", x"83", x"8c", x"7c", x"75", x"7e", x"84", x"84", x"7b", x"4f", x"37", x"25", x"17", x"0d", 
        x"07", x"03", x"03", x"0c", x"29", x"4e", x"67", x"6a", x"60", x"65", x"5f", x"84", x"ad", x"85", x"82", 
        x"85", x"86", x"80", x"78", x"7a", x"7f", x"80", x"86", x"86", x"95", x"85", x"66", x"44", x"35", x"36", 
        x"39", x"85", x"d9", x"de", x"df", x"db", x"d1", x"e0", x"db", x"cc", x"d0", x"d0", x"d0", x"cf", x"cf", 
        x"d0", x"d2", x"d1", x"d2", x"d1", x"d0", x"d1", x"d0", x"d0", x"d0", x"d1", x"d2", x"d2", x"d3", x"d2", 
        x"d2", x"d2", x"d2", x"d0", x"d0", x"d0", x"d2", x"d3", x"d3", x"d4", x"d3", x"d3", x"d3", x"d2", x"d3", 
        x"d4", x"d3", x"d2", x"d2", x"d3", x"d2", x"d2", x"d2", x"d7", x"d9", x"d1", x"d5", x"d4", x"d5", x"d4", 
        x"cf", x"e1", x"f0", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ef", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"e9", x"ee", x"f0", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"ef", x"ee", x"f0", x"f2", x"f2", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f1", x"f2", x"f1", x"f2", x"f3", x"f4", x"f0", x"e3", x"d5", 
        x"c6", x"b6", x"a8", x"a8", x"b7", x"ce", x"e5", x"f1", x"f3", x"f1", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"ef", x"f0", x"ef", x"eb", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f0", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"ef", x"ec", x"e6", x"df", x"db", 
        x"dd", x"e3", x"ee", x"f1", x"f3", x"f4", x"f4", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f5", 
        x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f3", x"f1", x"f1", x"f4", x"f3", x"f2", 
        x"f0", x"e6", x"d8", x"c9", x"c4", x"ca", x"dc", x"ee", x"f5", x"f2", x"ed", x"ee", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"ef", x"ef", x"ef", 
        x"f2", x"ef", x"ed", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f3", x"ed", 
        x"ee", x"e7", x"96", x"3e", x"40", x"73", x"8c", x"85", x"a2", x"97", x"8d", x"89", x"87", x"87", x"86", 
        x"84", x"82", x"83", x"82", x"77", x"76", x"83", x"6b", x"45", x"33", x"30", x"37", x"3a", x"38", x"35", 
        x"31", x"34", x"31", x"2c", x"27", x"69", x"a3", x"a0", x"a0", x"94", x"6e", x"6c", x"64", x"5c", x"58", 
        x"3d", x"2b", x"28", x"29", x"28", x"29", x"2c", x"2b", x"2c", x"2e", x"2b", x"1f", x"1d", x"2e", x"4b", 
        x"72", x"92", x"ae", x"c1", x"ce", x"d5", x"d8", x"d8", x"d5", x"d2", x"d6", x"d3", x"d4", x"d6", x"d5", 
        x"d5", x"d8", x"d6", x"d4", x"d7", x"d8", x"d9", x"d6", x"d6", x"d6", x"d4", x"d2", x"d3", x"d4", x"d5", 
        x"8d", x"8f", x"8e", x"8c", x"8c", x"8c", x"89", x"8a", x"8b", x"8d", x"8d", x"8d", x"8c", x"8b", x"8c", 
        x"8d", x"8c", x"8c", x"8c", x"8c", x"8b", x"8b", x"8a", x"8c", x"8b", x"8a", x"8a", x"8b", x"8c", x"8c", 
        x"8c", x"8b", x"8a", x"8c", x"8d", x"8a", x"8a", x"8a", x"89", x"8b", x"8c", x"8c", x"8b", x"8d", x"8c", 
        x"8f", x"8e", x"8c", x"8f", x"90", x"8d", x"8b", x"8d", x"8d", x"8d", x"8e", x"8d", x"8d", x"8d", x"8d", 
        x"8d", x"8d", x"8d", x"8d", x"8e", x"8f", x"8e", x"8e", x"8d", x"8d", x"8d", x"8c", x"8b", x"8c", x"8e", 
        x"8f", x"8f", x"8e", x"8d", x"8f", x"90", x"90", x"90", x"8f", x"8d", x"8c", x"8c", x"8d", x"8d", x"8e", 
        x"8e", x"8e", x"8e", x"8c", x"8c", x"8e", x"8c", x"8c", x"8f", x"8e", x"8e", x"8e", x"91", x"8f", x"8c", 
        x"90", x"91", x"7f", x"7d", x"73", x"79", x"85", x"7c", x"58", x"39", x"27", x"18", x"0a", x"05", x"03", 
        x"04", x"0b", x"26", x"54", x"69", x"68", x"78", x"73", x"7a", x"8c", x"65", x"81", x"aa", x"7f", x"82", 
        x"84", x"82", x"76", x"78", x"8f", x"96", x"87", x"8c", x"86", x"67", x"48", x"37", x"38", x"44", x"5b", 
        x"67", x"8e", x"dc", x"da", x"d8", x"dc", x"d9", x"e2", x"da", x"cf", x"d1", x"ce", x"cf", x"cd", x"ce", 
        x"d0", x"d2", x"d1", x"d2", x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"d0", x"d2", x"d1", x"d0", x"cf", 
        x"d0", x"d0", x"d1", x"d0", x"d1", x"d2", x"d4", x"d2", x"d3", x"d4", x"d3", x"d3", x"d2", x"d2", x"d3", 
        x"d4", x"d3", x"d2", x"d2", x"d3", x"d2", x"d0", x"d0", x"d6", x"d9", x"d1", x"d3", x"d2", x"d5", x"d5", 
        x"d0", x"e1", x"f0", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f2", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"ea", x"ee", x"f0", x"f1", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"f3", x"f2", x"ef", x"ef", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f2", x"f4", x"f4", x"f2", x"ee", x"ee", x"f1", x"f2", x"f1", 
        x"ef", x"eb", x"e3", x"d5", x"c1", x"b0", x"a8", x"b0", x"c2", x"d7", x"e9", x"ef", x"f0", x"f0", x"f2", 
        x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", x"f1", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"ef", x"f0", x"ef", x"ea", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"ee", 
        x"e5", x"dd", x"d7", x"dc", x"e4", x"eb", x"f0", x"f3", x"f4", x"f4", x"f3", x"f2", x"f1", x"f2", x"f3", 
        x"f4", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f1", x"f1", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f3", x"f4", x"f3", x"f3", x"f3", x"f0", x"f1", x"f2", 
        x"f0", x"f0", x"f1", x"ed", x"e4", x"d3", x"c6", x"c3", x"ce", x"e3", x"ef", x"f1", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"ef", x"ef", x"ef", 
        x"f2", x"ef", x"ed", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f1", x"ef", 
        x"ef", x"dd", x"8a", x"39", x"3e", x"6b", x"8b", x"85", x"a6", x"9d", x"93", x"8d", x"89", x"87", x"85", 
        x"82", x"81", x"80", x"82", x"82", x"79", x"76", x"82", x"86", x"6c", x"52", x"46", x"36", x"2f", x"35", 
        x"33", x"34", x"31", x"2b", x"29", x"65", x"a1", x"9f", x"9d", x"97", x"71", x"6a", x"65", x"5f", x"5c", 
        x"46", x"22", x"2a", x"49", x"47", x"35", x"2e", x"27", x"21", x"2a", x"44", x"6c", x"8e", x"ac", x"c2", 
        x"d1", x"d9", x"d7", x"d7", x"d8", x"d5", x"d3", x"d7", x"d8", x"d6", x"d9", x"d5", x"d5", x"d6", x"d8", 
        x"d6", x"d7", x"d5", x"d7", x"da", x"d4", x"d3", x"d3", x"d6", x"d8", x"d5", x"d3", x"d5", x"d5", x"d5", 
        x"8c", x"8d", x"8e", x"8e", x"8d", x"8c", x"8b", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8a", 
        x"8a", x"8c", x"8d", x"8e", x"8d", x"8c", x"8c", x"8b", x"8c", x"8c", x"8c", x"8c", x"8b", x"8c", x"8c", 
        x"8b", x"8b", x"8c", x"8c", x"8d", x"8e", x"8c", x"8c", x"8d", x"8d", x"8c", x"8c", x"8b", x"8e", x"8c", 
        x"8e", x"8e", x"8b", x"8f", x"8e", x"8b", x"8c", x"8c", x"8d", x"8c", x"8c", x"8e", x"8c", x"8c", x"8d", 
        x"8b", x"8c", x"8f", x"8f", x"8e", x"8e", x"8d", x"8f", x"8f", x"8d", x"8b", x"8c", x"8d", x"8d", x"8d", 
        x"8d", x"8d", x"8d", x"8d", x"8f", x"90", x"90", x"90", x"90", x"90", x"8f", x"90", x"8e", x"8d", x"8e", 
        x"90", x"90", x"8e", x"90", x"90", x"90", x"8f", x"90", x"91", x"90", x"8f", x"8e", x"8c", x"8e", x"8d", 
        x"90", x"8e", x"80", x"89", x"86", x"79", x"5d", x"3e", x"28", x"1d", x"0e", x"08", x"03", x"05", x"0b", 
        x"1e", x"40", x"63", x"7b", x"7a", x"79", x"85", x"77", x"8a", x"8d", x"53", x"7e", x"a9", x"83", x"83", 
        x"7c", x"79", x"89", x"b9", x"cf", x"a4", x"84", x"68", x"45", x"33", x"34", x"44", x"5c", x"72", x"7c", 
        x"77", x"90", x"db", x"da", x"d7", x"db", x"da", x"e2", x"da", x"d0", x"d1", x"d1", x"cf", x"cf", x"d0", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"cf", x"cf", x"d1", x"d2", x"d2", x"d2", x"d1", x"d1", 
        x"d2", x"d1", x"d0", x"d0", x"d1", x"d3", x"d4", x"d3", x"d4", x"d5", x"d2", x"d1", x"d2", x"d3", x"d2", 
        x"d3", x"d2", x"d2", x"d2", x"d1", x"d1", x"d2", x"d1", x"d6", x"da", x"cf", x"d3", x"d1", x"d4", x"d4", 
        x"d1", x"de", x"f1", x"ed", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ed", x"ec", x"ed", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"eb", x"ee", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"eb", x"e0", x"d0", x"bb", x"ab", x"ad", x"b9", x"cc", x"e0", x"ea", 
        x"ef", x"f2", x"f3", x"f1", x"ed", x"ee", x"f0", x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", x"f2", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"eb", x"f1", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"ed", x"e6", x"da", x"d4", x"d8", x"e3", x"ec", x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f3", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f4", 
        x"f4", x"f1", x"ee", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f3", x"f3", x"f1", x"f2", x"f2", 
        x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"eb", x"dd", x"cb", x"bf", x"c7", x"d9", x"e9", x"ef", x"f1", 
        x"f0", x"ef", x"f0", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"ef", x"f0", 
        x"f0", x"ef", x"ef", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f0", 
        x"f2", x"d9", x"8e", x"43", x"38", x"67", x"8e", x"86", x"a8", x"a1", x"93", x"8d", x"8b", x"8a", x"89", 
        x"83", x"84", x"84", x"81", x"82", x"83", x"7b", x"73", x"77", x"89", x"80", x"6a", x"55", x"43", x"35", 
        x"32", x"36", x"36", x"2d", x"2c", x"5d", x"9e", x"a4", x"a9", x"af", x"88", x"6c", x"6d", x"65", x"67", 
        x"52", x"2e", x"2a", x"34", x"33", x"2d", x"3f", x"61", x"86", x"a6", x"bf", x"d1", x"d4", x"d4", x"d7", 
        x"d9", x"d8", x"d7", x"d6", x"d7", x"d5", x"d5", x"d6", x"d6", x"d6", x"d8", x"d8", x"d7", x"d5", x"d7", 
        x"d6", x"d5", x"d5", x"d5", x"d6", x"d4", x"d4", x"d5", x"d5", x"d6", x"d6", x"d6", x"d6", x"d6", x"d5", 
        x"8e", x"8e", x"8d", x"8c", x"8c", x"8b", x"8b", x"8d", x"8c", x"8c", x"8c", x"8c", x"8c", x"8d", x"8b", 
        x"8b", x"8c", x"8d", x"8d", x"8d", x"8d", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8d", x"8f", 
        x"8c", x"8b", x"8b", x"8a", x"8b", x"8d", x"8e", x"8e", x"8d", x"8d", x"8c", x"8b", x"8b", x"8d", x"8c", 
        x"8e", x"8d", x"8b", x"8e", x"8d", x"8b", x"8d", x"8b", x"8c", x"8c", x"8d", x"8e", x"8c", x"8d", x"8e", 
        x"8d", x"8d", x"8e", x"8d", x"8c", x"8e", x"8e", x"8f", x"8f", x"8d", x"8c", x"8c", x"8e", x"8d", x"8c", 
        x"8c", x"8c", x"8e", x"8e", x"8f", x"90", x"90", x"90", x"90", x"91", x"91", x"90", x"8f", x"8e", x"8f", 
        x"90", x"90", x"8f", x"90", x"91", x"91", x"91", x"90", x"90", x"90", x"8f", x"8e", x"8d", x"8f", x"8e", 
        x"91", x"91", x"89", x"89", x"69", x"42", x"2d", x"21", x"0e", x"07", x"06", x"07", x"0d", x"1c", x"39", 
        x"58", x"6c", x"73", x"85", x"83", x"7a", x"80", x"76", x"8d", x"8b", x"51", x"7c", x"a5", x"7f", x"79", 
        x"8f", x"b2", x"cf", x"db", x"c6", x"84", x"4c", x"36", x"39", x"48", x"59", x"6c", x"7a", x"83", x"83", 
        x"78", x"91", x"dc", x"db", x"d8", x"da", x"d8", x"e1", x"da", x"d0", x"d1", x"d1", x"d0", x"cf", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", x"d2", x"d2", x"d3", x"d2", x"d1", x"d1", 
        x"d3", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d4", x"d3", x"d2", x"d2", x"d2", x"d1", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", x"d1", x"d0", x"d6", x"db", x"d0", x"d3", x"d0", x"d2", x"d3", 
        x"d0", x"de", x"f2", x"ed", x"f0", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ed", x"ed", x"ed", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f1", x"f0", 
        x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ea", x"ed", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f1", x"f2", x"f1", x"f1", x"f3", x"f2", x"ef", x"ec", x"e5", x"d8", x"c5", x"b8", x"b4", x"b7", 
        x"c7", x"d3", x"e0", x"ea", x"f0", x"f2", x"f3", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", 
        x"f4", x"f5", x"f3", x"f0", x"ef", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"eb", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f3", x"f0", x"ea", x"e4", x"dd", x"d7", x"da", x"e2", x"ea", x"f0", x"f2", x"f4", 
        x"f5", x"f1", x"f2", x"f4", x"f4", x"f2", x"f2", x"f4", x"f4", x"f3", x"f4", x"f4", x"f3", x"f2", x"f0", 
        x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f1", x"ed", x"f4", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"ef", x"e5", x"d6", x"c7", x"c5", x"d2", x"e1", 
        x"eb", x"ee", x"ef", x"f2", x"f3", x"f1", x"f0", x"ee", x"f0", x"f2", x"f2", x"ef", x"ef", x"ef", x"f1", 
        x"f1", x"ee", x"ed", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ed", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", 
        x"f2", x"da", x"84", x"42", x"39", x"67", x"90", x"85", x"ad", x"a5", x"95", x"90", x"8e", x"8c", x"8b", 
        x"86", x"84", x"83", x"83", x"82", x"82", x"80", x"7a", x"73", x"75", x"81", x"84", x"7a", x"67", x"53", 
        x"43", x"37", x"31", x"30", x"2a", x"5e", x"b7", x"c2", x"c1", x"c6", x"aa", x"7a", x"68", x"55", x"49", 
        x"36", x"2b", x"38", x"54", x"79", x"9e", x"b9", x"ca", x"d5", x"d8", x"d6", x"d8", x"d8", x"d7", x"d7", 
        x"d7", x"d7", x"d7", x"d7", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", x"d8", x"d8", x"d7", x"d5", x"d6", 
        x"d6", x"d5", x"d5", x"d5", x"d5", x"d4", x"d5", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", 
        x"8b", x"8c", x"8d", x"8e", x"8d", x"8d", x"8d", x"8d", x"8d", x"8c", x"8c", x"8c", x"8c", x"8d", x"8d", 
        x"8d", x"8d", x"8c", x"8c", x"8c", x"8d", x"8d", x"8d", x"8d", x"8c", x"8c", x"8c", x"8d", x"8d", x"8e", 
        x"8e", x"8c", x"8b", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8c", x"8d", x"8e", x"8e", x"8d", x"8c", 
        x"8d", x"8c", x"8c", x"8d", x"8d", x"8c", x"8d", x"8b", x"8d", x"8e", x"8e", x"8e", x"8d", x"8e", x"8f", 
        x"8f", x"8e", x"8d", x"8b", x"8a", x"8d", x"8f", x"90", x"8f", x"8f", x"8d", x"8c", x"8f", x"8e", x"8c", 
        x"8c", x"8c", x"8e", x"8f", x"90", x"90", x"90", x"90", x"90", x"91", x"91", x"90", x"8f", x"8f", x"90", 
        x"90", x"90", x"8f", x"90", x"91", x"91", x"91", x"90", x"90", x"90", x"8f", x"8e", x"8e", x"8f", x"8f", 
        x"91", x"95", x"7e", x"48", x"2c", x"21", x"15", x"08", x"04", x"04", x"05", x"0b", x"31", x"57", x"6a", 
        x"76", x"78", x"82", x"8b", x"83", x"7d", x"81", x"72", x"88", x"86", x"4f", x"78", x"9f", x"8e", x"af", 
        x"d3", x"dc", x"cf", x"9b", x"5e", x"3a", x"38", x"45", x"5b", x"70", x"7a", x"83", x"84", x"85", x"86", 
        x"7c", x"92", x"dd", x"dc", x"d8", x"da", x"d8", x"e0", x"d9", x"d0", x"d1", x"d1", x"d0", x"cf", x"d1", 
        x"d1", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", x"d2", x"d3", x"d2", x"d1", x"d0", x"d1", 
        x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d4", x"d3", x"d2", x"d1", x"d1", x"d2", x"d1", x"d0", x"d1", 
        x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"cf", x"d6", x"db", x"d0", x"d3", x"d0", x"d2", x"d3", 
        x"d0", x"de", x"f2", x"ee", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f1", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ea", x"ed", x"f0", x"f1", 
        x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f2", x"f3", x"f0", x"ef", x"f1", x"f3", x"f2", x"f1", x"f4", x"f5", x"f1", x"ee", x"e7", x"d5", 
        x"bd", x"b1", x"ae", x"b7", x"c9", x"da", x"e3", x"ea", x"ee", x"f1", x"f1", x"ef", x"ef", x"f1", x"f1", 
        x"f0", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"eb", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f3", x"f0", x"ef", x"f2", x"f2", x"f3", x"f4", x"f3", x"ee", x"e6", x"dc", x"d3", x"d3", x"de", x"e8", 
        x"ed", x"f3", x"f5", x"f5", x"f4", x"f3", x"f1", x"f1", x"ef", x"f0", x"f2", x"f3", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f1", x"f3", x"f3", x"f3", x"f2", x"f1", x"f3", 
        x"f3", x"f1", x"ed", x"f4", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f0", x"ed", x"ed", x"f0", x"f1", x"ee", x"e3", x"d2", x"c7", 
        x"c7", x"d6", x"e6", x"ed", x"ed", x"f0", x"f4", x"f2", x"ee", x"ee", x"f1", x"f1", x"f1", x"ef", x"ef", 
        x"f0", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ed", x"ee", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"db", x"89", x"49", x"39", x"60", x"8e", x"85", x"ac", x"a8", x"97", x"94", x"92", x"8f", x"8d", 
        x"8a", x"86", x"85", x"84", x"81", x"80", x"7f", x"7c", x"7b", x"7d", x"74", x"71", x"83", x"88", x"78", 
        x"67", x"53", x"41", x"31", x"29", x"64", x"c0", x"bf", x"ad", x"9b", x"7f", x"4c", x"34", x"34", x"46", 
        x"6c", x"93", x"b6", x"cc", x"d8", x"dc", x"d8", x"d7", x"db", x"da", x"d8", x"dc", x"dc", x"d8", x"d6", 
        x"d7", x"d7", x"d7", x"d7", x"d7", x"d7", x"d6", x"d6", x"d6", x"d6", x"d7", x"d7", x"d6", x"d6", x"d6", 
        x"d6", x"d6", x"d6", x"d5", x"d5", x"d4", x"d6", x"d7", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", 
        x"8b", x"8d", x"8e", x"90", x"8f", x"8d", x"8b", x"8c", x"8c", x"8d", x"8d", x"8d", x"8d", x"8c", x"8e", 
        x"8e", x"8d", x"8c", x"8b", x"8c", x"8c", x"8d", x"8e", x"8d", x"8c", x"8c", x"8d", x"8e", x"8c", x"89", 
        x"8c", x"8d", x"8d", x"8e", x"8d", x"8b", x"8d", x"8d", x"8c", x"8c", x"8d", x"8e", x"8f", x"8d", x"8c", 
        x"8c", x"8c", x"8c", x"8d", x"8d", x"8c", x"8d", x"8b", x"8e", x"8f", x"8f", x"8e", x"8d", x"8e", x"8e", 
        x"8e", x"8e", x"8d", x"8b", x"8b", x"8d", x"90", x"8f", x"8f", x"90", x"8e", x"8c", x"8f", x"8e", x"8e", 
        x"8d", x"8e", x"8e", x"8f", x"90", x"90", x"90", x"90", x"90", x"91", x"91", x"90", x"90", x"90", x"90", 
        x"90", x"90", x"90", x"90", x"91", x"92", x"91", x"8f", x"8f", x"90", x"90", x"8f", x"8d", x"8e", x"92", 
        x"93", x"94", x"79", x"30", x"17", x"0f", x"06", x"01", x"05", x"06", x"08", x"12", x"35", x"55", x"65", 
        x"76", x"81", x"82", x"8a", x"89", x"84", x"87", x"77", x"80", x"78", x"4d", x"80", x"c4", x"d1", x"dd", 
        x"c8", x"a0", x"66", x"39", x"35", x"46", x"59", x"6f", x"80", x"82", x"86", x"89", x"89", x"89", x"86", 
        x"7a", x"90", x"dd", x"dd", x"d9", x"db", x"d9", x"e1", x"da", x"d0", x"d1", x"d1", x"d0", x"cf", x"d1", 
        x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d2", x"d2", x"d2", x"d2", x"d0", x"d0", x"d1", 
        x"d2", x"d1", x"cf", x"cf", x"d1", x"d2", x"d3", x"d2", x"d1", x"d0", x"d1", x"d1", x"d0", x"cf", x"d1", 
        x"d1", x"d0", x"d0", x"d0", x"d1", x"d2", x"d1", x"cf", x"d5", x"da", x"cf", x"d3", x"d1", x"d3", x"d4", 
        x"d2", x"df", x"f2", x"ee", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"eb", x"ee", x"f0", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f3", x"f2", x"ef", x"ef", x"f0", x"f1", x"f0", x"f2", x"f3", x"f0", 
        x"f1", x"ec", x"dc", x"c8", x"b7", x"b6", x"b9", x"bb", x"c6", x"d7", x"e5", x"ef", x"f2", x"f4", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"eb", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", 
        x"f3", x"f1", x"f1", x"f1", x"ef", x"ef", x"f2", x"f2", x"f0", x"f1", x"f0", x"eb", x"e3", x"da", x"d5", 
        x"d4", x"de", x"e6", x"eb", x"f2", x"f5", x"f4", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"ee", x"f4", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f3", x"f2", x"eb", 
        x"dc", x"cc", x"c8", x"ce", x"d8", x"e4", x"ef", x"f3", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"ef", x"ee", x"ef", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"ee", x"ec", x"ee", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f0", 
        x"f1", x"e0", x"8a", x"47", x"3a", x"5d", x"8d", x"87", x"a7", x"a6", x"99", x"97", x"94", x"90", x"8e", 
        x"8b", x"8a", x"88", x"86", x"83", x"83", x"82", x"7d", x"7b", x"7f", x"7f", x"7c", x"72", x"78", x"84", 
        x"85", x"7f", x"76", x"53", x"36", x"49", x"6b", x"60", x"4c", x"44", x"51", x"69", x"8e", x"b2", x"ca", 
        x"d6", x"da", x"d6", x"d6", x"d5", x"d7", x"db", x"da", x"db", x"db", x"d8", x"d7", x"d7", x"d6", x"d6", 
        x"d8", x"d7", x"d7", x"d7", x"d7", x"d7", x"d6", x"d7", x"d7", x"d7", x"d6", x"d6", x"d6", x"d6", x"d6", 
        x"d6", x"d6", x"d6", x"d6", x"d5", x"d4", x"d7", x"d7", x"d7", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", 
        x"8f", x"8f", x"8e", x"8f", x"8e", x"8c", x"8b", x"8c", x"8c", x"8d", x"8e", x"8e", x"8d", x"8c", x"8e", 
        x"8f", x"8e", x"8c", x"8b", x"8c", x"8c", x"8d", x"8e", x"8d", x"8c", x"8c", x"8d", x"8e", x"8d", x"8c", 
        x"8d", x"8d", x"8d", x"8e", x"8e", x"8c", x"8e", x"8e", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8e", 
        x"8d", x"8d", x"8d", x"8d", x"8d", x"8c", x"8d", x"8c", x"8f", x"90", x"8f", x"8e", x"8d", x"8d", x"8d", 
        x"8d", x"8e", x"8d", x"8d", x"8e", x"8d", x"8f", x"8f", x"8f", x"90", x"8f", x"8e", x"8f", x"8f", x"8f", 
        x"8f", x"8f", x"8f", x"8e", x"8f", x"90", x"90", x"90", x"90", x"91", x"91", x"90", x"90", x"90", x"90", 
        x"90", x"90", x"90", x"90", x"91", x"92", x"91", x"90", x"8f", x"90", x"91", x"90", x"8d", x"8e", x"94", 
        x"94", x"91", x"8a", x"6b", x"54", x"43", x"34", x"19", x"0a", x"08", x"0b", x"1f", x"31", x"3b", x"47", 
        x"51", x"53", x"5e", x"74", x"79", x"76", x"7e", x"70", x"73", x"89", x"96", x"c4", x"db", x"c7", x"a3", 
        x"6f", x"4d", x"3c", x"4d", x"5c", x"69", x"7b", x"81", x"86", x"88", x"87", x"87", x"86", x"88", x"87", 
        x"7b", x"8f", x"dc", x"dd", x"da", x"dc", x"d9", x"e2", x"da", x"d0", x"d1", x"d1", x"d0", x"cf", x"d1", 
        x"d1", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d2", x"d2", x"d2", x"d2", x"d1", x"d0", x"d1", 
        x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"d0", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d3", x"d3", x"d2", x"cf", x"d5", x"d9", x"cf", x"d3", x"d2", x"d5", x"d6", 
        x"d2", x"de", x"f2", x"ed", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"eb", x"ee", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"ef", x"f1", x"f3", x"f1", x"f0", x"f0", x"ef", x"f1", x"f0", x"f0", x"f2", x"f0", 
        x"f0", x"ef", x"f1", x"f3", x"ef", x"e3", x"d4", x"bf", x"b7", x"b4", x"b6", x"c1", x"d0", x"de", x"e8", 
        x"ef", x"f4", x"f4", x"ef", x"ef", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"eb", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f2", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f3", x"f3", x"f0", x"f2", x"f2", x"f2", x"f3", x"f1", x"eb", 
        x"e5", x"df", x"d9", x"d5", x"d8", x"e1", x"eb", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", 
        x"f4", x"f3", x"ef", x"f4", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", 
        x"f0", x"ef", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", 
        x"f1", x"ef", x"e4", x"d3", x"c7", x"c8", x"cf", x"db", x"e8", x"ef", x"f0", x"ed", x"ee", x"f0", x"f0", 
        x"ee", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"ee", x"ec", x"ee", x"f0", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"e5", x"94", x"4b", x"3b", x"56", x"89", x"8b", x"a9", x"a8", x"9a", x"99", x"97", x"92", x"8f", 
        x"8c", x"8b", x"8a", x"87", x"83", x"81", x"80", x"7c", x"79", x"7e", x"83", x"82", x"80", x"7b", x"6f", 
        x"61", x"56", x"4d", x"3a", x"35", x"3f", x"50", x"62", x"81", x"a0", x"c0", x"d2", x"dd", x"dd", x"da", 
        x"d8", x"d9", x"d8", x"dd", x"db", x"d6", x"d9", x"d9", x"da", x"da", x"d9", x"d8", x"d9", x"d8", x"d7", 
        x"d8", x"d8", x"d8", x"d8", x"d7", x"d7", x"d7", x"d8", x"d8", x"d7", x"d5", x"d5", x"d5", x"d6", x"d6", 
        x"d7", x"d7", x"d7", x"d6", x"d5", x"d5", x"d7", x"d7", x"d7", x"d6", x"d6", x"d6", x"d6", x"d6", x"d7", 
        x"90", x"8f", x"8c", x"8c", x"8d", x"8e", x"8f", x"8e", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8e", 
        x"8f", x"8e", x"8d", x"8c", x"8c", x"8c", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8e", x"8f", 
        x"8e", x"8d", x"8d", x"8d", x"8d", x"8d", x"8c", x"8c", x"8c", x"8d", x"8d", x"8d", x"8d", x"8d", x"8f", 
        x"8d", x"8e", x"8f", x"8d", x"8e", x"8d", x"8e", x"8d", x"8e", x"8e", x"8e", x"8f", x"8d", x"8d", x"8c", 
        x"8e", x"8e", x"8d", x"8e", x"90", x"8e", x"8e", x"8f", x"8f", x"8f", x"90", x"90", x"8f", x"8f", x"8f", 
        x"8f", x"8f", x"8f", x"8e", x"8f", x"90", x"90", x"90", x"90", x"91", x"91", x"91", x"90", x"8f", x"90", 
        x"91", x"91", x"90", x"90", x"91", x"91", x"91", x"90", x"90", x"90", x"91", x"90", x"8f", x"8f", x"93", 
        x"94", x"8f", x"93", x"99", x"a0", x"98", x"91", x"51", x"1a", x"26", x"41", x"43", x"3f", x"3c", x"3b", 
        x"39", x"3b", x"3e", x"5d", x"57", x"36", x"4a", x"6e", x"a7", x"ce", x"e1", x"d5", x"a3", x"72", x"4a", 
        x"3c", x"4d", x"59", x"69", x"7b", x"83", x"8a", x"86", x"89", x"89", x"88", x"86", x"84", x"86", x"86", 
        x"7b", x"8e", x"dd", x"de", x"db", x"dc", x"d9", x"e3", x"da", x"d0", x"d1", x"d1", x"d0", x"cf", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d1", x"d1", x"d2", 
        x"d3", x"d4", x"d6", x"d6", x"d5", x"d5", x"d3", x"d2", x"d2", x"d2", x"d1", x"d0", x"d0", x"d0", x"d0", 
        x"d1", x"d1", x"d2", x"d2", x"d3", x"d3", x"d2", x"d0", x"d5", x"da", x"d0", x"d4", x"d3", x"d4", x"d4", 
        x"d2", x"de", x"f1", x"ed", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f1", x"f1", x"f1", x"eb", x"ee", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f1", x"f1", x"ef", x"ef", x"f1", x"f2", x"f3", x"f1", x"ef", x"f2", x"f1", x"f1", x"f2", x"f1", 
        x"f2", x"f3", x"f3", x"f2", x"f3", x"f3", x"f4", x"f4", x"eb", x"dd", x"ce", x"c0", x"b8", x"b2", x"b2", 
        x"bf", x"d4", x"e8", x"f1", x"f4", x"f6", x"f5", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"eb", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"f0", x"f1", 
        x"f2", x"f3", x"f2", x"f3", x"f2", x"f1", x"f2", x"f2", x"f0", x"f3", x"f4", x"f3", x"f1", x"f0", x"f1", 
        x"f3", x"f2", x"ec", x"e2", x"d4", x"cc", x"cd", x"d5", x"e2", x"ed", x"f4", x"f5", x"f3", x"f0", x"f1", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f5", x"f4", 
        x"f3", x"f3", x"ef", x"f3", x"f0", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"f1", x"f2", x"f1", x"ef", x"ef", x"f0", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"ec", x"dd", x"cd", x"c1", x"c3", x"ce", x"e1", x"ef", x"f2", x"f1", x"ee", 
        x"ef", x"f3", x"f2", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ec", x"ef", x"f1", x"f0", x"f0", x"f1", x"f3", x"f4", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"e8", x"9f", x"52", x"39", x"51", x"8f", x"93", x"aa", x"aa", x"9b", x"9a", x"98", x"95", x"91", 
        x"8d", x"8b", x"89", x"87", x"83", x"82", x"84", x"83", x"83", x"86", x"81", x"72", x"5d", x"47", x"32", 
        x"29", x"30", x"41", x"5a", x"7e", x"a0", x"bc", x"d0", x"da", x"de", x"db", x"d7", x"d8", x"d6", x"d9", 
        x"d7", x"d8", x"d9", x"db", x"d8", x"d6", x"da", x"dc", x"d9", x"d8", x"d8", x"d7", x"da", x"d9", x"d7", 
        x"d8", x"d8", x"d8", x"d8", x"d7", x"d7", x"d7", x"d8", x"d8", x"d7", x"d5", x"d4", x"d5", x"d6", x"d7", 
        x"d7", x"d6", x"d6", x"d6", x"d6", x"d5", x"d6", x"d7", x"d7", x"d7", x"d7", x"d7", x"d7", x"d7", x"d7", 
        x"90", x"8f", x"8d", x"8c", x"8d", x"8e", x"8e", x"8f", x"8e", x"8d", x"8c", x"8c", x"8d", x"8f", x"8f", 
        x"8e", x"8e", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8d", x"8e", x"8d", x"8c", x"8d", x"8d", 
        x"8d", x"8e", x"90", x"8e", x"8d", x"8e", x"8d", x"8d", x"8d", x"8d", x"8c", x"8b", x"8c", x"8d", x"90", 
        x"8e", x"8e", x"90", x"8e", x"8e", x"8e", x"8f", x"8d", x"8d", x"8c", x"8d", x"90", x"8f", x"8d", x"8d", 
        x"90", x"90", x"8e", x"8e", x"90", x"8e", x"8d", x"8e", x"8f", x"8e", x"8f", x"92", x"90", x"8f", x"8e", 
        x"8e", x"8e", x"8f", x"90", x"90", x"90", x"90", x"90", x"90", x"90", x"91", x"91", x"90", x"8f", x"90", 
        x"91", x"91", x"90", x"91", x"91", x"90", x"90", x"91", x"91", x"90", x"91", x"91", x"92", x"91", x"92", 
        x"93", x"90", x"91", x"8f", x"93", x"94", x"9f", x"5f", x"25", x"40", x"83", x"7e", x"74", x"6a", x"5d", 
        x"50", x"43", x"38", x"4b", x"4b", x"56", x"96", x"c5", x"df", x"d1", x"a3", x"72", x"4e", x"44", x"4e", 
        x"55", x"60", x"7c", x"a7", x"ac", x"8b", x"88", x"88", x"8d", x"8b", x"88", x"89", x"8a", x"8c", x"89", 
        x"7c", x"90", x"de", x"df", x"db", x"db", x"d8", x"e1", x"da", x"d0", x"d1", x"d1", x"cf", x"cf", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", 
        x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"d3", x"d3", x"d3", x"d2", x"d1", x"d0", x"d1", x"d1", x"cf", 
        x"cf", x"d0", x"d1", x"d1", x"d2", x"d2", x"d1", x"cf", x"d6", x"dc", x"d1", x"d5", x"d3", x"d3", x"d3", 
        x"d0", x"dd", x"f1", x"ed", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", 
        x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ea", x"ed", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"f0", x"ef", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"ef", x"f0", x"f2", x"f1", x"f0", x"f0", x"ef", x"f1", x"ef", x"f0", x"f2", x"f1", 
        x"f0", x"f0", x"f1", x"f3", x"f4", x"f2", x"f1", x"f0", x"f0", x"f1", x"f3", x"f0", x"e7", x"dd", x"ce", 
        x"c5", x"bb", x"b2", x"b5", x"c6", x"df", x"eb", x"ef", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"eb", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f3", x"f3", x"f2", x"f2", x"f4", x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"ec", x"e4", x"dc", x"d2", x"cf", x"d5", x"e2", x"ee", x"f3", x"f3", 
        x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f4", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"ef", x"f3", x"f1", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ee", x"ef", x"ee", x"eb", x"e6", x"d9", x"c8", x"c0", x"c5", x"d7", x"e5", x"f0", 
        x"f2", x"f1", x"f0", x"ee", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ed", x"ef", x"f1", x"f0", x"f0", x"f1", x"f3", x"f5", x"f3", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f0", 
        x"ef", x"e7", x"9a", x"54", x"3c", x"50", x"90", x"8e", x"a3", x"ac", x"9e", x"9b", x"9a", x"97", x"94", 
        x"90", x"8d", x"8b", x"8b", x"8d", x"8d", x"84", x"74", x"64", x"55", x"3e", x"2d", x"33", x"45", x"5d", 
        x"7a", x"9c", x"b4", x"c6", x"cf", x"d8", x"da", x"dc", x"dd", x"d8", x"da", x"d9", x"da", x"d5", x"d7", 
        x"d9", x"d7", x"d6", x"d8", x"d9", x"d9", x"da", x"da", x"d7", x"d8", x"d9", x"d6", x"d9", x"db", x"d9", 
        x"d9", x"d8", x"d8", x"d8", x"d8", x"d8", x"d7", x"d8", x"d8", x"d7", x"d5", x"d4", x"d5", x"d7", x"d7", 
        x"d7", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", x"d6", x"d7", x"d7", x"d7", x"d7", x"d7", x"d7", x"d7", 
        x"8f", x"8f", x"8f", x"8e", x"8f", x"8f", x"8f", x"8d", x"8e", x"8f", x"8e", x"8c", x"8c", x"8d", x"8e", 
        x"8e", x"8e", x"8e", x"8e", x"8d", x"8d", x"8f", x"8f", x"8f", x"8e", x"8d", x"8e", x"8d", x"8d", x"8e", 
        x"8d", x"8e", x"90", x"8e", x"8f", x"8d", x"8f", x"8e", x"8e", x"8f", x"8f", x"8e", x"8d", x"8f", x"8f", 
        x"8d", x"8d", x"8f", x"8e", x"8f", x"90", x"8f", x"8e", x"8d", x"8c", x"8d", x"8f", x"90", x"90", x"8f", 
        x"90", x"90", x"8f", x"8d", x"8e", x"91", x"91", x"90", x"8d", x"8c", x"8e", x"90", x"8f", x"8f", x"8f", 
        x"8f", x"8f", x"90", x"91", x"91", x"8e", x"8f", x"91", x"90", x"8e", x"90", x"8f", x"90", x"92", x"90", 
        x"8f", x"8f", x"90", x"90", x"91", x"91", x"91", x"91", x"91", x"93", x"92", x"91", x"92", x"92", x"91", 
        x"91", x"90", x"91", x"8f", x"8e", x"91", x"9c", x"5c", x"4e", x"63", x"80", x"85", x"83", x"82", x"82", 
        x"7f", x"72", x"5f", x"75", x"9b", x"c5", x"db", x"d5", x"a9", x"74", x"50", x"45", x"4b", x"56", x"66", 
        x"7a", x"9d", x"c0", x"d4", x"bd", x"8c", x"8c", x"8d", x"8d", x"89", x"88", x"89", x"8a", x"8c", x"89", 
        x"7c", x"91", x"dd", x"dd", x"dc", x"dc", x"d9", x"e2", x"d9", x"ce", x"cf", x"cf", x"cf", x"cf", x"d0", 
        x"d2", x"d1", x"d0", x"d1", x"d1", x"d2", x"d1", x"cf", x"d0", x"d2", x"d2", x"d2", x"d1", x"d1", x"d1", 
        x"d1", x"d1", x"d2", x"d2", x"d2", x"d3", x"d2", x"d3", x"d4", x"d0", x"d0", x"d1", x"d1", x"d1", x"ce", 
        x"d0", x"ce", x"cc", x"cf", x"d3", x"d2", x"d2", x"cf", x"d5", x"dc", x"d0", x"d5", x"d5", x"d7", x"d3", 
        x"ce", x"dd", x"f3", x"ed", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", 
        x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"eb", x"eb", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f0", 
        x"ec", x"e4", x"d7", x"c9", x"bd", x"b5", x"b5", x"bf", x"d3", x"e6", x"ef", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f5", x"f2", 
        x"f1", x"f2", x"f4", x"f4", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f1", x"f2", x"f2", x"ec", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f3", 
        x"f3", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f4", x"f3", x"f0", x"ea", x"e5", x"df", x"d5", x"cf", x"d5", x"e4", 
        x"ef", x"f4", x"f2", x"f0", x"f3", x"f3", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f4", x"f4", x"f3", 
        x"f2", x"f2", x"ef", x"f1", x"f2", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f2", x"f2", x"f1", x"ef", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ed", x"ec", x"f1", x"ef", x"ea", x"df", x"d3", x"c4", x"bf", x"cc", 
        x"e1", x"ef", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f3", x"f2", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"ef", x"ee", x"ed", x"ef", x"ef", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f2", x"f2", x"f3", x"f0", 
        x"f0", x"e9", x"a8", x"59", x"3c", x"4a", x"8b", x"92", x"a8", x"c4", x"aa", x"98", x"9b", x"98", x"97", 
        x"94", x"96", x"91", x"82", x"71", x"5f", x"48", x"36", x"32", x"41", x"59", x"71", x"8f", x"a7", x"b8", 
        x"c5", x"d3", x"da", x"dd", x"db", x"db", x"d9", x"da", x"da", x"d9", x"db", x"db", x"da", x"d8", x"d9", 
        x"d9", x"d7", x"d6", x"d7", x"d9", x"d8", x"d7", x"d8", x"d8", x"d7", x"d7", x"d8", x"d9", x"db", x"da", 
        x"db", x"da", x"d9", x"d8", x"d7", x"d7", x"d7", x"d8", x"d8", x"d7", x"d6", x"d6", x"d7", x"d8", x"d8", 
        x"d7", x"d6", x"d5", x"d6", x"d7", x"d8", x"d7", x"d8", x"d8", x"d8", x"d6", x"d6", x"d6", x"d7", x"d7", 
        x"8e", x"8e", x"8f", x"8f", x"90", x"90", x"90", x"8c", x"8c", x"8d", x"8d", x"8d", x"8c", x"8e", x"8e", 
        x"8e", x"8e", x"8e", x"8e", x"8d", x"8d", x"8e", x"8e", x"8e", x"8e", x"8f", x"91", x"8f", x"8e", x"8f", 
        x"8e", x"8e", x"90", x"8f", x"8f", x"8d", x"8d", x"8d", x"8d", x"8f", x"90", x"8f", x"8e", x"8f", x"8e", 
        x"8e", x"8e", x"8f", x"8f", x"8e", x"8f", x"8f", x"8f", x"8e", x"8e", x"8e", x"8d", x"8f", x"90", x"8f", 
        x"8f", x"90", x"90", x"8f", x"8f", x"91", x"92", x"91", x"8d", x"8c", x"8e", x"90", x"90", x"90", x"90", 
        x"90", x"90", x"90", x"90", x"91", x"8f", x"8f", x"91", x"8f", x"8f", x"91", x"8e", x"90", x"92", x"91", 
        x"8e", x"8e", x"91", x"91", x"92", x"92", x"92", x"91", x"91", x"92", x"92", x"92", x"92", x"92", x"92", 
        x"91", x"91", x"91", x"92", x"91", x"92", x"9c", x"60", x"6e", x"7c", x"7b", x"86", x"81", x"80", x"7b", 
        x"75", x"7c", x"a7", x"d0", x"e3", x"da", x"b1", x"7d", x"52", x"42", x"47", x"5c", x"65", x"74", x"9b", 
        x"c6", x"d5", x"d4", x"d7", x"b9", x"8c", x"8a", x"8b", x"8c", x"88", x"88", x"89", x"89", x"8a", x"87", 
        x"7b", x"93", x"de", x"de", x"db", x"dc", x"d8", x"e0", x"d8", x"cd", x"cf", x"cf", x"cf", x"cf", x"d0", 
        x"d3", x"d3", x"d0", x"d0", x"d1", x"d1", x"d1", x"cf", x"d0", x"d2", x"d3", x"d1", x"d1", x"d1", x"d1", 
        x"d1", x"d1", x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", x"d4", x"cf", x"d0", x"d2", x"d1", x"d1", x"d0", 
        x"d3", x"d2", x"ce", x"d0", x"d4", x"d3", x"d2", x"cf", x"d4", x"db", x"cf", x"d4", x"d5", x"d7", x"d2", 
        x"d0", x"dd", x"f1", x"ec", x"ed", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ee", x"f1", x"f1", x"f0", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"ef", x"ef", x"ec", x"ea", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f2", x"f1", x"ea", x"e1", x"d1", x"c4", x"b9", x"b1", x"b7", x"ca", x"e3", x"ef", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f4", x"f5", x"f5", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f0", x"f2", x"f2", x"ec", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", x"f3", 
        x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"ef", x"e6", x"da", x"cd", 
        x"ca", x"d4", x"e7", x"f0", x"f4", x"f1", x"ef", x"f3", x"f4", x"f2", x"f1", x"f2", x"f5", x"f4", x"ee", 
        x"f2", x"f5", x"f7", x"f6", x"f3", x"f2", x"f4", x"f1", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ed", x"ef", x"f0", x"f1", x"f2", x"ee", x"e8", x"d9", x"ca", 
        x"c3", x"c4", x"d7", x"eb", x"f1", x"f0", x"f0", x"f2", x"f0", x"ef", x"f1", x"f3", x"f0", x"ee", x"ef", 
        x"f1", x"ef", x"e9", x"ed", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f4", x"ef", x"f2", x"ef", 
        x"ed", x"ec", x"a7", x"55", x"3a", x"4b", x"90", x"9b", x"b3", x"d6", x"b8", x"9f", x"a4", x"a1", x"97", 
        x"85", x"72", x"56", x"3a", x"28", x"30", x"4f", x"6f", x"8c", x"a7", x"b9", x"c6", x"cb", x"d2", x"d7", 
        x"d8", x"d8", x"da", x"db", x"da", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"da", x"da", x"d9", x"d8", 
        x"d8", x"d7", x"d6", x"d7", x"d9", x"d8", x"d6", x"d7", x"d9", x"d7", x"d8", x"da", x"da", x"d9", x"da", 
        x"db", x"da", x"d9", x"d7", x"d7", x"d7", x"d7", x"d8", x"d7", x"d7", x"d7", x"d8", x"d8", x"d7", x"d7", 
        x"d6", x"d5", x"d5", x"d5", x"d7", x"d8", x"d8", x"d8", x"d8", x"d7", x"d6", x"d5", x"d5", x"d7", x"d7", 
        x"8f", x"8f", x"8f", x"8f", x"8f", x"90", x"90", x"90", x"90", x"8f", x"8f", x"8f", x"8f", x"8f", x"8f", 
        x"8e", x"8e", x"8e", x"8e", x"8e", x"8d", x"8e", x"8f", x"8f", x"8f", x"8f", x"90", x"8d", x"8d", x"8f", 
        x"8e", x"8e", x"90", x"8f", x"90", x"8d", x"8e", x"8e", x"8e", x"8f", x"91", x"91", x"90", x"8d", x"8d", 
        x"8e", x"8f", x"91", x"91", x"8f", x"8e", x"8f", x"8f", x"90", x"8f", x"8e", x"8d", x"8d", x"8d", x"8d", 
        x"8d", x"8f", x"8f", x"8f", x"8f", x"90", x"90", x"8e", x"8e", x"8e", x"90", x"91", x"92", x"91", x"90", 
        x"8f", x"8f", x"90", x"90", x"91", x"91", x"90", x"8f", x"90", x"91", x"91", x"8e", x"8f", x"90", x"8f", 
        x"8e", x"8e", x"8f", x"91", x"91", x"91", x"91", x"91", x"92", x"91", x"91", x"91", x"91", x"92", x"93", 
        x"93", x"92", x"91", x"92", x"92", x"94", x"9e", x"5b", x"71", x"7c", x"73", x"7e", x"7a", x"72", x"7e", 
        x"a3", x"cc", x"df", x"d4", x"ae", x"74", x"52", x"46", x"4f", x"5a", x"60", x"74", x"9c", x"c4", x"d4", 
        x"d1", x"d1", x"cf", x"d4", x"bb", x"90", x"8b", x"8b", x"8d", x"8a", x"89", x"8a", x"89", x"89", x"86", 
        x"7a", x"92", x"dd", x"de", x"dc", x"dd", x"d8", x"e0", x"d7", x"cc", x"cf", x"d0", x"d1", x"d0", x"d0", 
        x"d3", x"d3", x"d1", x"d1", x"d1", x"d0", x"d0", x"cf", x"d0", x"d1", x"d1", x"d1", x"d1", x"d2", x"d1", 
        x"d1", x"d2", x"d2", x"d3", x"d3", x"d3", x"d1", x"cf", x"d1", x"cf", x"d1", x"d3", x"d3", x"d2", x"d0", 
        x"d3", x"d5", x"d3", x"d2", x"d2", x"d1", x"d2", x"cf", x"d3", x"db", x"cf", x"d3", x"d4", x"d4", x"d3", 
        x"d3", x"dc", x"ef", x"ec", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ed", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ec", x"ea", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"f3", 
        x"f1", x"ee", x"ed", x"f0", x"f1", x"f0", x"f0", x"f0", x"ec", x"e2", x"d3", x"c0", x"af", x"b2", x"c2", 
        x"d4", x"e3", x"ec", x"f0", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f3", x"f5", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f0", x"f2", x"f2", x"ed", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"ef", x"ef", x"f2", x"f3", x"f0", 
        x"e8", x"db", x"cf", x"cc", x"d6", x"e5", x"ec", x"ee", x"f1", x"f4", x"f2", x"f0", x"f3", x"f2", x"ef", 
        x"f1", x"f2", x"f1", x"f2", x"f4", x"f5", x"f4", x"f1", x"f1", x"f2", x"f4", x"f4", x"f3", x"f2", x"f2", 
        x"f3", x"f2", x"f0", x"f1", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"e9", x"d9", x"c5", x"bc", x"cb", x"df", x"eb", x"ef", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", 
        x"f0", x"ee", x"eb", x"ef", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f4", x"f2", x"ef", x"f2", x"f1", 
        x"f0", x"f1", x"b5", x"68", x"3e", x"42", x"8b", x"a1", x"b9", x"d8", x"c2", x"97", x"7b", x"5b", x"40", 
        x"33", x"37", x"4a", x"6f", x"8e", x"a9", x"bc", x"c5", x"ca", x"cd", x"d5", x"da", x"da", x"d9", x"d9", 
        x"d9", x"db", x"db", x"da", x"d9", x"d9", x"da", x"db", x"da", x"d8", x"d7", x"d9", x"da", x"da", x"d7", 
        x"d8", x"d8", x"d8", x"d9", x"da", x"d9", x"d7", x"d8", x"da", x"da", x"da", x"db", x"da", x"d9", x"d9", 
        x"d9", x"d9", x"da", x"d9", x"d8", x"d8", x"d8", x"d9", x"d9", x"da", x"d9", x"d8", x"d7", x"d7", x"d7", 
        x"d6", x"d6", x"d6", x"d6", x"d7", x"d8", x"d9", x"d7", x"d7", x"d7", x"d7", x"d6", x"d5", x"d6", x"d7", 
        x"8f", x"8f", x"8f", x"8f", x"8f", x"8f", x"8f", x"8f", x"8e", x"8d", x"8e", x"8e", x"8e", x"8d", x"8e", 
        x"8f", x"8e", x"8e", x"8e", x"8e", x"8d", x"90", x"91", x"90", x"8e", x"8e", x"8f", x"8e", x"8e", x"90", 
        x"8f", x"8f", x"91", x"91", x"90", x"8e", x"8f", x"8f", x"8f", x"8f", x"90", x"91", x"91", x"92", x"91", 
        x"8f", x"8f", x"8f", x"8d", x"8b", x"8e", x"90", x"90", x"90", x"90", x"8f", x"8f", x"8e", x"8d", x"8d", 
        x"8e", x"8e", x"8f", x"8f", x"90", x"91", x"8f", x"8e", x"8e", x"8f", x"90", x"8f", x"92", x"91", x"8f", 
        x"8f", x"8f", x"91", x"91", x"91", x"91", x"90", x"90", x"90", x"91", x"91", x"91", x"92", x"92", x"92", 
        x"93", x"92", x"92", x"91", x"90", x"8f", x"90", x"92", x"93", x"93", x"91", x"91", x"91", x"92", x"93", 
        x"93", x"92", x"93", x"93", x"92", x"94", x"9d", x"58", x"6e", x"77", x"70", x"71", x"7b", x"9c", x"c8", 
        x"de", x"d9", x"b2", x"7d", x"57", x"48", x"4d", x"55", x"65", x"79", x"97", x"c3", x"d8", x"d4", x"d0", 
        x"d1", x"d0", x"d0", x"d4", x"b9", x"8f", x"8c", x"8d", x"8e", x"8b", x"89", x"8a", x"8a", x"8a", x"87", 
        x"79", x"90", x"db", x"dd", x"dd", x"de", x"da", x"e1", x"d6", x"cc", x"d0", x"d1", x"d2", x"d1", x"d1", 
        x"d3", x"d2", x"d1", x"d0", x"d1", x"d1", x"d0", x"d0", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d2", 
        x"d2", x"d2", x"d3", x"d3", x"d2", x"d2", x"d1", x"cf", x"d1", x"d0", x"d0", x"d2", x"d3", x"d1", x"d0", 
        x"d1", x"d4", x"d4", x"d1", x"cf", x"cf", x"d1", x"d0", x"d3", x"da", x"cf", x"d2", x"d3", x"d4", x"d3", 
        x"d2", x"dd", x"f0", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ed", x"ef", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ed", x"ee", x"ef", x"f0", x"ef", x"ef", x"ee", x"f0", x"ec", x"ea", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", x"f0", 
        x"f0", x"ee", x"ef", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"ee", x"e9", x"da", x"c7", 
        x"b9", x"b4", x"ba", x"cb", x"da", x"e2", x"ec", x"f4", x"f6", x"f4", x"f5", x"f5", x"f2", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f5", x"f5", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f0", x"f1", x"f3", x"ed", x"ef", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"ef", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"ef", x"e5", x"d8", x"ce", x"cf", x"d8", x"e7", x"ed", x"f1", x"f3", x"f3", x"f2", x"f0", 
        x"f2", x"f4", x"f4", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f4", x"f3", x"f1", x"f1", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"ee", x"ed", 
        x"f0", x"f1", x"ec", x"e3", x"cc", x"c5", x"cb", x"da", x"e8", x"ec", x"ef", x"f1", x"f1", x"ef", x"ee", 
        x"f0", x"f0", x"ec", x"ee", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f2", x"f1", x"f1", 
        x"ee", x"ef", x"c1", x"72", x"3c", x"45", x"86", x"96", x"86", x"7b", x"5e", x"39", x"36", x"42", x"5f", 
        x"80", x"9c", x"b7", x"ca", x"cf", x"d1", x"d5", x"da", x"dd", x"d8", x"db", x"dc", x"db", x"da", x"d9", 
        x"da", x"db", x"db", x"db", x"da", x"da", x"da", x"d9", x"d9", x"d8", x"d7", x"d9", x"d9", x"d9", x"d8", 
        x"d8", x"d8", x"d9", x"da", x"db", x"da", x"d8", x"d9", x"da", x"da", x"da", x"da", x"d9", x"d8", x"d8", 
        x"d8", x"d8", x"d9", x"d9", x"d9", x"d8", x"d9", x"da", x"da", x"d9", x"d8", x"d8", x"d7", x"d7", x"d7", 
        x"d7", x"d6", x"d6", x"d7", x"d7", x"d8", x"d9", x"d7", x"d6", x"d6", x"d7", x"d7", x"d6", x"d7", x"d7", 
        x"90", x"8f", x"8f", x"8f", x"8f", x"8f", x"8f", x"8c", x"8c", x"8d", x"8e", x"90", x"8f", x"8d", x"8e", 
        x"8f", x"8f", x"8f", x"8f", x"8e", x"8e", x"8f", x"8e", x"8e", x"8e", x"8f", x"91", x"8f", x"90", x"90", 
        x"8f", x"90", x"90", x"91", x"90", x"8f", x"8e", x"8e", x"8e", x"8d", x"8d", x"8e", x"8f", x"8f", x"8e", 
        x"8e", x"8e", x"8f", x"90", x"90", x"90", x"91", x"90", x"8f", x"90", x"90", x"91", x"90", x"8f", x"8f", 
        x"8f", x"8f", x"8e", x"8e", x"90", x"92", x"90", x"8e", x"8e", x"8f", x"8f", x"8e", x"90", x"90", x"8f", 
        x"8f", x"90", x"92", x"93", x"92", x"90", x"90", x"91", x"90", x"90", x"91", x"90", x"91", x"90", x"91", 
        x"91", x"91", x"91", x"91", x"91", x"8f", x"91", x"92", x"94", x"92", x"91", x"91", x"91", x"92", x"93", 
        x"93", x"93", x"93", x"92", x"8e", x"93", x"9d", x"5d", x"6a", x"73", x"7b", x"9a", x"c4", x"e0", x"d6", 
        x"b8", x"89", x"55", x"43", x"4b", x"56", x"5f", x"76", x"97", x"bd", x"d4", x"d4", x"cf", x"d0", x"d0", 
        x"cf", x"ce", x"d1", x"d4", x"b7", x"8b", x"8c", x"8e", x"8e", x"8b", x"8a", x"8b", x"8b", x"8b", x"88", 
        x"7a", x"8f", x"db", x"dd", x"dd", x"de", x"da", x"e1", x"d7", x"cc", x"d0", x"d1", x"d2", x"d1", x"d1", 
        x"d2", x"d1", x"d0", x"d0", x"d2", x"d2", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", 
        x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", x"d1", x"d2", x"d2", x"d0", x"ce", x"d0", x"d3", x"d2", x"d2", 
        x"d2", x"d4", x"d4", x"d0", x"cf", x"d0", x"d1", x"d1", x"d2", x"d9", x"d0", x"d2", x"d3", x"d4", x"d1", 
        x"cf", x"dc", x"f2", x"ed", x"ed", x"ed", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ee", x"f0", x"ed", x"eb", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"f1", x"f0", x"f1", x"f3", x"f4", x"f2", x"f0", x"f1", 
        x"ef", x"e3", x"d0", x"be", x"b5", x"b8", x"c6", x"d0", x"dc", x"e7", x"ee", x"f2", x"f4", x"f6", x"f3", 
        x"f0", x"f0", x"f2", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f3", x"f2", x"f0", x"f1", x"f3", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"ef", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f2", x"f0", x"f2", x"f2", x"ec", x"e1", x"d5", x"ce", x"ce", x"d7", x"e5", x"ec", x"ef", x"f1", 
        x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f3", x"f1", x"f1", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f2", x"f0", 
        x"ee", x"ed", x"ee", x"ee", x"ef", x"e9", x"d8", x"c9", x"c7", x"d3", x"de", x"e8", x"ef", x"f1", x"f0", 
        x"f0", x"f0", x"ec", x"ed", x"ef", x"f0", x"f0", x"f1", x"f2", x"f2", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"ee", x"f0", x"f2", x"f2", 
        x"ee", x"ef", x"ba", x"6c", x"3a", x"3e", x"4e", x"4a", x"3b", x"41", x"54", x"72", x"9c", x"af", x"bd", 
        x"c7", x"cd", x"d7", x"da", x"d8", x"da", x"db", x"da", x"da", x"dd", x"dd", x"dc", x"db", x"d9", x"da", 
        x"d9", x"dc", x"db", x"d9", x"d9", x"d9", x"da", x"d9", x"d8", x"da", x"db", x"d9", x"d8", x"d8", x"da", 
        x"d9", x"d9", x"d9", x"da", x"da", x"da", x"d8", x"d9", x"da", x"d9", x"d8", x"d8", x"d8", x"d9", x"d9", 
        x"d8", x"d8", x"d9", x"d9", x"d9", x"d9", x"d9", x"da", x"da", x"d8", x"d7", x"d7", x"d8", x"d8", x"d7", 
        x"d7", x"d7", x"d7", x"d7", x"d8", x"d9", x"d9", x"d7", x"d6", x"d6", x"d7", x"d8", x"d7", x"d8", x"d7", 
        x"90", x"90", x"8f", x"8f", x"8f", x"8e", x"8e", x"8e", x"8e", x"8f", x"90", x"8f", x"8e", x"8d", x"8e", 
        x"8f", x"8f", x"8f", x"8f", x"8e", x"8e", x"8f", x"8f", x"90", x"90", x"90", x"90", x"8d", x"8d", x"8f", 
        x"8f", x"90", x"90", x"91", x"8f", x"8f", x"90", x"90", x"8f", x"8e", x"8e", x"8f", x"90", x"8f", x"8e", 
        x"8d", x"8e", x"90", x"91", x"91", x"91", x"90", x"8f", x"8f", x"90", x"90", x"91", x"91", x"91", x"91", 
        x"91", x"8f", x"8e", x"8f", x"91", x"91", x"90", x"8e", x"8e", x"8f", x"8f", x"8e", x"91", x"91", x"90", 
        x"90", x"91", x"92", x"92", x"92", x"91", x"90", x"90", x"90", x"91", x"92", x"90", x"91", x"91", x"91", 
        x"91", x"91", x"91", x"92", x"93", x"92", x"92", x"92", x"92", x"92", x"91", x"92", x"92", x"93", x"93", 
        x"93", x"92", x"93", x"95", x"94", x"98", x"98", x"60", x"72", x"98", x"c5", x"df", x"d8", x"b8", x"83", 
        x"56", x"3d", x"4a", x"57", x"64", x"7b", x"9b", x"bd", x"d8", x"d6", x"d1", x"d0", x"d2", x"ce", x"cf", 
        x"d2", x"d0", x"d3", x"d7", x"b8", x"8d", x"8e", x"8f", x"8f", x"8b", x"8a", x"8b", x"8c", x"8c", x"88", 
        x"7b", x"90", x"dc", x"de", x"dd", x"de", x"d8", x"df", x"d9", x"ce", x"d0", x"d1", x"d1", x"d1", x"d1", 
        x"d3", x"d1", x"d0", x"d0", x"d2", x"d2", x"d2", x"d1", x"d1", x"d1", x"d1", x"d3", x"d3", x"d2", x"d1", 
        x"d2", x"d3", x"d3", x"d3", x"d2", x"d1", x"d1", x"d0", x"d0", x"d0", x"ce", x"d1", x"d6", x"d4", x"d4", 
        x"d4", x"d5", x"d4", x"d1", x"d1", x"d2", x"d1", x"d2", x"d2", x"da", x"d2", x"d2", x"d3", x"d3", x"d0", 
        x"cf", x"dd", x"f2", x"ee", x"ee", x"ed", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f1", x"ed", x"eb", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f3", x"f3", 
        x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"f2", 
        x"f2", x"f4", x"f7", x"f5", x"ef", x"e2", x"cb", x"ba", x"b5", x"ba", x"c4", x"d1", x"de", x"ea", x"f2", 
        x"f7", x"f6", x"f4", x"f3", x"f5", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f0", x"f0", x"f3", x"ee", x"ee", x"f0", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"f3", x"f3", x"f2", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", 
        x"f1", x"f0", x"f3", x"f5", x"f1", x"f0", x"f5", x"f4", x"ef", x"e3", x"da", x"d5", x"d2", x"d5", x"de", 
        x"e9", x"ec", x"f2", x"f8", x"f5", x"f3", x"f5", x"f3", x"f2", x"f4", x"f4", x"f4", x"f2", x"f0", x"f2", 
        x"f4", x"f3", x"f0", x"f0", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ee", x"f0", x"f1", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ee", x"ec", x"eb", x"ed", x"f1", x"f0", x"e2", x"d1", x"c7", x"ca", x"d7", x"e4", x"ec", 
        x"f0", x"f0", x"e8", x"eb", x"ef", x"ef", x"f0", x"f1", x"f2", x"f2", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f5", x"f3", x"f5", x"e7", 
        x"cc", x"e0", x"c7", x"7a", x"47", x"4c", x"57", x"70", x"98", x"b3", x"c3", x"ca", x"d7", x"d7", x"da", 
        x"dc", x"dd", x"df", x"da", x"d6", x"da", x"dd", x"db", x"db", x"de", x"de", x"db", x"d9", x"da", x"da", 
        x"da", x"dc", x"da", x"d8", x"d8", x"d9", x"db", x"db", x"d9", x"db", x"db", x"d9", x"d8", x"d9", x"db", 
        x"da", x"da", x"da", x"d9", x"d9", x"d9", x"da", x"da", x"da", x"da", x"d8", x"d7", x"d8", x"da", x"da", 
        x"d8", x"d8", x"d9", x"d9", x"d9", x"d9", x"d9", x"d9", x"d8", x"d7", x"d7", x"d7", x"d8", x"d8", x"d7", 
        x"d7", x"d8", x"d8", x"d8", x"d8", x"d9", x"d8", x"d7", x"d7", x"d7", x"d8", x"d8", x"d8", x"d9", x"d8", 
        x"90", x"90", x"90", x"8f", x"8f", x"8e", x"8e", x"8e", x"8f", x"90", x"8f", x"8e", x"8d", x"8f", x"90", 
        x"8f", x"8f", x"8f", x"8f", x"8f", x"8e", x"8f", x"8f", x"8f", x"8e", x"8f", x"90", x"8d", x"8e", x"8f", 
        x"8f", x"90", x"8f", x"91", x"8e", x"8e", x"8f", x"8f", x"8f", x"8d", x"8e", x"90", x"91", x"8e", x"8d", 
        x"8d", x"90", x"92", x"92", x"92", x"8f", x"8f", x"8f", x"90", x"91", x"91", x"91", x"90", x"91", x"92", 
        x"91", x"90", x"8f", x"90", x"91", x"8f", x"8f", x"8e", x"8e", x"90", x"91", x"91", x"92", x"92", x"91", 
        x"91", x"91", x"91", x"90", x"90", x"93", x"91", x"8f", x"91", x"93", x"91", x"90", x"91", x"91", x"91", 
        x"91", x"90", x"91", x"91", x"92", x"93", x"93", x"93", x"93", x"94", x"93", x"93", x"93", x"93", x"93", 
        x"92", x"91", x"91", x"91", x"8d", x"88", x"92", x"95", x"ba", x"db", x"d6", x"b0", x"84", x"5a", x"42", 
        x"49", x"54", x"62", x"80", x"9d", x"c0", x"d4", x"d5", x"d3", x"d0", x"d3", x"d0", x"d0", x"d0", x"d0", 
        x"d1", x"ce", x"cf", x"d4", x"ba", x"90", x"8d", x"8d", x"8f", x"8d", x"8c", x"8c", x"8c", x"8b", x"87", 
        x"7a", x"8f", x"db", x"de", x"de", x"df", x"da", x"e1", x"da", x"cf", x"d1", x"d0", x"d1", x"d1", x"d1", 
        x"d3", x"d3", x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", x"d0", x"d1", x"d2", x"d3", x"d3", x"d1", x"d0", 
        x"d2", x"d3", x"d3", x"d2", x"d1", x"d1", x"d1", x"d1", x"d1", x"d3", x"d0", x"d1", x"d4", x"d0", x"d1", 
        x"d3", x"d4", x"d3", x"d1", x"d0", x"d0", x"d1", x"d3", x"d3", x"da", x"d3", x"d2", x"d3", x"d3", x"d4", 
        x"d5", x"dd", x"f0", x"ef", x"f1", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", 
        x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"f0", x"f1", x"ef", x"ee", x"ef", x"f0", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"ef", x"f1", x"ed", x"eb", x"f2", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ee", x"f0", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f0", x"ed", x"e4", x"d6", x"c9", x"c1", x"be", x"c0", x"c6", 
        x"d0", x"e1", x"ee", x"f4", x"f5", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f0", x"f0", x"f3", x"ee", x"ee", x"f0", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"ef", x"f0", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"ef", x"ef", x"f0", 
        x"f3", x"f3", x"f0", x"f1", x"ef", x"f0", x"f2", x"ef", x"f1", x"f1", x"f1", x"ef", x"e5", x"dc", x"d8", 
        x"d1", x"ce", x"d5", x"e7", x"f0", x"f3", x"f6", x"f5", x"f4", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f4", x"f3", x"f0", x"f0", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ed", x"f0", x"f2", x"ee", x"ef", x"f0", x"ee", x"ee", 
        x"ef", x"ef", x"ed", x"ee", x"f1", x"f1", x"f0", x"ef", x"ef", x"ee", x"eb", x"de", x"d7", x"d1", x"d1", 
        x"de", x"ea", x"ec", x"ed", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f5", x"dd", 
        x"b7", x"d1", x"d5", x"aa", x"95", x"a3", x"b6", x"c3", x"cb", x"d2", x"d9", x"d8", x"dd", x"dc", x"db", 
        x"da", x"dc", x"dd", x"db", x"d8", x"da", x"db", x"da", x"da", x"da", x"de", x"dd", x"da", x"db", x"d9", 
        x"d6", x"da", x"d9", x"d8", x"da", x"db", x"db", x"da", x"db", x"da", x"d9", x"d9", x"da", x"db", x"db", 
        x"db", x"da", x"d9", x"d8", x"d8", x"d9", x"db", x"da", x"d9", x"db", x"db", x"da", x"da", x"db", x"dc", 
        x"d9", x"d9", x"d8", x"d8", x"d8", x"d9", x"d8", x"d7", x"d7", x"d8", x"d8", x"d8", x"d7", x"d7", x"d7", 
        x"d7", x"d8", x"d8", x"d9", x"d9", x"d8", x"d7", x"d8", x"d9", x"d9", x"d8", x"d8", x"d8", x"d8", x"d7", 
        x"91", x"92", x"91", x"8f", x"8f", x"8f", x"8f", x"8f", x"90", x"91", x"90", x"8f", x"8f", x"90", x"8e", 
        x"8e", x"8e", x"8d", x"8e", x"8d", x"8d", x"8f", x"8f", x"8e", x"8d", x"8f", x"90", x"90", x"90", x"90", 
        x"90", x"90", x"8f", x"8f", x"8e", x"8f", x"8f", x"8f", x"8e", x"8d", x"8e", x"8f", x"8f", x"90", x"8f", 
        x"8e", x"8f", x"90", x"90", x"8f", x"8f", x"90", x"90", x"91", x"91", x"91", x"90", x"90", x"90", x"90", 
        x"90", x"90", x"8f", x"90", x"91", x"8f", x"8f", x"8e", x"8f", x"90", x"92", x"93", x"91", x"91", x"91", 
        x"90", x"8f", x"90", x"90", x"90", x"93", x"91", x"8f", x"92", x"95", x"91", x"92", x"90", x"91", x"93", 
        x"91", x"92", x"92", x"90", x"91", x"94", x"95", x"93", x"91", x"92", x"92", x"92", x"94", x"95", x"93", 
        x"91", x"93", x"8b", x"87", x"8f", x"a3", x"be", x"d6", x"da", x"bb", x"84", x"5a", x"47", x"46", x"54", 
        x"63", x"76", x"9d", x"be", x"d4", x"db", x"d5", x"d3", x"d2", x"d2", x"d2", x"cf", x"cf", x"d0", x"d1", 
        x"d1", x"cd", x"cc", x"d4", x"bd", x"90", x"8b", x"8c", x"8e", x"8c", x"8d", x"8c", x"8c", x"8a", x"86", 
        x"7d", x"8e", x"db", x"dd", x"de", x"e0", x"d9", x"e2", x"d9", x"cf", x"d0", x"d0", x"d0", x"d0", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"cf", x"d0", x"d0", x"d1", x"d2", x"d3", x"d3", x"d1", x"d0", 
        x"d3", x"d3", x"d3", x"d1", x"d0", x"d0", x"d1", x"d1", x"d2", x"d2", x"d0", x"d0", x"d3", x"d1", x"d2", 
        x"d3", x"d2", x"d2", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"da", x"d1", x"d4", x"d4", x"d7", x"d1", 
        x"bb", x"ab", x"b5", x"bf", x"d1", x"e2", x"eb", x"f0", x"f1", x"ef", x"ed", x"ed", x"ed", x"ed", x"ec", 
        x"eb", x"eb", x"ec", x"ed", x"ee", x"ef", x"ed", x"ed", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"ee", x"ed", x"f3", x"f1", 
        x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f0", x"f3", x"f5", x"f6", x"f4", x"ea", x"dd", x"d0", x"c5", 
        x"ba", x"b6", x"bf", x"cd", x"da", x"ec", x"f2", x"f5", x"f6", x"f4", x"f2", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f0", x"f1", x"f2", x"ee", x"ed", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"ef", x"ef", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f4", x"f2", x"ee", 
        x"de", x"d5", x"cf", x"cb", x"cd", x"d7", x"e9", x"f2", x"f5", x"f3", x"ef", x"ef", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f0", x"f2", x"ef", x"ef", x"f1", x"ee", x"ed", 
        x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f2", x"ec", x"e2", x"d9", 
        x"d7", x"d6", x"d4", x"dd", x"e9", x"f0", x"f0", x"ee", x"ed", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", 
        x"ee", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f5", x"e4", 
        x"ce", x"cc", x"ce", x"cb", x"cf", x"d3", x"d8", x"dc", x"dc", x"dd", x"de", x"db", x"da", x"d9", x"da", 
        x"dd", x"df", x"dd", x"dc", x"da", x"db", x"db", x"dd", x"de", x"dc", x"de", x"dc", x"db", x"dc", x"db", 
        x"da", x"d9", x"d9", x"d9", x"da", x"db", x"da", x"d9", x"db", x"da", x"d8", x"d9", x"da", x"db", x"da", 
        x"d9", x"d8", x"d8", x"d8", x"d9", x"db", x"db", x"d9", x"d8", x"da", x"da", x"da", x"da", x"db", x"db", 
        x"d9", x"d9", x"d9", x"d8", x"d8", x"d9", x"d9", x"d7", x"d8", x"d9", x"d9", x"d9", x"d9", x"d8", x"d7", 
        x"d7", x"d7", x"d8", x"d9", x"d9", x"d9", x"d7", x"d9", x"d8", x"da", x"d9", x"d8", x"d8", x"d7", x"d7", 
        x"8f", x"92", x"92", x"8f", x"8f", x"90", x"8e", x"8f", x"91", x"91", x"8f", x"8f", x"90", x"8f", x"8e", 
        x"90", x"8f", x"8e", x"90", x"8f", x"8e", x"90", x"90", x"8e", x"8e", x"8f", x"90", x"8f", x"8f", x"90", 
        x"90", x"8f", x"8e", x"8f", x"90", x"91", x"90", x"8f", x"8f", x"90", x"92", x"91", x"8f", x"91", x"91", 
        x"8f", x"8f", x"90", x"90", x"90", x"90", x"90", x"90", x"90", x"91", x"90", x"8f", x"90", x"90", x"8f", 
        x"90", x"90", x"8f", x"90", x"92", x"91", x"92", x"92", x"91", x"91", x"91", x"92", x"92", x"93", x"93", 
        x"92", x"92", x"93", x"94", x"91", x"93", x"92", x"90", x"94", x"96", x"92", x"93", x"8f", x"90", x"94", 
        x"92", x"92", x"92", x"90", x"93", x"95", x"94", x"91", x"8f", x"90", x"93", x"93", x"93", x"93", x"96", 
        x"8e", x"85", x"8d", x"a9", x"ca", x"de", x"de", x"bb", x"82", x"58", x"3f", x"45", x"55", x"5d", x"76", 
        x"9c", x"c3", x"d4", x"d7", x"d6", x"d2", x"d3", x"d5", x"d2", x"d3", x"d3", x"d2", x"d1", x"d1", x"d2", 
        x"d2", x"d2", x"d0", x"d6", x"bb", x"8e", x"8b", x"8b", x"8a", x"8a", x"8d", x"89", x"89", x"8a", x"87", 
        x"7f", x"90", x"db", x"de", x"de", x"df", x"d5", x"dd", x"d6", x"cf", x"d0", x"cf", x"cf", x"d0", x"d1", 
        x"d0", x"d0", x"d2", x"d3", x"d2", x"d1", x"d0", x"d1", x"d1", x"d1", x"d2", x"d3", x"d4", x"d3", x"d2", 
        x"d3", x"d4", x"d3", x"d1", x"cf", x"d1", x"d1", x"d0", x"d2", x"d0", x"cf", x"d0", x"d1", x"d1", x"d3", 
        x"d4", x"d3", x"d3", x"d2", x"d2", x"d2", x"d1", x"d2", x"cf", x"d9", x"d8", x"da", x"d0", x"ab", x"91", 
        x"9b", x"b6", x"c1", x"b3", x"a8", x"9d", x"a1", x"ae", x"c7", x"dd", x"ed", x"f3", x"f2", x"ef", x"ed", 
        x"ec", x"ec", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", x"ed", x"ee", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f2", x"f1", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"ef", x"ed", x"f1", x"f1", x"ee", 
        x"f0", x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ee", x"ee", x"ed", 
        x"ef", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f4", x"f1", x"ee", 
        x"e7", x"dc", x"cf", x"c1", x"b6", x"b4", x"be", x"d0", x"e4", x"f1", x"f6", x"f6", x"f4", x"f4", x"f4", 
        x"f3", x"f1", x"f1", x"f2", x"f2", x"f0", x"ef", x"f0", x"f3", x"f5", x"f3", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f1", x"ef", x"ee", x"f1", x"f1", x"f1", x"f2", x"f1", x"ee", x"ec", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f4", x"f2", x"ef", x"f0", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ec", x"e5", x"d9", x"ce", x"c6", x"c4", x"d3", x"e8", x"f2", x"f5", x"f5", x"f2", x"f1", 
        x"f4", x"f3", x"ef", x"ed", x"ef", x"f1", x"f1", x"f2", x"f2", x"f2", x"f5", x"f4", x"f2", x"f0", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ee", x"ef", x"f0", x"ef", x"f0", x"f0", x"ee", x"ee", x"f0", x"ee", x"ed", x"ec", x"ef", x"f2", 
        x"f0", x"e4", x"d8", x"c7", x"c4", x"ce", x"e0", x"ee", x"f3", x"f1", x"ef", x"f1", x"f2", x"f1", x"f1", 
        x"ed", x"ef", x"f2", x"ee", x"ef", x"f1", x"f2", x"ef", x"ef", x"f1", x"f6", x"f4", x"ef", x"e7", x"d1", 
        x"cb", x"d2", x"d5", x"d7", x"db", x"de", x"df", x"de", x"dc", x"db", x"db", x"dc", x"db", x"da", x"db", 
        x"dc", x"dd", x"dd", x"dc", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", 
        x"db", x"db", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"da", x"da", x"da", x"da", x"da", x"da", 
        x"da", x"d9", x"d9", x"da", x"db", x"da", x"d8", x"d8", x"d8", x"d8", x"d9", x"d9", x"d9", x"da", x"da", 
        x"db", x"db", x"db", x"d9", x"d8", x"d8", x"d9", x"d8", x"d8", x"d9", x"d9", x"d9", x"d9", x"d9", x"d8", 
        x"d6", x"d6", x"d6", x"d8", x"d9", x"d8", x"d8", x"d8", x"d6", x"d8", x"d9", x"d8", x"d8", x"d8", x"d8", 
        x"90", x"93", x"94", x"92", x"91", x"91", x"8f", x"90", x"92", x"91", x"8d", x"8e", x"91", x"91", x"90", 
        x"8e", x"8f", x"8f", x"8e", x"8e", x"8f", x"8f", x"90", x"8e", x"8e", x"8f", x"90", x"8f", x"8f", x"8f", 
        x"8f", x"8f", x"8f", x"90", x"91", x"91", x"8f", x"8f", x"8f", x"90", x"92", x"91", x"90", x"90", x"91", 
        x"91", x"91", x"90", x"90", x"90", x"90", x"91", x"91", x"90", x"8f", x"8e", x"8e", x"90", x"90", x"90", 
        x"91", x"91", x"90", x"91", x"92", x"90", x"91", x"92", x"93", x"92", x"90", x"8f", x"92", x"92", x"92", 
        x"93", x"93", x"92", x"92", x"90", x"93", x"91", x"90", x"94", x"95", x"92", x"93", x"90", x"91", x"93", 
        x"92", x"92", x"92", x"92", x"93", x"93", x"92", x"91", x"92", x"95", x"95", x"92", x"96", x"90", x"8a", 
        x"8e", x"a5", x"c2", x"d4", x"d9", x"bd", x"87", x"5a", x"47", x"4c", x"55", x"61", x"78", x"9e", x"c5", 
        x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d4", x"d3", x"d0", x"d0", 
        x"d3", x"d2", x"d0", x"d4", x"b9", x"8f", x"8d", x"8b", x"89", x"8d", x"8e", x"8c", x"8a", x"8c", x"8b", 
        x"81", x"95", x"db", x"dd", x"dc", x"dd", x"d8", x"de", x"d7", x"cf", x"d0", x"cf", x"d0", x"d2", x"d3", 
        x"d1", x"d1", x"d2", x"d2", x"d2", x"d1", x"d1", x"d1", x"d1", x"d2", x"d3", x"d4", x"d4", x"d2", x"d2", 
        x"d4", x"d4", x"d4", x"d2", x"d2", x"d2", x"d2", x"d0", x"d1", x"cf", x"cf", x"d1", x"d2", x"d0", x"d3", 
        x"d3", x"d3", x"d4", x"d3", x"d2", x"d1", x"cf", x"ce", x"d4", x"e1", x"ca", x"b2", x"9c", x"a4", x"b6", 
        x"c8", x"dc", x"f0", x"e6", x"dc", x"d2", x"c8", x"b9", x"a6", x"9d", x"a2", x"b1", x"c3", x"d7", x"e2", 
        x"ea", x"ed", x"ef", x"f1", x"f0", x"eb", x"ee", x"ee", x"ec", x"ed", x"ef", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ea", x"ed", x"ee", x"f3", 
        x"f3", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f0", x"eb", x"e4", x"da", x"cf", x"c1", x"b8", x"bc", x"c9", x"d8", x"e7", x"ef", x"f3", 
        x"f3", x"f0", x"f1", x"f4", x"f5", x"f3", x"f2", x"f2", x"f4", x"f4", x"f2", x"f2", x"f4", x"f4", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"ee", x"ec", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"ef", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"ee", x"ee", x"f1", x"f1", x"eb", x"e3", x"da", x"d1", x"c5", x"c4", x"d2", x"e4", x"ed", x"f0", 
        x"f4", x"f3", x"ed", x"ec", x"f2", x"f4", x"f4", x"f4", x"f1", x"ef", x"ef", x"ee", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ee", x"ef", x"f0", x"ef", x"f0", x"f0", x"ee", x"ee", x"f0", x"ee", x"ef", x"ed", x"ed", x"f0", 
        x"f3", x"f1", x"ec", x"e4", x"dd", x"d2", x"c5", x"c7", x"d7", x"e7", x"ec", x"f0", x"f2", x"ef", x"f2", 
        x"ef", x"ef", x"ef", x"f1", x"f1", x"f1", x"f1", x"ed", x"e6", x"db", x"c3", x"aa", x"af", x"cc", x"d8", 
        x"d9", x"df", x"df", x"de", x"dd", x"dc", x"dc", x"dc", x"dd", x"db", x"db", x"dd", x"dc", x"db", x"dc", 
        x"dd", x"dd", x"dc", x"dd", x"dd", x"dc", x"db", x"da", x"da", x"db", x"db", x"db", x"db", x"db", x"db", 
        x"db", x"db", x"da", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"da", x"da", x"da", x"da", x"da", x"da", 
        x"da", x"d9", x"d9", x"da", x"da", x"da", x"d8", x"d8", x"d8", x"d8", x"d9", x"d9", x"d9", x"da", x"da", 
        x"db", x"db", x"da", x"d9", x"d9", x"d8", x"d8", x"d8", x"d9", x"d9", x"da", x"d9", x"d9", x"d8", x"d8", 
        x"d6", x"d6", x"d6", x"d8", x"d9", x"d8", x"d8", x"d8", x"d6", x"d8", x"d8", x"d7", x"d7", x"d8", x"d8", 
        x"91", x"93", x"94", x"92", x"91", x"90", x"8f", x"91", x"93", x"91", x"8d", x"8e", x"91", x"91", x"92", 
        x"90", x"91", x"92", x"8f", x"91", x"92", x"90", x"90", x"8f", x"8f", x"90", x"90", x"90", x"90", x"8f", 
        x"8f", x"90", x"8f", x"90", x"91", x"91", x"91", x"91", x"90", x"91", x"91", x"90", x"8f", x"8e", x"91", 
        x"92", x"92", x"90", x"90", x"90", x"90", x"91", x"91", x"91", x"8f", x"8e", x"8f", x"91", x"90", x"90", 
        x"92", x"92", x"90", x"91", x"91", x"8e", x"8f", x"91", x"93", x"93", x"91", x"90", x"91", x"90", x"91", 
        x"92", x"92", x"91", x"8f", x"91", x"93", x"93", x"91", x"94", x"94", x"92", x"93", x"92", x"92", x"93", 
        x"92", x"92", x"93", x"94", x"94", x"93", x"92", x"90", x"92", x"97", x"99", x"95", x"89", x"87", x"a2", 
        x"be", x"d6", x"d9", x"c6", x"89", x"52", x"33", x"41", x"54", x"61", x"70", x"98", x"c1", x"d5", x"cf", 
        x"d0", x"d1", x"d2", x"d1", x"d1", x"d2", x"d1", x"cf", x"d0", x"d2", x"d3", x"d4", x"d2", x"d1", x"d0", 
        x"d1", x"d2", x"d2", x"d8", x"bb", x"8e", x"8c", x"8c", x"89", x"89", x"8b", x"8b", x"87", x"89", x"8f", 
        x"86", x"91", x"df", x"de", x"db", x"da", x"d4", x"dc", x"d8", x"cf", x"d1", x"d0", x"d0", x"d3", x"d3", 
        x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d0", x"d1", x"d3", x"d5", x"d4", x"d1", x"d1", 
        x"d4", x"d4", x"d4", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"cf", x"cf", x"d0", x"d0", x"ce", x"d2", 
        x"d3", x"d3", x"d4", x"d3", x"d2", x"d2", x"d4", x"d0", x"d5", x"cb", x"9c", x"a7", x"bf", x"cf", x"d3", 
        x"d4", x"e0", x"f3", x"ed", x"ef", x"f2", x"ef", x"ea", x"e5", x"de", x"cf", x"b8", x"a4", x"98", x"9e", 
        x"ad", x"c0", x"d6", x"e6", x"ed", x"ee", x"ed", x"e9", x"e8", x"ec", x"ef", x"ee", x"ed", x"ef", x"ee", 
        x"ee", x"f0", x"f1", x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"ec", x"ef", x"ed", x"f0", 
        x"ef", x"ee", x"f1", x"f0", x"f0", x"f2", x"f3", x"f2", x"f1", x"f0", x"ef", x"ee", x"ee", x"ee", x"f0", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f5", x"f4", 
        x"f2", x"f0", x"f0", x"f1", x"f3", x"f2", x"f1", x"ed", x"e5", x"d7", x"c3", x"b2", x"ae", x"ba", x"d2", 
        x"e5", x"ef", x"f2", x"f3", x"f4", x"f2", x"ef", x"ef", x"f2", x"f4", x"f1", x"f0", x"f5", x"f6", x"f4", 
        x"f0", x"f1", x"f3", x"f4", x"f2", x"f1", x"f1", x"f2", x"f1", x"ee", x"ec", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f2", x"f2", x"f3", x"f5", 
        x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f2", x"f0", x"e5", x"d3", x"c5", x"be", x"bb", x"d0", 
        x"e7", x"f0", x"f0", x"ef", x"f0", x"f2", x"f3", x"f4", x"f2", x"f2", x"f4", x"f5", x"f6", x"f2", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"ee", x"ee", x"f0", x"ee", x"ed", x"ef", x"ee", x"ed", 
        x"ee", x"f0", x"f0", x"ef", x"f0", x"ef", x"e7", x"d8", x"ca", x"c1", x"cd", x"e0", x"ec", x"ee", x"ee", 
        x"ed", x"f2", x"f1", x"f3", x"ed", x"e1", x"cf", x"b1", x"96", x"84", x"8c", x"a9", x"c9", x"db", x"e0", 
        x"df", x"de", x"dd", x"dd", x"dd", x"de", x"de", x"dd", x"dd", x"dc", x"dc", x"dd", x"dd", x"dc", x"dd", 
        x"dd", x"de", x"dd", x"dd", x"dd", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", 
        x"db", x"db", x"db", x"db", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", 
        x"d9", x"d9", x"da", x"db", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"d9", x"da", x"da", x"da", x"da", 
        x"da", x"d9", x"d9", x"da", x"db", x"da", x"d9", x"d8", x"d9", x"da", x"da", x"d9", x"d9", x"d9", x"d8", 
        x"d7", x"d6", x"d7", x"d8", x"d9", x"d8", x"d8", x"d8", x"d7", x"d8", x"d8", x"d8", x"d8", x"d8", x"d8", 
        x"93", x"93", x"93", x"92", x"90", x"90", x"91", x"91", x"92", x"91", x"8f", x"8f", x"91", x"90", x"91", 
        x"90", x"91", x"92", x"90", x"91", x"93", x"91", x"91", x"90", x"90", x"90", x"90", x"91", x"91", x"90", 
        x"91", x"91", x"90", x"90", x"90", x"90", x"91", x"91", x"91", x"91", x"92", x"90", x"8f", x"8f", x"91", 
        x"92", x"92", x"91", x"90", x"90", x"8f", x"90", x"92", x"92", x"91", x"91", x"92", x"93", x"90", x"90", 
        x"92", x"92", x"90", x"91", x"92", x"90", x"8f", x"90", x"92", x"93", x"92", x"91", x"92", x"92", x"92", 
        x"93", x"94", x"92", x"90", x"92", x"94", x"95", x"93", x"93", x"93", x"92", x"94", x"93", x"92", x"93", 
        x"93", x"92", x"94", x"95", x"95", x"94", x"93", x"92", x"93", x"95", x"97", x"90", x"93", x"b8", x"d4", 
        x"d7", x"c3", x"8e", x"57", x"3c", x"43", x"4c", x"59", x"78", x"96", x"c2", x"d4", x"d6", x"d7", x"d4", 
        x"d2", x"d0", x"d2", x"d1", x"d2", x"d4", x"d3", x"d0", x"d1", x"d3", x"d3", x"d1", x"d2", x"d3", x"d3", 
        x"d1", x"d0", x"d1", x"d6", x"b7", x"8a", x"8b", x"8e", x"8c", x"8b", x"8c", x"8c", x"8f", x"8f", x"7b", 
        x"58", x"71", x"d6", x"db", x"dc", x"dd", x"d4", x"dd", x"d8", x"d0", x"d2", x"d0", x"d0", x"d3", x"d3", 
        x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d0", x"d2", x"d3", x"d5", x"d4", x"d1", x"d0", 
        x"d2", x"d3", x"d4", x"d4", x"d3", x"d2", x"d1", x"d2", x"d2", x"d0", x"cf", x"d1", x"d0", x"ce", x"d3", 
        x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"ce", x"d5", x"d9", x"c2", x"d2", x"d6", x"d6", x"d0", 
        x"ce", x"dc", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"ec", x"eb", x"eb", x"e9", x"e1", x"d3", 
        x"c1", x"b1", x"a9", x"a6", x"a9", x"b9", x"cb", x"db", x"e6", x"e9", x"ec", x"f0", x"f1", x"f2", x"f0", 
        x"ec", x"ee", x"f0", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f3", x"ec", x"e7", x"ee", x"f3", 
        x"f2", x"f5", x"f2", x"f0", x"ef", x"f0", x"f1", x"f3", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f3", x"f2", 
        x"f1", x"f2", x"f3", x"f3", x"f1", x"f2", x"f2", x"f3", x"f4", x"f3", x"ef", x"e8", x"dd", x"cd", x"b8", 
        x"ae", x"b4", x"c8", x"db", x"e7", x"ee", x"f1", x"f4", x"f3", x"f3", x"f4", x"f3", x"f1", x"f3", x"f1", 
        x"f1", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"ee", x"ec", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f0", x"f2", x"f4", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f5", 
        x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f1", x"f2", x"f1", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f2", x"f2", x"f1", x"f0", x"ef", x"e7", x"d5", x"c1", 
        x"b9", x"c3", x"d4", x"e3", x"ec", x"ef", x"f0", x"f3", x"f6", x"ec", x"de", x"e2", x"f0", x"f3", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"f0", x"ee", x"ee", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"ed", x"ee", x"f0", x"ed", x"ed", x"eb", x"e4", x"d3", x"c6", x"cb", x"d8", x"e4", 
        x"e5", x"db", x"d1", x"bb", x"9c", x"8d", x"91", x"a6", x"c0", x"d7", x"e6", x"ee", x"ed", x"e2", x"dc", 
        x"dd", x"e0", x"e0", x"e0", x"e0", x"df", x"df", x"df", x"df", x"dd", x"dd", x"dd", x"dd", x"dd", x"de", 
        x"de", x"de", x"de", x"dd", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", 
        x"dc", x"dc", x"dc", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", 
        x"db", x"dc", x"dc", x"db", x"da", x"d9", x"d9", x"d9", x"da", x"da", x"da", x"da", x"da", x"da", x"da", 
        x"da", x"d9", x"d9", x"da", x"db", x"da", x"d9", x"d8", x"d8", x"da", x"da", x"db", x"db", x"da", x"d9", 
        x"d8", x"d7", x"d7", x"d8", x"d9", x"d8", x"d9", x"d9", x"da", x"da", x"da", x"da", x"da", x"db", x"da", 
        x"95", x"94", x"94", x"94", x"92", x"91", x"93", x"93", x"91", x"91", x"92", x"91", x"90", x"91", x"90", 
        x"8f", x"90", x"90", x"8f", x"90", x"91", x"90", x"90", x"91", x"90", x"90", x"90", x"91", x"92", x"90", 
        x"91", x"92", x"91", x"91", x"90", x"8f", x"8f", x"90", x"90", x"91", x"93", x"92", x"91", x"91", x"91", 
        x"91", x"91", x"91", x"90", x"91", x"93", x"93", x"93", x"92", x"91", x"90", x"90", x"90", x"90", x"91", 
        x"93", x"93", x"91", x"91", x"92", x"92", x"92", x"91", x"91", x"92", x"92", x"91", x"91", x"92", x"91", 
        x"92", x"92", x"91", x"91", x"92", x"94", x"95", x"94", x"93", x"93", x"92", x"94", x"94", x"93", x"93", 
        x"94", x"92", x"94", x"93", x"91", x"92", x"93", x"95", x"95", x"96", x"95", x"8f", x"a8", x"cf", x"c7", 
        x"8e", x"4b", x"36", x"48", x"58", x"6c", x"73", x"8f", x"c3", x"dc", x"d5", x"d1", x"d1", x"d1", x"ce", 
        x"d3", x"d2", x"d1", x"d0", x"d2", x"d5", x"d4", x"d3", x"d4", x"d4", x"d3", x"d2", x"d2", x"d4", x"d4", 
        x"d1", x"cf", x"cf", x"d2", x"b7", x"8d", x"8c", x"8c", x"8b", x"8d", x"8e", x"90", x"7b", x"4b", x"20", 
        x"16", x"68", x"d9", x"dc", x"db", x"db", x"d2", x"dc", x"d8", x"d0", x"d1", x"d0", x"d0", x"d2", x"d2", 
        x"d1", x"d1", x"d1", x"d2", x"d2", x"d1", x"d1", x"d1", x"d0", x"d1", x"d3", x"d4", x"d4", x"d2", x"d0", 
        x"d1", x"d3", x"d4", x"d4", x"d3", x"d2", x"d1", x"d1", x"d1", x"d0", x"cf", x"d1", x"d1", x"d0", x"d4", 
        x"d3", x"d2", x"d2", x"d2", x"d2", x"d3", x"d2", x"d1", x"d1", x"da", x"d1", x"d4", x"d2", x"d0", x"d4", 
        x"d2", x"dc", x"f3", x"ed", x"ed", x"f1", x"f0", x"ed", x"ec", x"ec", x"ed", x"eb", x"ec", x"ee", x"ee", 
        x"f0", x"f1", x"ec", x"de", x"cc", x"b3", x"a3", x"9d", x"a5", x"b8", x"cb", x"da", x"e3", x"eb", x"ee", 
        x"ef", x"f1", x"f2", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"f4", x"dd", x"ad", x"c1", x"db", 
        x"e7", x"ee", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f4", 
        x"f4", x"f2", x"f0", x"f2", x"f4", x"f1", x"f3", x"f4", x"f4", x"f2", x"f1", x"f2", x"f6", x"f6", x"f2", 
        x"eb", x"db", x"c1", x"aa", x"af", x"c3", x"d1", x"df", x"ea", x"f1", x"f2", x"f2", x"f6", x"f5", x"f1", 
        x"f1", x"f5", x"f4", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"ee", x"ec", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f2", x"f4", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f2", x"ef", x"ef", x"f1", x"f2", x"f1", x"ef", 
        x"f2", x"f3", x"f3", x"f2", x"f0", x"f0", x"f0", x"f1", x"f3", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"ea", x"d5", x"c5", x"b9", x"ba", x"cf", x"e2", x"ef", x"f0", x"e8", x"d9", x"de", x"ef", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"f0", x"ee", x"ef", x"ef", x"ee", x"ef", 
        x"f1", x"f0", x"ed", x"ed", x"ee", x"ee", x"f0", x"f0", x"ee", x"ed", x"ed", x"e4", x"cc", x"b8", x"a9", 
        x"9d", x"82", x"83", x"90", x"b2", x"d3", x"eb", x"f5", x"f4", x"ee", x"e7", x"dc", x"d5", x"d8", x"df", 
        x"e1", x"de", x"dd", x"de", x"de", x"de", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", x"dd", x"df", 
        x"dd", x"de", x"de", x"dd", x"dc", x"dc", x"dc", x"dd", x"dd", x"dd", x"dd", x"dd", x"dd", x"dd", x"dd", 
        x"dd", x"dc", x"dc", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"da", 
        x"da", x"db", x"dc", x"db", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"d9", x"d9", x"da", 
        x"dc", x"dc", x"db", x"da", x"d9", x"d9", x"d8", x"d8", x"d9", x"da", x"da", x"da", x"da", x"da", x"da", 
        x"d8", x"d7", x"d8", x"d8", x"d8", x"d8", x"da", x"d9", x"dc", x"da", x"da", x"da", x"db", x"db", x"d9", 
        x"94", x"93", x"94", x"95", x"92", x"90", x"92", x"94", x"91", x"90", x"93", x"91", x"8f", x"91", x"91", 
        x"92", x"92", x"92", x"93", x"92", x"91", x"91", x"90", x"91", x"91", x"8f", x"8f", x"91", x"91", x"8f", 
        x"90", x"92", x"92", x"92", x"91", x"90", x"91", x"91", x"91", x"91", x"92", x"92", x"90", x"92", x"92", 
        x"90", x"90", x"91", x"91", x"91", x"92", x"92", x"91", x"91", x"91", x"90", x"90", x"8f", x"90", x"91", 
        x"93", x"93", x"91", x"91", x"91", x"91", x"93", x"93", x"92", x"92", x"92", x"92", x"93", x"93", x"92", 
        x"91", x"91", x"92", x"93", x"91", x"92", x"94", x"94", x"93", x"94", x"95", x"95", x"96", x"93", x"92", 
        x"94", x"92", x"95", x"93", x"91", x"92", x"93", x"94", x"95", x"95", x"93", x"91", x"9f", x"95", x"61", 
        x"37", x"3f", x"52", x"64", x"7d", x"9f", x"c0", x"d6", x"d6", x"d3", x"d2", x"d3", x"d3", x"d4", x"d2", 
        x"d1", x"d0", x"d1", x"d2", x"d3", x"d4", x"d4", x"d3", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d2", 
        x"d1", x"d2", x"d2", x"d4", x"b8", x"8c", x"8c", x"91", x"93", x"8e", x"74", x"4e", x"27", x"15", x"0f", 
        x"1a", x"6b", x"d9", x"db", x"db", x"db", x"d8", x"e0", x"d8", x"d0", x"d1", x"d0", x"d0", x"d2", x"d3", 
        x"d0", x"d0", x"d2", x"d2", x"d2", x"d1", x"d0", x"d1", x"d1", x"d1", x"d2", x"d3", x"d4", x"d2", x"d0", 
        x"d1", x"d5", x"d6", x"d4", x"d3", x"d3", x"d3", x"d2", x"d3", x"d1", x"ce", x"cf", x"d0", x"cf", x"d3", 
        x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", x"d3", x"d1", x"da", x"cf", x"d1", x"d1", x"d3", x"d3", 
        x"d0", x"d9", x"f1", x"ee", x"ee", x"f0", x"f0", x"f1", x"f1", x"ef", x"ef", x"ee", x"ee", x"ed", x"ee", 
        x"ed", x"ee", x"ef", x"ef", x"ee", x"eb", x"e8", x"de", x"ce", x"bc", x"b2", x"ad", x"b0", x"b9", x"c0", 
        x"c8", x"d6", x"e3", x"e9", x"f0", x"f3", x"f3", x"f1", x"f0", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f5", x"c0", x"5a", x"5f", x"76", 
        x"8e", x"a4", x"bc", x"cc", x"de", x"ec", x"f3", x"f4", x"f3", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f2", x"f3", x"f5", x"f5", x"f3", x"f1", x"f1", x"f1", x"f1", x"f4", x"f4", x"f3", 
        x"f3", x"f2", x"ef", x"eb", x"e0", x"d1", x"c4", x"bc", x"bf", x"ca", x"d4", x"dd", x"ea", x"f3", x"f5", 
        x"f3", x"f4", x"f2", x"ef", x"f1", x"f1", x"f1", x"f2", x"f1", x"ee", x"ec", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f2", x"f4", 
        x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f3", 
        x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"ef", x"f0", x"f2", x"ef", x"ef", x"f1", x"f2", x"f1", x"ef", 
        x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"ee", x"f0", x"f2", x"f2", x"f1", 
        x"f1", x"f3", x"f0", x"e2", x"ce", x"c2", x"c1", x"c5", x"cd", x"d4", x"d5", x"df", x"f1", x"f5", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"f0", x"ee", x"ed", x"ed", x"ed", x"f0", 
        x"f1", x"ef", x"f0", x"ee", x"f0", x"f3", x"f0", x"e9", x"dc", x"ca", x"b6", x"a5", x"9c", x"8e", x"7e", 
        x"aa", x"bf", x"c8", x"d0", x"e2", x"ea", x"e7", x"d8", x"c7", x"b9", x"ae", x"a9", x"b5", x"d4", x"e0", 
        x"e2", x"df", x"de", x"de", x"de", x"de", x"de", x"dc", x"dc", x"dc", x"dc", x"db", x"dc", x"dd", x"df", 
        x"dd", x"dd", x"de", x"de", x"dd", x"dd", x"dc", x"dc", x"dd", x"de", x"de", x"de", x"de", x"de", x"de", 
        x"de", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"da", 
        x"d8", x"d9", x"db", x"dc", x"db", x"db", x"dc", x"dc", x"db", x"db", x"da", x"da", x"d9", x"d9", x"d9", 
        x"db", x"dc", x"dc", x"da", x"d9", x"d9", x"da", x"db", x"db", x"db", x"da", x"d9", x"d8", x"d8", x"db", 
        x"d9", x"d8", x"d8", x"d8", x"d8", x"d8", x"da", x"d9", x"dc", x"d9", x"d9", x"d9", x"da", x"da", x"d9", 
        x"93", x"94", x"95", x"96", x"92", x"90", x"92", x"94", x"91", x"90", x"91", x"90", x"8e", x"92", x"91", 
        x"91", x"91", x"91", x"92", x"90", x"8e", x"90", x"90", x"90", x"90", x"8f", x"8f", x"90", x"90", x"8f", 
        x"8f", x"90", x"92", x"92", x"91", x"90", x"91", x"92", x"91", x"90", x"91", x"91", x"8f", x"92", x"92", 
        x"90", x"90", x"91", x"92", x"91", x"91", x"90", x"8f", x"8f", x"91", x"92", x"92", x"92", x"92", x"91", 
        x"92", x"93", x"91", x"92", x"92", x"91", x"92", x"93", x"93", x"93", x"93", x"94", x"94", x"94", x"94", 
        x"94", x"93", x"94", x"96", x"91", x"91", x"92", x"93", x"93", x"94", x"96", x"95", x"95", x"93", x"93", 
        x"94", x"92", x"95", x"96", x"95", x"95", x"94", x"94", x"93", x"94", x"95", x"95", x"8d", x"80", x"73", 
        x"64", x"66", x"76", x"91", x"c1", x"de", x"dc", x"d7", x"d2", x"d1", x"d2", x"d3", x"d2", x"cf", x"d2", 
        x"d4", x"d0", x"d3", x"d3", x"d3", x"d4", x"d3", x"d2", x"d1", x"d0", x"d0", x"d3", x"d4", x"d0", x"d0", 
        x"d2", x"d3", x"d0", x"d3", x"b8", x"91", x"96", x"90", x"77", x"4b", x"1f", x"09", x"10", x"1f", x"27", 
        x"32", x"70", x"d8", x"db", x"db", x"d8", x"d6", x"dc", x"d7", x"cf", x"d0", x"d0", x"d1", x"d3", x"d2", 
        x"d0", x"d0", x"d2", x"d2", x"d2", x"d1", x"d0", x"cf", x"d0", x"d0", x"d2", x"d3", x"d3", x"d2", x"d0", 
        x"d2", x"d4", x"d5", x"d4", x"d3", x"d4", x"d4", x"d1", x"d2", x"d1", x"cf", x"cf", x"d1", x"d1", x"d3", 
        x"d4", x"d4", x"d4", x"d3", x"d2", x"d1", x"d4", x"d2", x"d1", x"d8", x"cc", x"d3", x"d3", x"d4", x"d4", 
        x"d1", x"dd", x"f4", x"ee", x"ec", x"ef", x"f0", x"f1", x"f0", x"ee", x"ee", x"ee", x"ef", x"ee", x"f0", 
        x"f1", x"f1", x"f0", x"ed", x"ec", x"ed", x"f0", x"f1", x"f3", x"f4", x"f0", x"e9", x"d2", x"c4", x"b2", 
        x"a3", x"a6", x"b3", x"be", x"cc", x"d5", x"df", x"ea", x"f0", x"f3", x"f2", x"f0", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", x"f1", x"f1", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"f5", x"cc", x"66", x"6c", x"67", 
        x"5c", x"57", x"5f", x"6c", x"83", x"9d", x"b4", x"ca", x"dc", x"e8", x"f0", x"f5", x"f4", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f0", x"f0", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f0", x"f1", x"f2", x"f2", x"f1", x"f2", x"f3", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f4", x"f5", 
        x"f4", x"f3", x"f1", x"f1", x"f2", x"f3", x"f4", x"f5", x"f3", x"f1", x"f1", x"f4", x"f3", x"f3", x"f5", 
        x"f5", x"f3", x"f2", x"f2", x"f4", x"f7", x"f4", x"ea", x"d6", x"c2", x"b8", x"b8", x"c4", x"cf", x"d9", 
        x"e5", x"ef", x"f4", x"f3", x"f1", x"f1", x"f0", x"f2", x"f3", x"f0", x"ec", x"f1", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f0", x"ef", x"f1", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f3", x"f1", x"f0", x"f1", x"f2", x"f1", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f1", x"f3", x"f4", x"f1", x"f2", 
        x"f4", x"f2", x"f3", x"f3", x"f6", x"f5", x"e9", x"d1", x"c1", x"be", x"c2", x"cf", x"e1", x"eb", x"f2", 
        x"f3", x"f2", x"f1", x"f0", x"f1", x"f3", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"f0", x"ef", x"ed", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"ef", x"ee", x"ed", x"ec", x"ee", 
        x"ef", x"f1", x"f3", x"ee", x"e4", x"d5", x"c1", x"ad", x"99", x"8e", x"92", x"a2", x"c5", x"d1", x"a8", 
        x"df", x"f3", x"de", x"bf", x"b3", x"b0", x"aa", x"9b", x"9a", x"a8", x"c4", x"de", x"eb", x"e8", x"de", 
        x"df", x"df", x"df", x"df", x"df", x"df", x"e0", x"e1", x"e1", x"df", x"dd", x"dc", x"dc", x"dd", x"de", 
        x"dd", x"dd", x"de", x"de", x"dd", x"dd", x"dc", x"dc", x"dc", x"dd", x"de", x"de", x"dd", x"dc", x"dc", 
        x"dd", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"db", x"da", x"da", x"db", x"db", x"da", x"da", x"da", 
        x"d9", x"da", x"db", x"db", x"db", x"db", x"db", x"db", x"da", x"da", x"da", x"da", x"da", x"d9", x"d9", 
        x"da", x"dc", x"dc", x"da", x"d9", x"db", x"dc", x"db", x"dc", x"dc", x"da", x"d8", x"d8", x"d8", x"da", 
        x"da", x"d9", x"d8", x"d9", x"d8", x"d7", x"d9", x"da", x"dc", x"db", x"dc", x"da", x"db", x"db", x"da", 
        x"93", x"94", x"94", x"93", x"91", x"91", x"92", x"92", x"92", x"91", x"90", x"90", x"91", x"93", x"92", 
        x"91", x"91", x"92", x"91", x"91", x"90", x"91", x"90", x"8f", x"91", x"93", x"92", x"90", x"91", x"92", 
        x"90", x"90", x"91", x"92", x"91", x"91", x"90", x"91", x"90", x"90", x"92", x"93", x"91", x"93", x"93", 
        x"92", x"91", x"91", x"93", x"94", x"93", x"93", x"92", x"91", x"91", x"92", x"93", x"94", x"94", x"92", 
        x"91", x"92", x"93", x"94", x"94", x"93", x"93", x"93", x"93", x"93", x"93", x"92", x"92", x"91", x"92", 
        x"93", x"93", x"93", x"94", x"93", x"92", x"91", x"91", x"92", x"93", x"95", x"96", x"93", x"94", x"95", 
        x"94", x"93", x"94", x"95", x"96", x"96", x"95", x"94", x"94", x"95", x"94", x"94", x"96", x"99", x"99", 
        x"94", x"9f", x"bf", x"d5", x"d8", x"d4", x"d6", x"d7", x"d1", x"d2", x"d1", x"d2", x"d3", x"d3", x"d4", 
        x"d3", x"d2", x"d5", x"d2", x"d1", x"d3", x"d4", x"d3", x"d5", x"d0", x"d3", x"d6", x"d3", x"cd", x"d5", 
        x"d4", x"d2", x"ce", x"da", x"c8", x"94", x"67", x"3d", x"1d", x"0c", x"11", x"1c", x"2d", x"3e", x"46", 
        x"44", x"74", x"d8", x"da", x"db", x"d8", x"d4", x"da", x"d8", x"ce", x"d1", x"d0", x"d2", x"d4", x"d2", 
        x"d2", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"cf", x"ce", x"d0", x"d2", x"d2", x"d2", x"d1", x"d1", 
        x"d4", x"d3", x"d3", x"d2", x"d3", x"d3", x"d3", x"d3", x"d2", x"d1", x"cf", x"ce", x"cf", x"d2", x"d3", 
        x"d5", x"d5", x"d4", x"d2", x"d2", x"d2", x"d0", x"d1", x"d2", x"db", x"d0", x"d2", x"d2", x"d4", x"d3", 
        x"d0", x"da", x"f1", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", x"f0", x"f2", x"f3", x"f1", 
        x"eb", x"df", x"d2", x"c7", x"bf", x"b6", x"ae", x"ac", x"b5", x"c3", x"d2", x"e2", x"ee", x"f2", x"f1", 
        x"ef", x"ef", x"ec", x"ed", x"ee", x"ec", x"ee", x"ef", x"ed", x"ee", x"f0", x"ef", x"ee", x"ed", x"ed", 
        x"ed", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"f1", x"f3", x"f3", x"f1", x"ef", x"f0", x"f7", x"c6", x"46", x"41", x"57", 
        x"6b", x"7b", x"7d", x"75", x"6f", x"6a", x"68", x"6e", x"79", x"87", x"9a", x"ba", x"d5", x"e9", x"f4", 
        x"f7", x"f7", x"f6", x"f1", x"ef", x"ef", x"f1", x"f1", x"ec", x"ef", x"f2", x"f0", x"f0", x"f2", x"f1", 
        x"ef", x"f1", x"f2", x"f1", x"f2", x"f5", x"f4", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f3", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f5", x"f7", x"f3", x"eb", x"e2", x"d6", x"ca", x"bf", 
        x"bc", x"c0", x"cc", x"da", x"e9", x"f0", x"f4", x"f4", x"f3", x"ef", x"ec", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f1", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f0", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f4", x"f4", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f1", x"f3", x"ef", x"f3", x"f2", x"f2", x"f2", x"f0", x"e9", x"da", x"cd", x"c6", x"c3", x"c8", 
        x"d8", x"e9", x"f3", x"f4", x"f2", x"f0", x"ef", x"f2", x"f3", x"f0", x"f0", x"f1", x"f1", x"f1", x"f3", 
        x"f1", x"ef", x"f1", x"f3", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"ef", x"e5", x"e8", x"f5", x"f4", x"f0", x"ef", x"ef", x"ec", 
        x"ed", x"ee", x"ee", x"f2", x"ef", x"ed", x"f2", x"ef", x"ea", x"eb", x"ed", x"ec", x"f0", x"f3", x"f0", 
        x"e6", x"cf", x"b2", x"9b", x"97", x"99", x"9f", x"b0", x"c4", x"dc", x"ed", x"f5", x"f5", x"e3", x"91", 
        x"aa", x"ac", x"a8", x"a6", x"a9", x"b5", x"bf", x"bf", x"c6", x"d7", x"f2", x"f5", x"ee", x"e3", x"de", 
        x"df", x"e3", x"e0", x"de", x"de", x"de", x"df", x"df", x"de", x"de", x"de", x"de", x"dd", x"dd", x"dd", 
        x"dd", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", x"dc", x"db", x"dd", x"dd", x"dc", x"db", x"dc", 
        x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", x"db", x"d9", x"da", x"dc", x"db", x"da", x"da", x"da", 
        x"da", x"da", x"d9", x"da", x"dc", x"dc", x"db", x"da", x"d9", x"d9", x"da", x"da", x"db", x"da", x"db", 
        x"db", x"dc", x"dc", x"da", x"d8", x"da", x"dc", x"db", x"dc", x"dc", x"db", x"da", x"db", x"dc", x"da", 
        x"dc", x"dc", x"da", x"db", x"da", x"d8", x"d9", x"dd", x"da", x"d9", x"dc", x"da", x"db", x"d9", x"d8", 
        x"93", x"95", x"95", x"94", x"92", x"91", x"93", x"92", x"91", x"91", x"91", x"90", x"91", x"91", x"92", 
        x"93", x"90", x"90", x"91", x"92", x"92", x"92", x"8f", x"8f", x"92", x"94", x"93", x"92", x"92", x"92", 
        x"92", x"92", x"92", x"92", x"92", x"92", x"90", x"90", x"92", x"92", x"92", x"92", x"92", x"93", x"93", 
        x"91", x"91", x"91", x"92", x"93", x"92", x"92", x"91", x"91", x"92", x"93", x"94", x"93", x"92", x"91", 
        x"91", x"92", x"93", x"94", x"95", x"94", x"94", x"94", x"93", x"93", x"93", x"92", x"92", x"92", x"92", 
        x"92", x"93", x"93", x"92", x"92", x"93", x"94", x"94", x"94", x"95", x"95", x"95", x"94", x"94", x"96", 
        x"95", x"93", x"92", x"94", x"96", x"96", x"95", x"94", x"94", x"94", x"92", x"94", x"96", x"96", x"91", 
        x"99", x"d0", x"dc", x"d7", x"d3", x"d2", x"d6", x"d8", x"d1", x"d3", x"d2", x"d2", x"d3", x"d4", x"d3", 
        x"d2", x"d1", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d2", x"d3", x"d2", x"d2", x"ce", x"d5", 
        x"d5", x"d8", x"d9", x"c7", x"8d", x"47", x"1f", x"11", x"14", x"1e", x"2c", x"3c", x"44", x"47", x"45", 
        x"40", x"74", x"d9", x"da", x"dc", x"d9", x"d6", x"db", x"da", x"cf", x"d1", x"d0", x"d2", x"d4", x"d3", 
        x"d3", x"d4", x"d3", x"d2", x"d2", x"d2", x"d2", x"d1", x"d0", x"d0", x"d1", x"d1", x"d1", x"d1", x"d2", 
        x"d5", x"d5", x"d4", x"d4", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d0", x"cf", x"d0", x"d1", x"d2", 
        x"d4", x"d4", x"d4", x"d2", x"d2", x"d3", x"d2", x"d1", x"d1", x"da", x"cf", x"d2", x"d2", x"d3", x"d3", 
        x"d0", x"da", x"f1", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f1", x"f1", x"eb", x"e2", x"d5", x"c7", x"be", x"b7", x"b1", x"b3", x"b8", x"c1", x"cf", 
        x"dd", x"e8", x"ed", x"f0", x"f1", x"f0", x"f0", x"ef", x"ee", x"ef", x"f1", x"ee", x"ee", x"ed", x"ed", 
        x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f7", x"c4", x"32", x"0d", x"15", 
        x"27", x"36", x"45", x"56", x"6b", x"79", x"7c", x"78", x"71", x"6a", x"6a", x"72", x"7f", x"8f", x"a6", 
        x"bc", x"d3", x"e2", x"ec", x"ef", x"f1", x"f2", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f1", x"f2", x"f4", x"f3", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f2", x"f2", x"f5", x"f0", x"e6", 
        x"d9", x"ce", x"c7", x"c3", x"c2", x"ca", x"d6", x"e4", x"ee", x"ef", x"ec", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f0", x"ef", x"f3", x"f2", x"f3", x"f3", x"f1", x"ef", x"f0", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f3", x"ef", x"f3", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"e5", x"d7", x"cd", 
        x"cc", x"ce", x"d3", x"dc", x"e7", x"ef", x"f2", x"f3", x"f2", x"f0", x"f0", x"f1", x"ef", x"f0", x"f3", 
        x"f2", x"f1", x"f3", x"f4", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f0", x"f0", x"ef", x"f0", x"f2", x"ec", x"c1", x"b6", x"d0", x"e5", x"ed", x"f2", x"f2", x"ee", 
        x"ed", x"ee", x"ef", x"f2", x"ed", x"ed", x"ee", x"ed", x"ef", x"ee", x"eb", x"e5", x"d9", x"c3", x"ab", 
        x"9d", x"9b", x"9b", x"a4", x"bb", x"d1", x"e3", x"ef", x"f2", x"eb", x"de", x"cc", x"b8", x"a9", x"74", 
        x"9d", x"b3", x"c2", x"d0", x"e1", x"ef", x"f4", x"e6", x"d3", x"c4", x"bc", x"b2", x"b1", x"cc", x"e3", 
        x"df", x"e0", x"df", x"de", x"de", x"de", x"de", x"df", x"df", x"de", x"de", x"dd", x"dd", x"dd", x"dd", 
        x"dd", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"db", x"db", x"dd", x"de", x"de", x"dd", x"dc", x"dc", 
        x"dd", x"dc", x"dc", x"dc", x"dc", x"db", x"db", x"db", x"d9", x"da", x"dc", x"db", x"da", x"da", x"da", 
        x"da", x"da", x"d9", x"da", x"dc", x"dc", x"db", x"db", x"db", x"da", x"da", x"d9", x"da", x"db", x"dc", 
        x"db", x"dc", x"db", x"da", x"d9", x"da", x"dc", x"dd", x"db", x"db", x"dc", x"dc", x"db", x"da", x"db", 
        x"dd", x"db", x"da", x"db", x"da", x"da", x"db", x"dc", x"da", x"d9", x"da", x"da", x"da", x"dc", x"dc", 
        x"94", x"95", x"96", x"95", x"93", x"93", x"94", x"94", x"93", x"92", x"92", x"93", x"93", x"90", x"91", 
        x"91", x"90", x"90", x"92", x"93", x"93", x"91", x"90", x"90", x"93", x"95", x"93", x"93", x"91", x"90", 
        x"92", x"94", x"93", x"92", x"91", x"91", x"91", x"91", x"93", x"94", x"92", x"91", x"93", x"91", x"91", 
        x"92", x"93", x"92", x"91", x"91", x"92", x"93", x"93", x"93", x"93", x"93", x"92", x"92", x"92", x"91", 
        x"91", x"92", x"93", x"94", x"94", x"94", x"94", x"94", x"94", x"93", x"93", x"93", x"93", x"94", x"93", 
        x"92", x"93", x"94", x"92", x"93", x"94", x"95", x"96", x"96", x"95", x"95", x"95", x"94", x"95", x"96", 
        x"95", x"93", x"92", x"92", x"93", x"93", x"95", x"95", x"96", x"95", x"92", x"94", x"96", x"97", x"92", 
        x"9a", x"da", x"d3", x"d3", x"d3", x"d4", x"d6", x"d5", x"d1", x"d4", x"d2", x"d2", x"d3", x"d4", x"d3", 
        x"d1", x"d1", x"d3", x"d4", x"d4", x"d4", x"d2", x"d2", x"d4", x"d2", x"d4", x"d5", x"d4", x"d1", x"db", 
        x"e0", x"cd", x"96", x"4b", x"1f", x"13", x"12", x"16", x"2a", x"3d", x"47", x"4b", x"45", x"40", x"41", 
        x"41", x"74", x"d9", x"db", x"db", x"da", x"d7", x"db", x"db", x"d0", x"d1", x"cf", x"d2", x"d5", x"d3", 
        x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d0", x"d0", x"d1", x"d1", x"d1", 
        x"d4", x"d5", x"d6", x"d6", x"d4", x"d2", x"d1", x"d2", x"d3", x"d3", x"d1", x"cf", x"d0", x"d0", x"d1", 
        x"d3", x"d4", x"d4", x"d3", x"d3", x"d3", x"d2", x"d0", x"d1", x"db", x"d1", x"d3", x"d2", x"d3", x"d3", 
        x"d0", x"da", x"f1", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"ef", x"ee", x"ef", x"f1", x"ef", x"ee", x"ee", x"ef", x"f1", 
        x"f1", x"f0", x"ee", x"ed", x"ef", x"ef", x"ee", x"ee", x"ec", x"e8", x"e1", x"d6", x"c7", x"b8", x"ae", 
        x"a6", x"a6", x"b3", x"c6", x"d8", x"e9", x"f5", x"f8", x"f3", x"ee", x"ed", x"ee", x"ef", x"f1", x"f1", 
        x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", x"ed", x"ef", x"f1", x"f0", x"ef", x"f0", x"ef", x"ef", 
        x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f6", x"c7", x"35", x"08", x"03", 
        x"04", x"01", x"07", x"10", x"1b", x"2c", x"43", x"5b", x"70", x"80", x"86", x"85", x"7d", x"73", x"6d", 
        x"6c", x"6f", x"7a", x"97", x"ba", x"da", x"ee", x"f6", x"f7", x"f5", x"f3", x"f1", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f4", 
        x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f0", x"f4", x"f5", 
        x"f3", x"f0", x"ec", x"e6", x"db", x"d0", x"bf", x"b8", x"bf", x"cc", x"d9", x"eb", x"f1", x"f3", x"f2", 
        x"f1", x"f0", x"f1", x"f4", x"f2", x"f2", x"f3", x"f0", x"ef", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f3", x"ef", x"f3", x"f1", x"f0", x"f1", x"f4", x"f1", x"ee", x"f1", x"f5", x"f5", x"f1", 
        x"e9", x"e0", x"d5", x"cc", x"c4", x"c4", x"db", x"eb", x"f6", x"f3", x"ed", x"ed", x"f1", x"ee", x"ef", 
        x"f1", x"f2", x"f3", x"f1", x"ef", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f0", x"ef", x"f0", x"f0", x"ee", x"ef", x"f2", x"c0", x"9d", x"a1", x"ab", x"bb", x"d5", x"ed", x"f6", 
        x"f3", x"ee", x"ec", x"ea", x"ea", x"f0", x"f4", x"f4", x"e9", x"c8", x"a8", x"8c", x"8c", x"9b", x"ae", 
        x"c2", x"d3", x"e3", x"ee", x"f7", x"f7", x"ea", x"d3", x"b7", x"9e", x"9a", x"a4", x"b7", x"c5", x"99", 
        x"c6", x"ef", x"f5", x"f9", x"f6", x"e9", x"d2", x"b4", x"9f", x"96", x"9c", x"af", x"b8", x"cd", x"e4", 
        x"e3", x"e1", x"df", x"df", x"e0", x"df", x"de", x"de", x"df", x"de", x"dd", x"dd", x"dd", x"dc", x"dc", 
        x"dc", x"dc", x"dc", x"dd", x"dd", x"dd", x"dc", x"db", x"dc", x"df", x"df", x"df", x"dd", x"db", x"da", 
        x"db", x"db", x"dc", x"db", x"db", x"db", x"db", x"da", x"d9", x"da", x"dc", x"db", x"da", x"da", x"db", 
        x"db", x"da", x"d9", x"da", x"db", x"db", x"da", x"db", x"dc", x"db", x"da", x"da", x"da", x"da", x"dc", 
        x"dc", x"db", x"db", x"db", x"da", x"db", x"db", x"dc", x"d9", x"d8", x"da", x"db", x"d9", x"d7", x"d8", 
        x"da", x"da", x"d8", x"da", x"db", x"d9", x"db", x"d9", x"d7", x"d7", x"db", x"de", x"e2", x"e7", x"dc", 
        x"94", x"96", x"97", x"96", x"94", x"94", x"95", x"96", x"95", x"94", x"94", x"94", x"94", x"92", x"91", 
        x"90", x"90", x"91", x"92", x"92", x"92", x"92", x"92", x"93", x"93", x"93", x"93", x"93", x"91", x"91", 
        x"92", x"93", x"92", x"91", x"91", x"92", x"93", x"93", x"93", x"93", x"91", x"91", x"94", x"92", x"91", 
        x"93", x"94", x"94", x"92", x"91", x"92", x"94", x"94", x"93", x"93", x"92", x"92", x"92", x"92", x"92", 
        x"92", x"92", x"92", x"93", x"93", x"92", x"93", x"93", x"94", x"95", x"95", x"94", x"94", x"95", x"94", 
        x"94", x"95", x"96", x"95", x"96", x"95", x"94", x"94", x"94", x"94", x"94", x"95", x"96", x"95", x"94", 
        x"94", x"94", x"94", x"92", x"92", x"93", x"94", x"96", x"96", x"95", x"93", x"94", x"97", x"97", x"90", 
        x"96", x"d9", x"d5", x"d4", x"d5", x"d5", x"d3", x"d4", x"d2", x"d2", x"d1", x"d1", x"d2", x"d4", x"d3", 
        x"d3", x"d2", x"d2", x"d1", x"d3", x"d5", x"d2", x"d1", x"d4", x"d3", x"d3", x"d4", x"d7", x"d9", x"c4", 
        x"86", x"49", x"24", x"1a", x"17", x"20", x"35", x"42", x"4a", x"49", x"46", x"45", x"41", x"43", x"42", 
        x"3e", x"72", x"d8", x"d9", x"da", x"d9", x"d6", x"da", x"db", x"d0", x"d1", x"cf", x"d1", x"d4", x"d2", 
        x"d0", x"d1", x"d2", x"d3", x"d2", x"d1", x"d0", x"d1", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d1", 
        x"d2", x"d4", x"d6", x"d7", x"d5", x"d3", x"d2", x"d2", x"d3", x"d3", x"d1", x"d0", x"d0", x"d0", x"d0", 
        x"d2", x"d4", x"d4", x"d3", x"d2", x"d2", x"d2", x"d0", x"d1", x"dc", x"d2", x"d4", x"d1", x"d3", x"d3", 
        x"d0", x"da", x"f1", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"ee", x"ed", x"ef", x"f1", x"ef", x"ed", x"ee", x"ef", x"f0", 
        x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ed", x"ee", x"f0", x"f0", x"ef", x"ee", x"ed", x"ec", x"e5", 
        x"de", x"d3", x"c2", x"b5", x"ad", x"aa", x"ae", x"bb", x"cf", x"e0", x"ea", x"ee", x"ef", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f5", x"ce", x"51", x"36", x"2f", 
        x"23", x"13", x"0c", x"09", x"07", x"05", x"09", x"10", x"19", x"23", x"36", x"4f", x"62", x"73", x"80", 
        x"83", x"7a", x"73", x"71", x"71", x"73", x"7e", x"91", x"ae", x"cc", x"e2", x"eb", x"f0", x"f4", x"f3", 
        x"f2", x"f4", x"f3", x"f1", x"f3", x"f5", x"f3", x"ef", x"f0", x"f1", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f6", x"f3", x"f1", 
        x"f2", x"f5", x"f4", x"f2", x"f2", x"f1", x"eb", x"e5", x"dc", x"ce", x"c0", x"b9", x"c1", x"d0", x"de", 
        x"ea", x"ef", x"f1", x"f2", x"f3", x"f3", x"ef", x"ed", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f3", x"ef", x"f3", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f4", x"f1", x"eb", x"e1", x"d9", x"cd", x"cd", x"d3", x"de", x"e8", x"ef", x"f2", x"f1", x"ef", 
        x"ee", x"f1", x"f4", x"f4", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"ca", x"ab", x"a6", x"9d", x"9d", x"9d", x"a5", x"ba", 
        x"d3", x"e8", x"ee", x"ea", x"e1", x"cc", x"af", x"90", x"87", x"95", x"a9", x"c5", x"d5", x"e2", x"ed", 
        x"f1", x"ee", x"e6", x"d2", x"bb", x"a3", x"9b", x"a7", x"b6", x"c9", x"d8", x"e4", x"ed", x"e7", x"aa", 
        x"be", x"e5", x"d4", x"ba", x"a2", x"99", x"a2", x"b8", x"cb", x"d9", x"e3", x"ea", x"ef", x"e7", x"de", 
        x"df", x"de", x"de", x"df", x"e0", x"df", x"de", x"de", x"df", x"de", x"dd", x"dd", x"dd", x"dc", x"dc", 
        x"dc", x"dc", x"dc", x"dd", x"de", x"de", x"dc", x"db", x"da", x"db", x"dd", x"dd", x"dc", x"db", x"db", 
        x"dc", x"dc", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"dc", x"db", x"da", x"da", x"dc", 
        x"dc", x"da", x"da", x"da", x"db", x"db", x"da", x"da", x"dc", x"dc", x"db", x"db", x"da", x"da", x"db", 
        x"dc", x"db", x"db", x"db", x"db", x"db", x"da", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"d8", 
        x"d9", x"d9", x"d9", x"db", x"db", x"d8", x"dc", x"df", x"e0", x"dd", x"d2", x"c5", x"b9", x"a6", x"98", 
        x"95", x"96", x"97", x"96", x"94", x"94", x"95", x"96", x"95", x"94", x"95", x"94", x"94", x"94", x"92", 
        x"92", x"92", x"90", x"90", x"91", x"93", x"93", x"93", x"94", x"92", x"91", x"93", x"93", x"92", x"92", 
        x"92", x"90", x"8f", x"90", x"91", x"93", x"94", x"93", x"93", x"93", x"92", x"91", x"93", x"94", x"93", 
        x"93", x"92", x"92", x"93", x"93", x"92", x"93", x"93", x"93", x"93", x"94", x"94", x"94", x"93", x"92", 
        x"92", x"93", x"93", x"93", x"92", x"93", x"93", x"93", x"94", x"94", x"95", x"95", x"93", x"94", x"94", 
        x"95", x"96", x"97", x"96", x"96", x"95", x"95", x"94", x"94", x"94", x"94", x"94", x"95", x"94", x"93", 
        x"93", x"95", x"95", x"94", x"94", x"94", x"95", x"95", x"95", x"95", x"94", x"95", x"98", x"98", x"92", 
        x"97", x"d5", x"d7", x"d5", x"d4", x"d3", x"d3", x"d6", x"d3", x"d0", x"d1", x"d2", x"d3", x"d4", x"d4", 
        x"d4", x"d3", x"d4", x"d2", x"d2", x"d3", x"d1", x"d0", x"d1", x"d6", x"d9", x"d9", x"be", x"85", x"44", 
        x"1e", x"18", x"1b", x"28", x"3a", x"42", x"44", x"46", x"46", x"41", x"42", x"44", x"41", x"41", x"41", 
        x"3e", x"70", x"d8", x"d9", x"d8", x"d9", x"d7", x"da", x"db", x"d0", x"d1", x"d0", x"d1", x"d3", x"d1", 
        x"d0", x"d1", x"d2", x"d2", x"d2", x"d1", x"d0", x"d1", x"d1", x"d0", x"d0", x"d3", x"d4", x"d2", x"d0", 
        x"d2", x"d4", x"d6", x"d6", x"d5", x"d4", x"d2", x"d3", x"d3", x"d3", x"d1", x"d0", x"d1", x"d1", x"d0", 
        x"d2", x"d4", x"d4", x"d2", x"d1", x"d1", x"d3", x"d2", x"d1", x"db", x"d1", x"d4", x"d3", x"d4", x"d3", 
        x"d0", x"da", x"f1", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"ee", x"ed", x"ee", x"f1", x"ef", x"ed", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f2", x"f1", x"ef", x"ed", x"ee", x"ef", x"ef", x"ee", x"eb", x"ed", x"f3", x"f1", 
        x"ef", x"ed", x"eb", x"e8", x"e4", x"d9", x"ca", x"b9", x"ab", x"a8", x"af", x"c0", x"ce", x"dc", x"e8", 
        x"ee", x"f1", x"f3", x"f1", x"f1", x"f0", x"ee", x"ec", x"ed", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f6", x"d0", x"5c", x"51", x"54", 
        x"50", x"48", x"3d", x"2f", x"21", x"16", x"0d", x"08", x"04", x"03", x"07", x"0d", x"12", x"1d", x"37", 
        x"53", x"6b", x"78", x"86", x"88", x"81", x"77", x"74", x"6c", x"6f", x"7c", x"95", x"b7", x"d0", x"df", 
        x"e8", x"f1", x"f6", x"f5", x"f2", x"f2", x"f3", x"f1", x"f0", x"f1", x"f3", x"f3", x"f3", x"f2", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f1", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"f3", x"f3", x"f2", x"f3", x"f3", x"ee", x"e7", x"e4", x"db", x"c9", x"b8", 
        x"b4", x"c2", x"d4", x"e2", x"ec", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f3", x"ef", x"f3", x"f1", x"f2", x"f2", x"f2", x"f4", x"f4", x"f2", x"f3", x"f4", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f0", x"ee", x"ee", x"e4", x"d6", x"cc", x"ca", x"d3", x"e1", x"ee", x"f0", 
        x"f1", x"f0", x"ef", x"ef", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"cc", x"ac", x"ab", x"a9", x"a8", x"a7", x"a0", x"9e", 
        x"a4", x"ad", x"a9", x"9a", x"8b", x"93", x"9b", x"94", x"bb", x"e3", x"ea", x"ee", x"ee", x"e9", x"de", 
        x"c8", x"b2", x"a0", x"a0", x"af", x"c3", x"d7", x"e5", x"e8", x"ea", x"eb", x"eb", x"e6", x"d3", x"95", 
        x"82", x"9b", x"9f", x"ae", x"c4", x"d7", x"e4", x"eb", x"ee", x"ed", x"eb", x"e5", x"da", x"d6", x"e0", 
        x"e4", x"e1", x"df", x"df", x"df", x"df", x"de", x"de", x"df", x"de", x"dd", x"dd", x"dd", x"dd", x"dc", 
        x"dc", x"dc", x"dc", x"dd", x"dd", x"dc", x"dc", x"db", x"da", x"da", x"dc", x"dd", x"dc", x"db", x"db", 
        x"dc", x"dc", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"dc", x"db", x"da", x"da", x"db", x"dc", 
        x"dc", x"db", x"da", x"db", x"dc", x"db", x"da", x"da", x"db", x"db", x"dc", x"dc", x"db", x"da", x"db", 
        x"dc", x"db", x"db", x"da", x"da", x"da", x"db", x"dc", x"dc", x"dc", x"db", x"da", x"da", x"db", x"db", 
        x"db", x"da", x"db", x"df", x"e0", x"dd", x"d7", x"c6", x"b3", x"9f", x"92", x"93", x"96", x"9b", x"9f", 
        x"95", x"96", x"97", x"95", x"93", x"93", x"95", x"94", x"94", x"95", x"95", x"94", x"94", x"93", x"93", 
        x"94", x"95", x"94", x"92", x"91", x"93", x"93", x"91", x"94", x"92", x"91", x"93", x"93", x"93", x"93", 
        x"92", x"91", x"92", x"93", x"93", x"93", x"92", x"93", x"94", x"94", x"94", x"92", x"90", x"94", x"94", 
        x"93", x"92", x"92", x"94", x"95", x"94", x"93", x"93", x"92", x"93", x"94", x"94", x"94", x"92", x"92", 
        x"93", x"94", x"94", x"94", x"94", x"95", x"94", x"94", x"94", x"94", x"93", x"93", x"93", x"93", x"93", 
        x"95", x"94", x"95", x"95", x"94", x"95", x"96", x"97", x"97", x"97", x"96", x"93", x"94", x"94", x"93", 
        x"95", x"97", x"96", x"94", x"95", x"95", x"95", x"94", x"94", x"97", x"97", x"96", x"94", x"98", x"92", 
        x"98", x"d4", x"d7", x"d4", x"d2", x"d3", x"d4", x"d6", x"d4", x"d1", x"d2", x"d3", x"d3", x"d5", x"d5", 
        x"d4", x"d3", x"d4", x"d5", x"d4", x"d1", x"d3", x"d6", x"d4", x"d5", x"bd", x"84", x"41", x"21", x"19", 
        x"20", x"29", x"36", x"43", x"4c", x"4b", x"44", x"42", x"42", x"41", x"43", x"45", x"42", x"41", x"3f", 
        x"3b", x"70", x"d9", x"d9", x"d9", x"da", x"d8", x"da", x"da", x"d0", x"d1", x"d0", x"d1", x"d2", x"d0", 
        x"d1", x"d3", x"d3", x"d2", x"d2", x"d1", x"d2", x"d2", x"d1", x"cf", x"d0", x"d3", x"d4", x"d3", x"d1", 
        x"d2", x"d3", x"d5", x"d5", x"d4", x"d2", x"d2", x"d4", x"d3", x"d2", x"d0", x"d0", x"d1", x"d2", x"d1", 
        x"d3", x"d5", x"d5", x"d2", x"d0", x"d0", x"d2", x"d1", x"d2", x"db", x"d0", x"d3", x"d3", x"d4", x"d3", 
        x"d0", x"da", x"f1", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"ee", x"ee", x"ef", x"f1", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"ec", x"ed", x"ef", x"f0", x"ee", x"f1", x"ef", x"ec", x"ee", 
        x"f0", x"ef", x"ee", x"f1", x"f1", x"ea", x"ea", x"eb", x"e4", x"db", x"d0", x"be", x"b7", x"af", x"ae", 
        x"b9", x"cc", x"dc", x"e4", x"ea", x"ef", x"f1", x"ef", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ed", x"f3", x"d1", x"5b", x"4d", x"4f", 
        x"53", x"58", x"58", x"56", x"51", x"4a", x"41", x"30", x"20", x"18", x"11", x"0a", x"08", x"07", x"09", 
        x"0d", x"14", x"20", x"37", x"4f", x"64", x"76", x"84", x"89", x"81", x"76", x"6e", x"6b", x"71", x"7f", 
        x"99", x"b3", x"ca", x"de", x"e8", x"f0", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f4", x"f0", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f4", x"f4", x"f4", x"ef", x"eb", x"ee", x"ef", x"ee", x"eb", 
        x"e3", x"cf", x"c0", x"b2", x"bb", x"cb", x"d9", x"e4", x"eb", x"f0", x"f4", x"f4", x"f4", x"f2", x"f0", 
        x"f0", x"f2", x"f1", x"ef", x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f3", x"ef", x"f3", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"ee", x"e4", x"d4", x"cc", x"cf", x"d6", 
        x"e3", x"ef", x"f2", x"f1", x"ef", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"ef", 
        x"ef", x"f1", x"f1", x"ef", x"ef", x"f2", x"f3", x"cf", x"a5", x"a8", x"ab", x"a5", x"a0", x"93", x"83", 
        x"70", x"65", x"73", x"84", x"97", x"b6", x"ca", x"b1", x"c9", x"e9", x"df", x"cd", x"b8", x"a6", x"a3", 
        x"aa", x"ba", x"d0", x"df", x"e7", x"ec", x"ed", x"ec", x"e4", x"d6", x"c6", x"b4", x"a0", x"9e", x"8a", 
        x"96", x"d3", x"e2", x"eb", x"ee", x"ed", x"eb", x"e5", x"d9", x"cb", x"b2", x"9b", x"94", x"b8", x"e0", 
        x"e4", x"e2", x"e0", x"de", x"de", x"de", x"df", x"df", x"de", x"de", x"de", x"de", x"de", x"dd", x"dd", 
        x"dd", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", x"db", x"db", x"dd", x"dd", x"dd", x"dc", x"dc", 
        x"dc", x"dc", x"dd", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"db", x"da", x"da", x"db", x"dd", 
        x"dd", x"dd", x"db", x"dc", x"dc", x"dc", x"da", x"da", x"db", x"db", x"db", x"db", x"dc", x"db", x"dc", 
        x"db", x"dc", x"dc", x"da", x"d9", x"da", x"dc", x"db", x"da", x"da", x"dd", x"de", x"de", x"dd", x"de", 
        x"de", x"d9", x"d0", x"c4", x"b2", x"a2", x"97", x"93", x"98", x"9b", x"9e", x"a4", x"a7", x"aa", x"ae", 
        x"95", x"96", x"97", x"94", x"93", x"93", x"94", x"91", x"91", x"94", x"95", x"94", x"93", x"93", x"92", 
        x"94", x"98", x"97", x"94", x"92", x"93", x"91", x"90", x"93", x"93", x"93", x"94", x"94", x"93", x"92", 
        x"93", x"94", x"96", x"96", x"93", x"90", x"8f", x"92", x"93", x"94", x"95", x"93", x"8f", x"93", x"94", 
        x"94", x"94", x"94", x"94", x"94", x"95", x"94", x"93", x"93", x"93", x"92", x"93", x"93", x"92", x"93", 
        x"94", x"95", x"95", x"95", x"95", x"96", x"95", x"95", x"94", x"93", x"92", x"92", x"94", x"92", x"93", 
        x"94", x"93", x"93", x"94", x"94", x"95", x"97", x"98", x"99", x"98", x"97", x"93", x"94", x"95", x"94", 
        x"95", x"97", x"96", x"94", x"94", x"95", x"95", x"95", x"96", x"99", x"99", x"96", x"96", x"9b", x"92", 
        x"97", x"d3", x"d6", x"d4", x"d2", x"d5", x"d5", x"d3", x"d3", x"d4", x"d4", x"d4", x"d5", x"d5", x"d5", 
        x"d4", x"d3", x"d1", x"d3", x"d3", x"d6", x"db", x"d1", x"b3", x"75", x"35", x"15", x"1b", x"28", x"27", 
        x"3b", x"49", x"4c", x"46", x"42", x"43", x"42", x"44", x"46", x"40", x"42", x"42", x"3e", x"3b", x"38", 
        x"35", x"70", x"da", x"db", x"da", x"db", x"d9", x"db", x"d9", x"ce", x"cf", x"cf", x"d0", x"d1", x"cf", 
        x"d2", x"d4", x"d3", x"d2", x"d2", x"d2", x"d3", x"d3", x"d1", x"ce", x"d0", x"d2", x"d4", x"d3", x"d3", 
        x"d3", x"d4", x"d4", x"d3", x"d2", x"d1", x"d1", x"d4", x"d4", x"d2", x"d1", x"d0", x"d1", x"d3", x"d1", 
        x"d3", x"d4", x"d4", x"d1", x"d0", x"cf", x"d0", x"d1", x"d3", x"dd", x"d1", x"d3", x"d3", x"d3", x"d2", 
        x"d0", x"d9", x"f0", x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"f0", x"f1", x"ef", x"ef", x"ef", x"f1", x"f0", x"ef", x"ed", x"ed", x"ee", 
        x"ef", x"f0", x"ee", x"ec", x"ed", x"ed", x"ed", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"ee", x"ef", x"f0", x"ed", x"ec", x"ef", x"f4", x"f1", x"e9", x"d8", 
        x"c5", x"b5", x"ab", x"ad", x"b7", x"c6", x"d4", x"df", x"e8", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f5", x"d0", x"58", x"4f", x"54", 
        x"53", x"55", x"54", x"54", x"51", x"52", x"58", x"5a", x"56", x"52", x"4c", x"3b", x"28", x"1e", x"18", 
        x"10", x"0d", x"08", x"06", x"07", x"07", x"14", x"2a", x"43", x"5c", x"73", x"83", x"8c", x"87", x"7a", 
        x"6b", x"66", x"66", x"71", x"8b", x"a9", x"c4", x"d7", x"e4", x"ed", x"f2", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f0", x"f0", x"f0", x"f2", 
        x"f3", x"f2", x"f2", x"f3", x"f1", x"f2", x"f1", x"f3", x"f5", x"f4", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f4", x"f5", x"f4", x"ed", x"dd", x"c7", x"b7", x"b1", x"bc", x"cc", x"db", x"e4", x"ec", x"f1", x"f2", 
        x"f2", x"f2", x"f0", x"ee", x"f0", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f0", x"f2", x"ef", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f4", x"f2", x"f0", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f5", x"f1", x"ee", x"f0", x"f1", x"f0", x"ef", x"e4", x"d7", 
        x"cd", x"d0", x"d8", x"e3", x"eb", x"ef", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f1", x"f0", x"f2", x"f0", x"f1", x"f1", x"ee", x"cf", x"a0", x"94", x"89", x"76", x"68", x"6b", x"7e", 
        x"94", x"a6", x"ac", x"a7", x"99", x"8e", x"96", x"81", x"90", x"a2", x"9b", x"a3", x"b6", x"d0", x"e5", 
        x"f2", x"f4", x"f2", x"e9", x"e3", x"d9", x"c5", x"b2", x"a2", x"9c", x"a4", x"b8", x"d3", x"e7", x"c1", 
        x"b4", x"f0", x"eb", x"e0", x"d5", x"c5", x"ae", x"98", x"8f", x"92", x"ac", x"c9", x"e1", x"ea", x"e4", 
        x"de", x"e0", x"e0", x"df", x"de", x"de", x"df", x"df", x"de", x"de", x"de", x"de", x"dd", x"de", x"de", 
        x"dd", x"dd", x"de", x"dd", x"dc", x"dc", x"dc", x"dd", x"dc", x"d9", x"dc", x"dd", x"de", x"de", x"de", 
        x"df", x"dd", x"dd", x"dc", x"dc", x"db", x"dc", x"dc", x"dc", x"dc", x"db", x"da", x"da", x"db", x"dd", 
        x"de", x"dd", x"db", x"db", x"dc", x"dd", x"da", x"da", x"db", x"dc", x"dc", x"db", x"dc", x"dc", x"dc", 
        x"dc", x"dd", x"dd", x"da", x"d8", x"da", x"dc", x"dd", x"dc", x"dc", x"db", x"dc", x"d4", x"cc", x"be", 
        x"ae", x"9b", x"8f", x"8d", x"92", x"95", x"a3", x"a8", x"aa", x"aa", x"a9", x"ab", x"a8", x"9b", x"84", 
        x"97", x"96", x"97", x"93", x"93", x"92", x"93", x"94", x"92", x"94", x"95", x"94", x"96", x"96", x"93", 
        x"94", x"95", x"94", x"92", x"92", x"93", x"93", x"92", x"91", x"94", x"95", x"94", x"95", x"95", x"93", 
        x"93", x"94", x"95", x"94", x"93", x"93", x"91", x"92", x"93", x"93", x"93", x"93", x"92", x"92", x"93", 
        x"93", x"94", x"93", x"92", x"92", x"93", x"93", x"93", x"95", x"95", x"94", x"95", x"95", x"95", x"96", 
        x"95", x"95", x"95", x"95", x"96", x"94", x"94", x"97", x"94", x"93", x"94", x"91", x"95", x"94", x"94", 
        x"93", x"94", x"94", x"95", x"96", x"95", x"97", x"95", x"97", x"95", x"95", x"95", x"95", x"95", x"95", 
        x"96", x"97", x"96", x"95", x"95", x"96", x"97", x"98", x"98", x"98", x"96", x"95", x"96", x"96", x"92", 
        x"98", x"d5", x"d5", x"d4", x"d5", x"d4", x"d4", x"d3", x"d2", x"d2", x"d3", x"d3", x"d4", x"d5", x"d6", 
        x"d4", x"d4", x"d2", x"d9", x"d6", x"ce", x"a6", x"6e", x"36", x"1a", x"1b", x"25", x"2f", x"3a", x"43", 
        x"49", x"49", x"46", x"44", x"43", x"44", x"44", x"46", x"44", x"3f", x"3f", x"3c", x"39", x"39", x"36", 
        x"35", x"6a", x"db", x"de", x"da", x"da", x"d7", x"dd", x"d9", x"cd", x"cc", x"ce", x"d1", x"d1", x"d1", 
        x"d1", x"d2", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", x"d0", x"cf", x"d2", x"d4", x"d3", x"d3", x"d3", 
        x"d2", x"d3", x"d5", x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"d4", x"d2", x"d1", x"d1", x"d3", x"d1", 
        x"d2", x"d3", x"d2", x"d0", x"d0", x"d0", x"d0", x"d1", x"d0", x"db", x"ce", x"d2", x"d4", x"d3", x"d1", 
        x"d0", x"d8", x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"eb", 
        x"ed", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"ee", x"ea", x"db", x"d0", x"c4", x"bc", x"bb", x"bf", x"c4", x"c7", x"cf", x"dc", x"e7", x"ee", 
        x"f0", x"f0", x"f0", x"f1", x"ef", x"ef", x"f1", x"f1", x"f0", x"ef", x"f3", x"d2", x"5c", x"54", x"57", 
        x"51", x"55", x"56", x"54", x"53", x"54", x"56", x"55", x"54", x"55", x"59", x"59", x"51", x"4d", x"49", 
        x"3e", x"39", x"2e", x"1f", x"19", x"13", x"0d", x"09", x"0a", x"0d", x"17", x"2c", x"44", x"58", x"68", 
        x"7a", x"83", x"83", x"78", x"70", x"6c", x"6c", x"7b", x"8c", x"a1", x"b9", x"cd", x"df", x"ed", x"f1", 
        x"f2", x"f4", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"ef", x"f0", x"f3", x"f0", x"f0", x"f3", x"f2", 
        x"f4", x"f3", x"f1", x"f2", x"f4", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f1", x"f2", x"f3", x"f2", x"f1", x"f2", x"ed", x"ef", x"f2", x"f1", x"f1", 
        x"f2", x"f3", x"f0", x"ee", x"f0", x"f2", x"ef", x"e5", x"d3", x"c5", x"ba", x"bb", x"c2", x"cd", x"d8", 
        x"e4", x"ec", x"f1", x"f3", x"f4", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f4", x"f5", x"f4", x"f2", 
        x"f3", x"f4", x"f2", x"f1", x"f0", x"f0", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"ee", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"ef", x"e8", x"db", x"d3", x"d5", x"d8", x"df", x"e7", x"ee", x"f2", x"f4", x"f2", x"f1", x"ef", x"f1", 
        x"f4", x"f0", x"ee", x"e3", x"d1", x"c3", x"b8", x"a2", x"82", x"75", x"80", x"8e", x"9f", x"a9", x"a8", 
        x"a9", x"a1", x"96", x"8e", x"86", x"81", x"7b", x"5f", x"66", x"8e", x"9d", x"be", x"de", x"f0", x"ee", 
        x"e2", x"d4", x"c3", x"b4", x"ad", x"aa", x"ac", x"ba", x"cf", x"e4", x"ed", x"ef", x"ee", x"e7", x"b8", 
        x"92", x"bb", x"ad", x"a2", x"9b", x"a1", x"b2", x"c8", x"da", x"e8", x"e8", x"e0", x"d3", x"d2", x"df", 
        x"e1", x"e0", x"e0", x"df", x"de", x"de", x"de", x"df", x"df", x"de", x"dd", x"dc", x"dd", x"de", x"df", 
        x"de", x"de", x"de", x"de", x"dd", x"dd", x"de", x"de", x"dd", x"dc", x"dc", x"dd", x"dd", x"dc", x"dc", 
        x"dc", x"dc", x"dc", x"dc", x"da", x"da", x"dc", x"de", x"db", x"da", x"da", x"db", x"dc", x"dd", x"dd", 
        x"dc", x"dc", x"da", x"d9", x"da", x"dc", x"db", x"da", x"dc", x"dd", x"dc", x"da", x"db", x"de", x"de", 
        x"db", x"dc", x"dd", x"de", x"e0", x"df", x"db", x"d7", x"d0", x"c1", x"b1", x"a8", x"9d", x"98", x"95", 
        x"95", x"9c", x"a4", x"a8", x"ad", x"aa", x"a8", x"a7", x"9d", x"89", x"70", x"5a", x"46", x"29", x"1e", 
        x"98", x"97", x"97", x"93", x"94", x"94", x"94", x"95", x"94", x"94", x"95", x"93", x"96", x"96", x"94", 
        x"92", x"93", x"94", x"94", x"94", x"94", x"93", x"93", x"93", x"95", x"94", x"92", x"94", x"96", x"94", 
        x"94", x"93", x"93", x"93", x"94", x"95", x"93", x"93", x"94", x"94", x"94", x"94", x"93", x"93", x"94", 
        x"94", x"94", x"94", x"93", x"93", x"95", x"94", x"94", x"95", x"95", x"94", x"97", x"97", x"95", x"94", 
        x"94", x"95", x"94", x"94", x"95", x"95", x"94", x"96", x"95", x"95", x"95", x"93", x"96", x"96", x"94", 
        x"94", x"94", x"94", x"95", x"94", x"94", x"97", x"96", x"97", x"95", x"95", x"96", x"96", x"96", x"96", 
        x"97", x"97", x"97", x"96", x"95", x"96", x"98", x"98", x"99", x"98", x"97", x"96", x"97", x"96", x"93", 
        x"98", x"d5", x"d5", x"d2", x"d6", x"d2", x"d4", x"d5", x"d2", x"d0", x"d2", x"d5", x"d4", x"d4", x"d6", 
        x"d5", x"d7", x"d6", x"cf", x"a8", x"6a", x"36", x"15", x"1a", x"24", x"30", x"3e", x"44", x"46", x"46", 
        x"43", x"43", x"44", x"43", x"42", x"41", x"41", x"40", x"3f", x"3c", x"3c", x"3a", x"39", x"3a", x"38", 
        x"36", x"69", x"d9", x"de", x"d9", x"da", x"d8", x"de", x"da", x"ce", x"cd", x"cf", x"d2", x"d2", x"d3", 
        x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"d3", x"d3", x"d1", x"d0", x"d2", x"d4", x"d3", x"d2", x"d2", 
        x"d2", x"d3", x"d4", x"d4", x"d3", x"d3", x"d4", x"d4", x"d5", x"d4", x"d2", x"d1", x"d2", x"d3", x"d1", 
        x"d2", x"d3", x"d2", x"d0", x"d0", x"d1", x"d0", x"d1", x"d0", x"db", x"ce", x"d2", x"d4", x"d2", x"d1", 
        x"d1", x"da", x"f2", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ec", 
        x"ee", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"ec", x"e1", x"d3", x"c6", x"b8", x"b5", x"b7", x"bd", x"c7", 
        x"d1", x"d8", x"e3", x"eb", x"f0", x"f2", x"f2", x"f1", x"f0", x"ef", x"f1", x"d3", x"5f", x"58", x"58", 
        x"54", x"58", x"58", x"57", x"56", x"56", x"56", x"55", x"52", x"51", x"53", x"54", x"50", x"4a", x"52", 
        x"55", x"52", x"53", x"4a", x"45", x"3e", x"32", x"27", x"1e", x"14", x"0c", x"08", x"07", x"0d", x"17", 
        x"2e", x"45", x"56", x"66", x"79", x"84", x"83", x"7f", x"74", x"6e", x"6f", x"7a", x"8b", x"a2", x"b6", 
        x"cb", x"e0", x"ec", x"f2", x"f5", x"f4", x"f1", x"f0", x"ef", x"f2", x"f5", x"f0", x"ef", x"f2", x"f1", 
        x"f2", x"f2", x"f2", x"f1", x"ef", x"ed", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f1", x"f2", x"f3", x"f2", x"f1", x"f3", x"ec", x"ef", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f1", x"f0", x"f2", x"f3", x"f4", x"f4", x"f4", x"f2", x"e8", x"da", x"ca", x"bd", x"b9", 
        x"bf", x"c8", x"d2", x"e1", x"ed", x"f2", x"f3", x"f5", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f0", x"f1", x"f1", x"ee", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"ef", 
        x"f2", x"f5", x"f3", x"eb", x"e6", x"d9", x"d1", x"d2", x"d8", x"e1", x"e9", x"ee", x"f1", x"f4", x"ef", 
        x"ee", x"cd", x"b7", x"b1", x"a0", x"a3", x"b1", x"ba", x"ac", x"a9", x"ac", x"ad", x"a9", x"9c", x"8f", 
        x"8d", x"84", x"7c", x"7b", x"7a", x"86", x"94", x"7f", x"7d", x"9e", x"8e", x"8b", x"9c", x"ae", x"b2", 
        x"ab", x"a8", x"aa", x"b1", x"c5", x"dc", x"ec", x"f3", x"f2", x"ea", x"e1", x"cf", x"bd", x"b3", x"8f", 
        x"6a", x"9f", x"a9", x"bd", x"d4", x"e5", x"ec", x"e5", x"d5", x"c7", x"b9", x"ac", x"a5", x"b7", x"db", 
        x"e5", x"e0", x"df", x"df", x"df", x"df", x"df", x"df", x"e0", x"de", x"dd", x"dd", x"de", x"df", x"e0", 
        x"de", x"de", x"df", x"df", x"de", x"de", x"dd", x"dc", x"dc", x"dd", x"dd", x"dd", x"dd", x"dc", x"db", 
        x"db", x"dc", x"dc", x"dc", x"da", x"da", x"dc", x"dd", x"d9", x"da", x"dc", x"dd", x"de", x"dd", x"db", 
        x"d9", x"da", x"da", x"d9", x"d9", x"db", x"da", x"db", x"dd", x"dd", x"db", x"da", x"dc", x"e0", x"e1", 
        x"df", x"df", x"df", x"da", x"d0", x"c4", x"b9", x"a9", x"a2", x"9b", x"95", x"96", x"9b", x"a4", x"aa", 
        x"a9", x"ae", x"ac", x"a6", x"9c", x"8a", x"6e", x"5a", x"42", x"27", x"19", x"1d", x"26", x"2f", x"3f", 
        x"9a", x"97", x"96", x"95", x"96", x"96", x"95", x"94", x"94", x"95", x"95", x"94", x"95", x"95", x"93", 
        x"92", x"93", x"95", x"96", x"96", x"94", x"93", x"93", x"94", x"94", x"93", x"92", x"93", x"95", x"95", 
        x"94", x"93", x"93", x"93", x"94", x"95", x"94", x"94", x"93", x"94", x"94", x"95", x"95", x"94", x"94", 
        x"95", x"95", x"95", x"95", x"94", x"97", x"95", x"94", x"95", x"94", x"94", x"97", x"97", x"95", x"93", 
        x"93", x"95", x"95", x"94", x"94", x"95", x"94", x"95", x"96", x"96", x"95", x"93", x"97", x"97", x"97", 
        x"95", x"94", x"94", x"95", x"95", x"94", x"94", x"93", x"95", x"96", x"97", x"97", x"96", x"96", x"97", 
        x"97", x"98", x"98", x"95", x"96", x"98", x"98", x"98", x"99", x"98", x"97", x"98", x"99", x"99", x"96", 
        x"9a", x"d6", x"d2", x"c9", x"d3", x"d1", x"d2", x"d6", x"d2", x"cf", x"d5", x"d2", x"d2", x"d4", x"dc", 
        x"de", x"d1", x"9c", x"59", x"2c", x"0f", x"23", x"30", x"2b", x"33", x"40", x"48", x"46", x"42", x"43", 
        x"46", x"46", x"45", x"44", x"42", x"40", x"3d", x"3b", x"3a", x"38", x"37", x"37", x"3a", x"3f", x"3f", 
        x"3c", x"6b", x"da", x"df", x"d9", x"d9", x"d7", x"dc", x"dc", x"d1", x"cf", x"d0", x"d1", x"d1", x"d2", 
        x"d4", x"d5", x"d4", x"d3", x"d3", x"d3", x"d4", x"d3", x"d2", x"d0", x"d2", x"d3", x"d2", x"d2", x"d1", 
        x"d2", x"d3", x"d4", x"d3", x"d3", x"d3", x"d3", x"d5", x"d5", x"d4", x"d3", x"d2", x"d3", x"d3", x"d1", 
        x"d3", x"d3", x"d2", x"d1", x"d1", x"d1", x"d1", x"d1", x"cf", x"db", x"cf", x"d3", x"d4", x"d2", x"d1", 
        x"d1", x"da", x"f1", x"ee", x"ed", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ed", 
        x"ef", x"f1", x"f1", x"ef", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f1", x"ef", x"ef", 
        x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"f0", x"f1", x"ef", 
        x"ed", x"ec", x"ed", x"f0", x"ee", x"ec", x"ec", x"ee", x"f1", x"f3", x"ee", x"e7", x"db", x"ce", x"c3", 
        x"ba", x"b6", x"b8", x"bc", x"c3", x"d0", x"e1", x"ee", x"f4", x"f2", x"f5", x"d2", x"59", x"4f", x"55", 
        x"56", x"56", x"57", x"58", x"58", x"55", x"56", x"58", x"5a", x"5a", x"59", x"55", x"58", x"4a", x"63", 
        x"6a", x"4d", x"52", x"51", x"53", x"58", x"55", x"52", x"4b", x"42", x"37", x"29", x"1f", x"16", x"0b", 
        x"05", x"05", x"09", x"11", x"23", x"39", x"4e", x"62", x"74", x"86", x"8f", x"85", x"74", x"6c", x"6e", 
        x"73", x"80", x"93", x"ac", x"c9", x"e1", x"f0", x"f6", x"f7", x"f4", x"f1", x"ef", x"ef", x"f1", x"f0", 
        x"f0", x"f2", x"f4", x"f3", x"f1", x"f1", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f1", x"f2", x"f3", x"f2", x"f1", x"f3", x"ec", x"ee", x"f1", x"f1", x"f1", 
        x"f2", x"f4", x"f2", x"f3", x"f6", x"f5", x"f3", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f1", x"e6", 
        x"d7", x"c8", x"bb", x"b4", x"b5", x"c2", x"d6", x"e6", x"f1", x"f6", x"f6", x"f5", x"f4", x"f3", x"f3", 
        x"f4", x"f4", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f1", x"ee", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"f1", x"f4", x"f6", x"ef", x"e5", x"db", x"d2", x"cf", x"d3", x"d9", x"e7", x"f3", 
        x"e6", x"7c", x"9e", x"be", x"d7", x"eb", x"f7", x"ea", x"b7", x"9c", x"90", x"8a", x"84", x"7f", x"7c", 
        x"81", x"86", x"91", x"9c", x"a2", x"a5", x"a8", x"8b", x"73", x"86", x"7b", x"76", x"74", x"77", x"7f", 
        x"88", x"a1", x"cd", x"ed", x"f8", x"f6", x"e5", x"d1", x"b7", x"a3", x"a1", x"a2", x"a4", x"b3", x"ae", 
        x"88", x"e4", x"f2", x"ec", x"d8", x"bd", x"a9", x"a3", x"a4", x"a6", x"b1", x"bf", x"d1", x"e1", x"e8", 
        x"df", x"df", x"e0", x"df", x"df", x"df", x"df", x"df", x"e0", x"de", x"dd", x"de", x"df", x"e0", x"e0", 
        x"de", x"de", x"e0", x"df", x"de", x"de", x"dd", x"dc", x"dd", x"df", x"df", x"de", x"de", x"dd", x"dc", 
        x"db", x"dd", x"dd", x"dd", x"db", x"db", x"dc", x"dd", x"db", x"dc", x"dd", x"dc", x"dc", x"db", x"dc", 
        x"dc", x"dc", x"db", x"da", x"dc", x"dd", x"dd", x"da", x"d9", x"db", x"df", x"e4", x"e3", x"de", x"d7", 
        x"ca", x"bb", x"ae", x"a4", x"9c", x"98", x"96", x"93", x"9a", x"a2", x"a8", x"af", x"b1", x"b0", x"a7", 
        x"91", x"79", x"5e", x"4a", x"35", x"1c", x"10", x"17", x"26", x"35", x"45", x"4d", x"52", x"51", x"52", 
        x"99", x"97", x"95", x"96", x"96", x"96", x"95", x"95", x"96", x"96", x"96", x"95", x"95", x"95", x"95", 
        x"94", x"94", x"96", x"97", x"96", x"93", x"92", x"93", x"92", x"92", x"93", x"94", x"92", x"92", x"94", 
        x"95", x"95", x"95", x"95", x"95", x"95", x"95", x"94", x"93", x"92", x"92", x"93", x"93", x"94", x"94", 
        x"95", x"96", x"96", x"95", x"95", x"95", x"94", x"94", x"96", x"94", x"93", x"94", x"96", x"96", x"94", 
        x"94", x"96", x"96", x"95", x"94", x"95", x"95", x"95", x"97", x"97", x"95", x"95", x"98", x"98", x"98", 
        x"96", x"96", x"94", x"94", x"96", x"97", x"97", x"97", x"97", x"96", x"96", x"96", x"96", x"97", x"97", 
        x"98", x"97", x"98", x"96", x"97", x"99", x"98", x"98", x"9a", x"98", x"98", x"99", x"99", x"9a", x"96", 
        x"99", x"d5", x"d4", x"cd", x"d5", x"d4", x"d3", x"d4", x"d5", x"d7", x"d7", x"d1", x"d8", x"db", x"c4", 
        x"97", x"5b", x"2b", x"14", x"18", x"28", x"32", x"4d", x"51", x"39", x"37", x"40", x"46", x"44", x"43", 
        x"45", x"45", x"44", x"41", x"3f", x"3c", x"3b", x"3a", x"3a", x"3d", x"3c", x"3b", x"3e", x"41", x"41", 
        x"3d", x"6c", x"d9", x"df", x"d8", x"d8", x"d7", x"da", x"db", x"d1", x"d0", x"d0", x"d0", x"d0", x"d1", 
        x"d3", x"d4", x"d3", x"d2", x"d1", x"d2", x"d2", x"d2", x"d2", x"d1", x"d2", x"d3", x"d3", x"d2", x"d0", 
        x"d2", x"d3", x"d4", x"d3", x"d3", x"d3", x"d4", x"d5", x"d4", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", 
        x"d3", x"d4", x"d3", x"d1", x"d1", x"d2", x"d1", x"d1", x"cf", x"da", x"cf", x"d3", x"d3", x"d2", x"d0", 
        x"cf", x"d7", x"ef", x"ed", x"ed", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"ef", 
        x"f0", x"f1", x"f0", x"ef", x"ef", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ee", x"ef", x"f1", x"f0", x"ee", x"f0", x"f1", x"ef", 
        x"ee", x"ed", x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", 
        x"e7", x"df", x"d4", x"cd", x"c7", x"bf", x"bb", x"be", x"c5", x"ce", x"e0", x"c9", x"62", x"55", x"57", 
        x"59", x"53", x"50", x"4f", x"51", x"54", x"57", x"59", x"5a", x"57", x"5b", x"67", x"5e", x"45", x"61", 
        x"7a", x"4e", x"51", x"51", x"51", x"55", x"54", x"53", x"54", x"55", x"55", x"51", x"4d", x"46", x"3b", 
        x"33", x"28", x"1b", x"12", x"0d", x"09", x"0b", x"13", x"22", x"30", x"47", x"5c", x"6e", x"7b", x"80", 
        x"7f", x"7c", x"77", x"75", x"77", x"82", x"94", x"a9", x"c1", x"d9", x"e8", x"ef", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f2", x"f1", x"f3", x"ec", x"ee", x"f1", x"f1", x"f1", 
        x"f3", x"f4", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f1", x"f2", x"f4", x"f3", x"f2", x"f3", x"f5", 
        x"f4", x"f0", x"e7", x"db", x"d1", x"c7", x"be", x"b8", x"bd", x"cd", x"de", x"e9", x"f3", x"f6", x"f4", 
        x"f2", x"f3", x"f4", x"f2", x"f2", x"f3", x"f5", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f1", x"ee", x"f0", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"ef", x"ec", x"e5", x"de", x"d5", x"ce", x"cf", 
        x"c5", x"5b", x"bc", x"ec", x"ed", x"e1", x"d3", x"b9", x"8d", x"88", x"8a", x"8d", x"94", x"98", x"99", 
        x"9d", x"a3", x"a2", x"9d", x"96", x"8c", x"83", x"68", x"5b", x"7a", x"7e", x"8b", x"90", x"95", x"97", 
        x"96", x"98", x"9c", x"a6", x"ac", x"a5", x"9d", x"a3", x"ad", x"b9", x"c7", x"d5", x"e3", x"e8", x"d3", 
        x"80", x"b5", x"ad", x"a5", x"ab", x"b0", x"b6", x"c3", x"d4", x"e1", x"e9", x"e6", x"d7", x"cc", x"dd", 
        x"e2", x"e0", x"e0", x"e0", x"df", x"df", x"df", x"df", x"e0", x"df", x"de", x"dd", x"de", x"df", x"e0", 
        x"df", x"df", x"de", x"de", x"de", x"de", x"dd", x"dd", x"de", x"de", x"de", x"de", x"de", x"dd", x"dd", 
        x"dd", x"dd", x"dd", x"dd", x"db", x"db", x"dc", x"dc", x"dc", x"dd", x"dd", x"dc", x"dc", x"dc", x"dd", 
        x"de", x"dd", x"da", x"db", x"dd", x"de", x"dd", x"df", x"df", x"db", x"d3", x"c5", x"b6", x"a8", x"a1", 
        x"9e", x"9a", x"98", x"9a", x"a0", x"a5", x"aa", x"ad", x"b2", x"ab", x"9c", x"8a", x"71", x"5a", x"44", 
        x"2e", x"1d", x"13", x"1d", x"2a", x"34", x"3f", x"44", x"49", x"4b", x"48", x"48", x"4d", x"57", x"62", 
        x"97", x"97", x"95", x"97", x"96", x"96", x"95", x"96", x"97", x"94", x"92", x"93", x"93", x"95", x"95", 
        x"95", x"95", x"96", x"97", x"95", x"93", x"93", x"94", x"92", x"91", x"94", x"96", x"93", x"91", x"94", 
        x"95", x"96", x"96", x"96", x"95", x"93", x"93", x"93", x"93", x"92", x"92", x"93", x"94", x"93", x"93", 
        x"95", x"95", x"96", x"96", x"96", x"95", x"94", x"94", x"96", x"94", x"92", x"93", x"95", x"96", x"95", 
        x"94", x"96", x"96", x"95", x"94", x"95", x"96", x"95", x"97", x"97", x"95", x"96", x"97", x"97", x"97", 
        x"97", x"96", x"95", x"95", x"97", x"98", x"98", x"99", x"97", x"96", x"95", x"96", x"96", x"97", x"97", 
        x"97", x"97", x"97", x"96", x"98", x"9a", x"97", x"98", x"9a", x"99", x"97", x"98", x"97", x"98", x"95", 
        x"97", x"d3", x"d6", x"d4", x"d3", x"d5", x"d5", x"d1", x"d2", x"d5", x"d8", x"de", x"cb", x"97", x"53", 
        x"2b", x"17", x"17", x"29", x"39", x"45", x"34", x"4f", x"61", x"3c", x"36", x"41", x"46", x"41", x"41", 
        x"44", x"41", x"3f", x"3c", x"3a", x"39", x"39", x"3a", x"3b", x"3e", x"40", x"41", x"43", x"44", x"41", 
        x"3c", x"6a", x"d6", x"dd", x"d8", x"d9", x"da", x"db", x"d8", x"ce", x"ce", x"cf", x"d0", x"d1", x"d2", 
        x"d3", x"d4", x"d2", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d1", x"d2", x"d4", x"d2", x"d0", 
        x"d2", x"d3", x"d4", x"d4", x"d3", x"d4", x"d4", x"d5", x"d4", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", 
        x"d3", x"d4", x"d3", x"d2", x"d1", x"d2", x"d1", x"d1", x"ce", x"da", x"cf", x"d3", x"d3", x"d3", x"d1", 
        x"ce", x"d6", x"ed", x"ec", x"ed", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", 
        x"f0", x"f1", x"ef", x"ef", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"ee", x"ef", x"ef", x"f0", x"ee", 
        x"ee", x"f0", x"ef", x"ef", x"ed", x"e6", x"dc", x"d1", x"cb", x"c2", x"bf", x"ab", x"5f", x"4d", x"49", 
        x"52", x"58", x"57", x"58", x"57", x"53", x"50", x"52", x"54", x"54", x"64", x"7a", x"63", x"4a", x"65", 
        x"78", x"4d", x"50", x"50", x"52", x"55", x"56", x"56", x"51", x"4f", x"4e", x"4f", x"54", x"56", x"55", 
        x"56", x"54", x"49", x"40", x"34", x"29", x"1e", x"11", x"0b", x"07", x"0b", x"14", x"20", x"2d", x"3e", 
        x"58", x"6d", x"7e", x"89", x"87", x"7c", x"73", x"6f", x"72", x"7f", x"93", x"ad", x"c8", x"e0", x"ec", 
        x"f2", x"f5", x"f4", x"f3", x"f2", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f2", x"f1", x"f3", x"ec", x"ef", x"f1", x"f2", x"f2", 
        x"f3", x"f4", x"f2", x"f4", x"f5", x"f4", x"f2", x"f2", x"f3", x"f5", x"f3", x"f2", x"f5", x"f5", x"f2", 
        x"f1", x"f1", x"f3", x"f3", x"f3", x"ef", x"e6", x"d9", x"cb", x"bf", x"b5", x"b6", x"c3", x"d7", x"ea", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f2", x"ee", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f0", x"f2", 
        x"f2", x"f0", x"ef", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"ee", x"e9", x"e4", x"dc", 
        x"c6", x"56", x"84", x"b9", x"aa", x"aa", x"b3", x"ba", x"9f", x"a1", x"a2", x"a2", x"a5", x"a8", x"a8", 
        x"9c", x"8f", x"80", x"76", x"74", x"7a", x"82", x"70", x"65", x"95", x"99", x"98", x"a0", x"a0", x"95", 
        x"88", x"79", x"69", x"64", x"6f", x"79", x"86", x"a8", x"d3", x"ed", x"ea", x"dc", x"c4", x"aa", x"99", 
        x"5c", x"a1", x"b4", x"c5", x"d6", x"e3", x"ea", x"e8", x"dd", x"cf", x"bd", x"b1", x"a6", x"ae", x"d9", 
        x"e5", x"e0", x"e0", x"e0", x"e0", x"df", x"df", x"e0", x"e0", x"df", x"de", x"dc", x"dc", x"de", x"df", 
        x"df", x"df", x"de", x"de", x"de", x"de", x"de", x"de", x"de", x"dd", x"dd", x"de", x"de", x"de", x"de", 
        x"de", x"de", x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", x"e1", x"e0", x"dd", x"db", x"dc", x"dd", x"dd", 
        x"df", x"df", x"e0", x"e4", x"e3", x"db", x"d3", x"c7", x"b6", x"a6", x"9c", x"9b", x"9d", x"9a", x"9c", 
        x"a2", x"a3", x"a7", x"ae", x"b2", x"ad", x"a1", x"8e", x"74", x"51", x"3a", x"28", x"1a", x"0f", x"0b", 
        x"07", x"06", x"1a", x"4a", x"50", x"45", x"3f", x"43", x"4e", x"59", x"62", x"6b", x"77", x"7f", x"82", 
        x"94", x"96", x"95", x"97", x"95", x"95", x"94", x"95", x"97", x"94", x"94", x"96", x"94", x"95", x"96", 
        x"96", x"96", x"96", x"95", x"95", x"95", x"93", x"92", x"94", x"93", x"94", x"95", x"95", x"94", x"95", 
        x"95", x"96", x"96", x"96", x"95", x"95", x"95", x"96", x"95", x"94", x"93", x"92", x"91", x"92", x"93", 
        x"94", x"95", x"96", x"96", x"96", x"96", x"95", x"95", x"96", x"94", x"93", x"93", x"95", x"96", x"95", 
        x"95", x"95", x"95", x"95", x"93", x"94", x"96", x"95", x"96", x"95", x"95", x"97", x"96", x"96", x"97", 
        x"97", x"97", x"96", x"95", x"98", x"98", x"96", x"96", x"95", x"97", x"98", x"96", x"96", x"96", x"96", 
        x"97", x"97", x"97", x"95", x"99", x"9b", x"98", x"97", x"9b", x"99", x"97", x"98", x"97", x"98", x"95", 
        x"96", x"d2", x"d6", x"d2", x"d3", x"d2", x"d0", x"d7", x"de", x"d9", x"c4", x"89", x"4b", x"21", x"15", 
        x"1c", x"2a", x"3b", x"47", x"4f", x"4a", x"35", x"48", x"5e", x"44", x"38", x"3d", x"48", x"43", x"3e", 
        x"3d", x"3b", x"3a", x"3a", x"3a", x"3b", x"3c", x"3e", x"40", x"42", x"45", x"45", x"44", x"44", x"40", 
        x"3b", x"68", x"d4", x"dc", x"d8", x"da", x"dc", x"dc", x"d9", x"cf", x"cf", x"d0", x"d0", x"d1", x"d3", 
        x"d4", x"d4", x"d3", x"d3", x"d2", x"d1", x"d0", x"d0", x"d1", x"d1", x"d0", x"d2", x"d5", x"d3", x"d2", 
        x"d3", x"d4", x"d5", x"d4", x"d4", x"d4", x"d5", x"d4", x"d3", x"d1", x"d2", x"d2", x"d2", x"d1", x"d2", 
        x"d3", x"d4", x"d3", x"d2", x"d2", x"d2", x"d2", x"d1", x"ce", x"d9", x"cf", x"d3", x"d3", x"d3", x"d2", 
        x"cf", x"d7", x"ee", x"ed", x"ee", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ec", x"ed", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ed", x"ef", x"f1", x"f0", x"ed", x"e8", x"e4", x"dd", x"c3", x"b7", x"9b", 
        x"7d", x"62", x"4d", x"4b", x"4d", x"52", x"57", x"59", x"5a", x"5f", x"6d", x"75", x"59", x"47", x"66", 
        x"61", x"50", x"52", x"50", x"52", x"52", x"55", x"56", x"51", x"50", x"50", x"50", x"4e", x"50", x"53", 
        x"5a", x"60", x"60", x"5d", x"54", x"51", x"51", x"46", x"3c", x"30", x"24", x"18", x"0f", x"0c", x"0e", 
        x"11", x"18", x"25", x"3b", x"58", x"70", x"7f", x"85", x"83", x"7b", x"72", x"6a", x"6c", x"75", x"8f", 
        x"a6", x"c1", x"dd", x"eb", x"f1", x"f5", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f2", x"f1", x"f3", x"ec", x"f0", x"f3", x"f2", x"f2", 
        x"f3", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f4", x"f2", x"f2", x"f3", 
        x"f3", x"f4", x"f2", x"f1", x"f2", x"ef", x"f0", x"f3", x"f2", x"eb", x"e4", x"da", x"c7", x"b7", x"b2", 
        x"bb", x"cb", x"e4", x"ed", x"f2", x"f4", x"f3", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"ef", x"f2", x"f2", x"ef", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f1", x"f0", x"f2", x"f3", x"f0", x"f0", x"f3", x"f4", x"f2", x"ee", x"ee", x"f1", x"f0", x"f0", x"f1", 
        x"e2", x"6d", x"66", x"a2", x"b8", x"bf", x"d2", x"df", x"b5", x"ab", x"a6", x"a4", x"96", x"86", x"7b", 
        x"6f", x"70", x"7d", x"8b", x"98", x"99", x"9e", x"89", x"70", x"98", x"99", x"8e", x"7d", x"6d", x"65", 
        x"69", x"77", x"85", x"88", x"89", x"91", x"8d", x"82", x"88", x"98", x"94", x"93", x"a2", x"b6", x"c0", 
        x"81", x"cd", x"e8", x"ea", x"e5", x"d6", x"c2", x"b2", x"ab", x"a9", x"a8", x"aa", x"ab", x"b5", x"db", 
        x"e5", x"e1", x"e1", x"e1", x"e0", x"e0", x"e0", x"e1", x"e1", x"df", x"dd", x"dc", x"dc", x"dd", x"df", 
        x"de", x"de", x"df", x"de", x"de", x"de", x"de", x"de", x"de", x"df", x"df", x"df", x"df", x"df", x"df", 
        x"df", x"df", x"dd", x"dd", x"dd", x"dd", x"dc", x"db", x"df", x"dd", x"dc", x"de", x"e1", x"e1", x"df", 
        x"e1", x"dd", x"d1", x"c1", x"ad", x"9e", x"9d", x"9b", x"98", x"97", x"99", x"9e", x"a5", x"ab", x"b3", 
        x"b6", x"ad", x"9e", x"87", x"6a", x"48", x"2d", x"20", x"15", x"0b", x"0b", x"0c", x"12", x"11", x"0a", 
        x"0f", x"0b", x"22", x"5f", x"65", x"65", x"6f", x"73", x"79", x"81", x"85", x"84", x"82", x"7e", x"7d", 
        x"94", x"96", x"96", x"97", x"94", x"95", x"94", x"92", x"95", x"95", x"96", x"97", x"93", x"91", x"94", 
        x"95", x"96", x"96", x"95", x"95", x"97", x"94", x"91", x"96", x"95", x"93", x"94", x"95", x"96", x"96", 
        x"95", x"95", x"94", x"94", x"95", x"96", x"95", x"95", x"96", x"96", x"95", x"94", x"93", x"92", x"93", 
        x"95", x"95", x"96", x"96", x"96", x"97", x"96", x"95", x"96", x"94", x"93", x"95", x"96", x"95", x"95", 
        x"94", x"94", x"93", x"94", x"93", x"93", x"97", x"95", x"96", x"94", x"94", x"97", x"96", x"96", x"97", 
        x"98", x"97", x"96", x"96", x"95", x"97", x"96", x"98", x"97", x"98", x"98", x"96", x"96", x"96", x"96", 
        x"96", x"97", x"97", x"96", x"99", x"9b", x"97", x"97", x"9b", x"99", x"98", x"9a", x"98", x"9a", x"97", 
        x"97", x"d4", x"d7", x"d2", x"d3", x"d5", x"d8", x"d7", x"b9", x"83", x"3e", x"1a", x"14", x"1a", x"2c", 
        x"43", x"4d", x"4d", x"4c", x"4b", x"49", x"36", x"4b", x"5e", x"46", x"3c", x"3d", x"40", x"3b", x"3a", 
        x"3a", x"3a", x"3a", x"3b", x"3e", x"40", x"43", x"43", x"42", x"3f", x"42", x"42", x"43", x"45", x"46", 
        x"43", x"69", x"d5", x"dd", x"d9", x"da", x"dc", x"db", x"dc", x"d3", x"d3", x"d1", x"d1", x"d0", x"d1", 
        x"d3", x"d4", x"d5", x"d4", x"d3", x"d2", x"d1", x"d0", x"d1", x"d2", x"d0", x"d2", x"d5", x"d4", x"d2", 
        x"d4", x"d5", x"d5", x"d5", x"d4", x"d5", x"d4", x"d3", x"d2", x"d0", x"d1", x"d1", x"d1", x"d0", x"d2", 
        x"d3", x"d4", x"d3", x"d2", x"d2", x"d2", x"d3", x"d1", x"ce", x"da", x"d0", x"d3", x"d3", x"d4", x"d3", 
        x"d1", x"d8", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f1", 
        x"f0", x"ee", x"ed", x"ed", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ee", x"ed", x"eb", x"ed", x"f0", x"f0", x"f0", 
        x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ec", x"f0", x"eb", 
        x"e3", x"d8", x"c4", x"ad", x"8d", x"70", x"5d", x"50", x"4b", x"52", x"59", x"67", x"5d", x"58", x"69", 
        x"5c", x"56", x"56", x"55", x"58", x"56", x"56", x"56", x"55", x"51", x"4e", x"51", x"53", x"50", x"4f", 
        x"53", x"58", x"5b", x"60", x"5b", x"58", x"5b", x"59", x"59", x"57", x"51", x"4c", x"46", x"36", x"28", 
        x"1e", x"13", x"0c", x"0c", x"0f", x"14", x"1e", x"34", x"4e", x"64", x"74", x"82", x"85", x"7f", x"73", 
        x"6c", x"6b", x"73", x"83", x"9c", x"ba", x"d6", x"e4", x"ea", x"f1", x"f3", x"f4", x"f3", x"f3", x"f2", 
        x"f1", x"f0", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f2", x"f1", x"f2", x"ec", x"f0", x"f3", x"f3", x"f2", 
        x"f3", x"f3", x"f1", x"f2", x"f2", x"f2", x"f3", x"f5", x"f4", x"f3", x"f2", x"f4", x"f5", x"f4", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f1", x"ec", x"e3", 
        x"d1", x"c1", x"ae", x"b0", x"be", x"d1", x"e3", x"eb", x"ef", x"f2", x"f4", x"f3", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"ef", x"f2", x"f2", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f2", x"f3", x"ef", x"f2", x"f2", x"f1", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"f2", 
        x"ea", x"7b", x"9a", x"bf", x"e7", x"de", x"cd", x"ba", x"8d", x"84", x"79", x"78", x"78", x"7f", x"90", 
        x"97", x"9d", x"9b", x"97", x"9b", x"9a", x"98", x"81", x"60", x"6a", x"67", x"68", x"71", x"80", x"8f", 
        x"92", x"91", x"93", x"8d", x"7f", x"77", x"6f", x"62", x"66", x"6f", x"76", x"84", x"97", x"bf", x"d6", 
        x"96", x"bd", x"c7", x"b9", x"aa", x"a7", x"ab", x"ae", x"b1", x"b4", x"b2", x"b3", x"b1", x"b5", x"d8", 
        x"e2", x"e1", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"de", x"dd", x"dd", x"de", x"df", x"df", 
        x"de", x"de", x"df", x"df", x"de", x"de", x"de", x"de", x"de", x"e0", x"df", x"df", x"de", x"dd", x"dd", 
        x"de", x"df", x"de", x"dd", x"dd", x"df", x"df", x"de", x"e1", x"e2", x"e1", x"e0", x"da", x"ce", x"c3", 
        x"b4", x"a5", x"98", x"94", x"96", x"9e", x"a6", x"a9", x"a9", x"ab", x"ae", x"aa", x"9e", x"90", x"7c", 
        x"5d", x"3f", x"23", x"17", x"11", x"0e", x"0c", x"0e", x"17", x"21", x"2c", x"34", x"39", x"2b", x"15", 
        x"1f", x"13", x"30", x"85", x"90", x"89", x"86", x"85", x"83", x"81", x"7f", x"7d", x"7c", x"78", x"76", 
        x"96", x"96", x"95", x"94", x"94", x"94", x"94", x"93", x"94", x"95", x"96", x"96", x"95", x"94", x"96", 
        x"93", x"94", x"97", x"96", x"96", x"96", x"93", x"92", x"94", x"94", x"96", x"95", x"93", x"93", x"94", 
        x"94", x"95", x"96", x"94", x"95", x"93", x"95", x"96", x"96", x"96", x"96", x"96", x"96", x"95", x"96", 
        x"98", x"97", x"98", x"97", x"97", x"96", x"96", x"96", x"97", x"95", x"95", x"96", x"9a", x"97", x"94", 
        x"94", x"96", x"95", x"94", x"93", x"93", x"95", x"96", x"97", x"97", x"96", x"97", x"99", x"98", x"99", 
        x"99", x"97", x"97", x"9a", x"97", x"98", x"97", x"96", x"98", x"99", x"98", x"95", x"96", x"96", x"97", 
        x"98", x"98", x"99", x"97", x"98", x"99", x"96", x"96", x"98", x"98", x"97", x"98", x"98", x"97", x"95", 
        x"94", x"d3", x"d7", x"d6", x"d7", x"d8", x"c4", x"80", x"3b", x"1c", x"14", x"1b", x"2b", x"3f", x"4d", 
        x"52", x"50", x"4e", x"4b", x"4a", x"4a", x"34", x"4a", x"61", x"4c", x"43", x"3b", x"39", x"3c", x"3b", 
        x"37", x"3c", x"40", x"3e", x"41", x"43", x"42", x"42", x"41", x"3f", x"42", x"45", x"47", x"47", x"46", 
        x"42", x"63", x"d3", x"dd", x"dc", x"de", x"dc", x"dc", x"db", x"d3", x"d4", x"d3", x"d3", x"d4", x"d2", 
        x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d3", x"d2", x"d3", x"d4", x"d2", x"d3", x"d4", x"d4", x"d3", 
        x"d4", x"d5", x"d5", x"d2", x"d4", x"d6", x"d2", x"d1", x"d2", x"d0", x"cf", x"d1", x"d1", x"cf", x"d3", 
        x"d4", x"d4", x"d3", x"d1", x"d1", x"d2", x"d4", x"d0", x"cf", x"de", x"d3", x"d3", x"d4", x"d3", x"d2", 
        x"d1", x"d5", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"ef", x"f0", x"f2", x"f1", 
        x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"f1", x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ed", x"ed", x"e9", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"ee", x"e9", x"df", x"d0", x"b5", x"96", x"7a", x"60", x"49", x"5a", x"6e", x"65", 
        x"5b", x"55", x"53", x"55", x"58", x"57", x"57", x"53", x"55", x"53", x"51", x"51", x"50", x"4f", x"50", 
        x"50", x"50", x"54", x"59", x"5a", x"5c", x"5d", x"5e", x"61", x"5c", x"57", x"59", x"5c", x"5a", x"54", 
        x"4d", x"41", x"31", x"24", x"1c", x"12", x"0b", x"0b", x"0e", x"13", x"1d", x"38", x"52", x"65", x"73", 
        x"7c", x"85", x"83", x"76", x"6e", x"6c", x"78", x"89", x"9e", x"bb", x"d2", x"e2", x"ec", x"f3", x"f5", 
        x"f3", x"f1", x"f3", x"f2", x"f1", x"f4", x"f5", x"f3", x"f3", x"f4", x"f2", x"f1", x"f2", x"f2", x"f4", 
        x"f4", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f4", x"f5", x"f4", x"f2", x"f3", x"f4", x"f5", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f1", x"eb", x"ef", x"f3", x"f2", x"f2", 
        x"f4", x"f3", x"f0", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", 
        x"f2", x"f0", x"e7", x"d8", x"c2", x"b0", x"ab", x"b9", x"ca", x"dd", x"e7", x"ed", x"f2", x"f3", x"f4", 
        x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f2", x"f3", x"f2", x"f2", 
        x"f2", x"f1", x"f2", x"f2", x"f3", x"f5", x"f4", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ed", x"ef", x"f3", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"ef", x"f0", x"ee", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f1", x"f0", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f3", x"f1", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f3", x"f4", x"f3", x"f2", x"f1", x"f0", x"ef", x"f1", x"f1", x"f1", 
        x"ea", x"87", x"9a", x"b9", x"c1", x"c6", x"af", x"a1", x"95", x"7b", x"6b", x"81", x"94", x"9b", x"a0", 
        x"a1", x"9e", x"99", x"8e", x"85", x"74", x"6b", x"58", x"47", x"75", x"8f", x"93", x"91", x"90", x"8e", 
        x"86", x"7f", x"76", x"65", x"5f", x"67", x"77", x"7f", x"80", x"7b", x"75", x"75", x"86", x"a5", x"b5", 
        x"b5", x"b4", x"ae", x"b4", x"b2", x"b2", x"b4", x"b5", x"b6", x"b4", x"b2", x"b5", x"b3", x"b3", x"d5", 
        x"e3", x"e1", x"e0", x"e1", x"e0", x"e0", x"e1", x"df", x"de", x"e0", x"df", x"df", x"df", x"e0", x"e0", 
        x"df", x"df", x"de", x"de", x"de", x"de", x"df", x"e0", x"e0", x"dd", x"dd", x"df", x"df", x"dc", x"dc", 
        x"dd", x"dc", x"e0", x"e1", x"df", x"e1", x"e4", x"df", x"da", x"d4", x"c0", x"b3", x"a4", x"97", x"95", 
        x"9a", x"a2", x"a4", x"a8", x"aa", x"af", x"b0", x"aa", x"9c", x"8b", x"79", x"5b", x"39", x"21", x"14", 
        x"10", x"0e", x"0b", x"0e", x"17", x"24", x"2f", x"36", x"3d", x"41", x"49", x"53", x"61", x"51", x"25", 
        x"27", x"17", x"33", x"89", x"93", x"8a", x"85", x"84", x"81", x"7f", x"7d", x"72", x"69", x"65", x"6c", 
        x"96", x"96", x"94", x"94", x"93", x"93", x"94", x"94", x"94", x"96", x"96", x"97", x"96", x"95", x"96", 
        x"94", x"94", x"97", x"96", x"96", x"96", x"95", x"95", x"94", x"92", x"95", x"95", x"96", x"96", x"93", 
        x"94", x"95", x"97", x"95", x"95", x"94", x"94", x"95", x"95", x"95", x"95", x"96", x"96", x"97", x"95", 
        x"96", x"96", x"99", x"97", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"93", x"91", 
        x"94", x"96", x"96", x"95", x"94", x"93", x"95", x"97", x"98", x"97", x"97", x"96", x"98", x"98", x"98", 
        x"98", x"96", x"97", x"9a", x"98", x"99", x"99", x"97", x"98", x"98", x"96", x"96", x"97", x"97", x"98", 
        x"98", x"99", x"9a", x"99", x"9a", x"9a", x"98", x"97", x"98", x"98", x"99", x"9a", x"98", x"98", x"92", 
        x"96", x"d5", x"d8", x"d9", x"c1", x"8c", x"48", x"1a", x"12", x"1e", x"2f", x"42", x"4e", x"50", x"51", 
        x"50", x"4b", x"48", x"48", x"4b", x"48", x"34", x"49", x"5e", x"49", x"45", x"3f", x"38", x"3a", x"3d", 
        x"3b", x"3f", x"42", x"42", x"43", x"44", x"41", x"3f", x"40", x"42", x"45", x"47", x"48", x"47", x"46", 
        x"3f", x"5a", x"cc", x"d7", x"d7", x"d9", x"d7", x"d9", x"dd", x"d3", x"d3", x"d0", x"d1", x"d3", x"d1", 
        x"d3", x"d4", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d4", x"d4", x"d3", x"d3", x"d4", x"d4", x"d3", 
        x"d4", x"d5", x"d5", x"d2", x"d4", x"d7", x"d2", x"d2", x"d3", x"d2", x"d0", x"d2", x"d2", x"d0", x"d3", 
        x"d5", x"d4", x"d3", x"d1", x"d1", x"d2", x"d4", x"d0", x"cf", x"de", x"d2", x"d2", x"d3", x"d2", x"d2", 
        x"d1", x"d6", x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", 
        x"ef", x"ef", x"f0", x"f0", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"ee", x"ee", x"e9", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"f0", x"ee", x"f0", x"f4", x"f1", x"eb", x"e8", x"da", x"bb", x"a0", x"84", x"68", 
        x"5f", x"51", x"4b", x"4c", x"4c", x"4c", x"52", x"54", x"50", x"52", x"54", x"52", x"50", x"51", x"4f", 
        x"4e", x"4e", x"50", x"52", x"51", x"55", x"58", x"58", x"5d", x"5d", x"59", x"5a", x"5e", x"5d", x"58", 
        x"5a", x"59", x"57", x"52", x"4c", x"40", x"34", x"28", x"1e", x"17", x"11", x"0b", x"0b", x"0f", x"19", 
        x"30", x"51", x"67", x"74", x"7e", x"88", x"83", x"7a", x"6c", x"67", x"6f", x"87", x"a4", x"bc", x"d0", 
        x"e1", x"ea", x"ee", x"f0", x"f2", x"f5", x"f5", x"f3", x"f1", x"f1", x"f5", x"f5", x"f4", x"f2", x"f1", 
        x"f2", x"f3", x"f2", x"f2", x"f3", x"f2", x"f1", x"f3", x"f7", x"f6", x"f3", x"f2", x"f4", x"f4", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f1", x"ec", x"ee", x"f3", x"f3", x"f2", 
        x"f4", x"f3", x"f1", x"f2", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"f2", x"f3", x"f3", x"f3", 
        x"f4", x"f5", x"f2", x"f3", x"f2", x"ec", x"dd", x"c8", x"b8", x"ae", x"b1", x"be", x"d0", x"e0", x"eb", 
        x"f2", x"f5", x"f5", x"f4", x"f1", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f3", 
        x"f3", x"f2", x"f4", x"f2", x"f1", x"f2", x"f3", x"f3", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"ef", x"f1", x"f4", x"f3", x"f3", x"f2", x"f1", 
        x"f2", x"f2", x"ef", x"f0", x"ed", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f3", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f1", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f0", x"f3", 
        x"ee", x"8b", x"70", x"97", x"8e", x"ad", x"c8", x"da", x"dc", x"b3", x"98", x"92", x"7c", x"73", x"7f", 
        x"86", x"75", x"6a", x"66", x"6c", x"7a", x"8f", x"88", x"64", x"86", x"91", x"8a", x"81", x"77", x"6c", 
        x"65", x"6c", x"73", x"7b", x"7d", x"7b", x"79", x"7e", x"91", x"ac", x"c4", x"d3", x"de", x"db", x"c1", 
        x"b7", x"b8", x"b9", x"b9", x"b9", x"b8", x"b7", x"b7", x"b7", x"b6", x"b5", x"b5", x"b5", x"b5", x"d3", 
        x"e4", x"e1", x"e1", x"e2", x"df", x"de", x"e0", x"de", x"e0", x"e0", x"df", x"e0", x"e0", x"e0", x"e0", 
        x"df", x"e0", x"e0", x"df", x"df", x"df", x"de", x"de", x"de", x"dd", x"df", x"df", x"de", x"df", x"df", 
        x"e0", x"e3", x"e3", x"e0", x"d7", x"cc", x"c1", x"b3", x"a8", x"9d", x"92", x"98", x"a1", x"a7", x"a8", 
        x"aa", x"ad", x"ac", x"a9", x"9f", x"89", x"71", x"52", x"32", x"1b", x"0f", x"0b", x"0b", x"11", x"16", 
        x"1c", x"24", x"2d", x"36", x"41", x"4b", x"51", x"56", x"62", x"6f", x"7a", x"82", x"85", x"68", x"25", 
        x"29", x"1e", x"2e", x"83", x"92", x"84", x"80", x"79", x"71", x"72", x"79", x"81", x"8f", x"ad", x"c4", 
        x"9a", x"9a", x"99", x"98", x"97", x"97", x"97", x"95", x"95", x"96", x"96", x"96", x"95", x"95", x"96", 
        x"94", x"95", x"97", x"96", x"96", x"96", x"96", x"96", x"94", x"93", x"95", x"97", x"97", x"97", x"93", 
        x"93", x"94", x"95", x"94", x"94", x"93", x"96", x"96", x"96", x"96", x"96", x"95", x"96", x"98", x"95", 
        x"95", x"95", x"98", x"97", x"96", x"95", x"96", x"96", x"95", x"97", x"97", x"96", x"97", x"96", x"94", 
        x"97", x"98", x"96", x"93", x"94", x"95", x"96", x"98", x"98", x"98", x"97", x"97", x"97", x"97", x"97", 
        x"97", x"95", x"97", x"98", x"97", x"98", x"99", x"98", x"98", x"98", x"97", x"98", x"99", x"98", x"98", 
        x"98", x"98", x"98", x"99", x"9b", x"9b", x"99", x"99", x"99", x"98", x"98", x"9b", x"9c", x"99", x"92", 
        x"9c", x"c8", x"ae", x"7f", x"3c", x"18", x"10", x"21", x"31", x"42", x"52", x"54", x"50", x"4b", x"4b", 
        x"4b", x"4a", x"4a", x"49", x"49", x"42", x"33", x"4a", x"5f", x"48", x"49", x"45", x"3c", x"3d", x"42", 
        x"42", x"44", x"44", x"41", x"41", x"43", x"44", x"46", x"46", x"45", x"46", x"47", x"47", x"46", x"46", 
        x"40", x"5c", x"cf", x"dd", x"d9", x"da", x"d8", x"db", x"dd", x"d1", x"cf", x"cd", x"d0", x"d2", x"d2", 
        x"d4", x"d5", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d4", x"d4", x"d3", x"d3", x"d4", x"d4", x"d3", 
        x"d4", x"d5", x"d5", x"d2", x"d4", x"d7", x"d3", x"d4", x"d4", x"d3", x"d2", x"d2", x"d2", x"d1", x"d3", 
        x"d4", x"d3", x"d3", x"d2", x"d1", x"d2", x"d3", x"d0", x"cf", x"dc", x"d2", x"d1", x"d2", x"d2", x"d2", 
        x"d2", x"d6", x"f0", x"ef", x"ef", x"f1", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"ee", x"f0", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"f0", x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ed", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ea", x"f0", x"ef", 
        x"f1", x"f0", x"ef", x"f1", x"f0", x"ed", x"f0", x"f0", x"ef", x"f1", x"ef", x"f3", x"f5", x"f1", x"e3", 
        x"d1", x"b4", x"95", x"77", x"60", x"52", x"4d", x"48", x"42", x"46", x"4c", x"51", x"53", x"53", x"52", 
        x"52", x"53", x"56", x"56", x"51", x"51", x"53", x"53", x"53", x"53", x"52", x"54", x"57", x"56", x"53", 
        x"54", x"54", x"52", x"54", x"57", x"57", x"56", x"56", x"4d", x"43", x"39", x"2d", x"20", x"16", x"0c", 
        x"08", x"07", x"09", x"1a", x"32", x"49", x"58", x"6a", x"7c", x"86", x"84", x"7a", x"6b", x"67", x"6e", 
        x"85", x"99", x"b1", x"ca", x"dd", x"ea", x"f5", x"f7", x"f5", x"f4", x"f5", x"f3", x"f0", x"f5", x"f3", 
        x"f3", x"f5", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f4", x"f4", x"f4", x"f3", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f4", x"f1", x"ed", x"ee", x"f3", x"f3", x"f2", 
        x"f4", x"f3", x"f1", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f2", x"f3", x"f1", x"f1", x"f2", x"f4", x"f6", x"f5", x"eb", x"d6", x"bf", x"af", x"ab", x"b6", 
        x"c5", x"d4", x"de", x"e9", x"f3", x"f7", x"f6", x"f3", x"ef", x"f0", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f2", x"f5", x"f3", x"f0", x"f0", x"f2", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f4", x"f3", x"f3", x"f2", x"f1", 
        x"f2", x"f2", x"ef", x"f0", x"ed", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"ee", x"f1", 
        x"ef", x"8e", x"74", x"c9", x"c9", x"d6", x"f3", x"ed", x"e3", x"bc", x"8e", x"87", x"81", x"67", x"5a", 
        x"5d", x"5d", x"76", x"8b", x"96", x"97", x"94", x"81", x"59", x"6b", x"6f", x"63", x"65", x"6e", x"79", 
        x"7f", x"84", x"85", x"7f", x"8c", x"a9", x"c6", x"d8", x"e1", x"e6", x"e2", x"de", x"e0", x"dc", x"c4", 
        x"ba", x"bd", x"bc", x"ba", x"b9", x"b7", x"b6", x"b6", x"b6", x"b6", x"b5", x"b4", x"b4", x"b1", x"d2", 
        x"e7", x"e0", x"e1", x"e2", x"de", x"dc", x"de", x"de", x"e1", x"de", x"dd", x"de", x"df", x"df", x"df", 
        x"df", x"e0", x"df", x"de", x"de", x"df", x"de", x"df", x"e0", x"e3", x"e3", x"e2", x"e2", x"e3", x"dd", 
        x"d3", x"c8", x"be", x"b2", x"a4", x"9b", x"99", x"99", x"a2", x"a7", x"b1", x"b0", x"b0", x"ab", x"a1", 
        x"93", x"83", x"67", x"4b", x"2c", x"11", x"09", x"09", x"0b", x"12", x"1a", x"20", x"24", x"2e", x"3c", 
        x"4a", x"55", x"5a", x"5e", x"67", x"72", x"7d", x"88", x"85", x"7c", x"7a", x"7b", x"7c", x"62", x"25", 
        x"24", x"1b", x"26", x"70", x"86", x"7f", x"84", x"91", x"a5", x"bd", x"d5", x"e3", x"ed", x"ee", x"ea", 
        x"9a", x"9a", x"99", x"98", x"98", x"97", x"97", x"97", x"96", x"96", x"96", x"96", x"95", x"95", x"95", 
        x"95", x"96", x"96", x"95", x"96", x"96", x"95", x"96", x"96", x"95", x"97", x"98", x"96", x"97", x"95", 
        x"95", x"95", x"95", x"94", x"94", x"94", x"97", x"97", x"97", x"97", x"96", x"95", x"95", x"98", x"96", 
        x"96", x"95", x"97", x"95", x"96", x"96", x"97", x"96", x"95", x"97", x"98", x"97", x"97", x"97", x"96", 
        x"98", x"98", x"97", x"96", x"97", x"96", x"96", x"97", x"97", x"97", x"98", x"97", x"97", x"97", x"97", 
        x"96", x"96", x"97", x"98", x"97", x"97", x"97", x"98", x"99", x"99", x"99", x"99", x"99", x"98", x"98", 
        x"97", x"97", x"96", x"98", x"99", x"99", x"99", x"99", x"99", x"98", x"97", x"99", x"9a", x"9a", x"9b", 
        x"9c", x"9b", x"61", x"1f", x"15", x"20", x"2f", x"44", x"51", x"53", x"50", x"4c", x"4c", x"4f", x"4e", 
        x"4a", x"4a", x"49", x"42", x"42", x"3e", x"32", x"48", x"5c", x"4a", x"48", x"46", x"41", x"43", x"43", 
        x"43", x"46", x"46", x"44", x"44", x"45", x"47", x"48", x"48", x"47", x"47", x"47", x"45", x"45", x"46", 
        x"40", x"5a", x"cd", x"de", x"d8", x"d8", x"d7", x"da", x"dd", x"d0", x"cf", x"cf", x"d1", x"d3", x"d4", 
        x"d3", x"d4", x"d3", x"d3", x"d3", x"d2", x"d2", x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", 
        x"d4", x"d5", x"d5", x"d2", x"d4", x"d7", x"d3", x"d4", x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", 
        x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d0", x"cf", x"dc", x"d2", x"d2", x"d2", x"d2", x"d3", 
        x"d2", x"d7", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"ef", 
        x"f1", x"f2", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"f1", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ed", x"ee", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"ea", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"f1", x"ef", x"ef", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"ef", x"ef", x"f2", 
        x"f3", x"f0", x"ea", x"e2", x"d1", x"b6", x"9d", x"88", x"73", x"5f", x"51", x"48", x"44", x"45", x"49", 
        x"52", x"55", x"58", x"5a", x"56", x"53", x"54", x"54", x"53", x"53", x"56", x"56", x"52", x"51", x"51", 
        x"52", x"52", x"52", x"53", x"52", x"51", x"4e", x"4d", x"52", x"58", x"5c", x"5e", x"55", x"46", x"36", 
        x"2d", x"25", x"1b", x"13", x"0c", x"0b", x"0f", x"1c", x"2e", x"43", x"56", x"6a", x"7a", x"80", x"82", 
        x"7d", x"73", x"71", x"7b", x"89", x"99", x"af", x"c4", x"da", x"e9", x"f1", x"f5", x"f5", x"f4", x"f3", 
        x"f3", x"f4", x"f5", x"f5", x"f4", x"f1", x"f2", x"f4", x"f3", x"f2", x"f2", x"f4", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f2", x"ee", x"ed", x"f3", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f3", x"f4", x"f6", x"f5", x"f1", x"e9", x"d9", x"c8", 
        x"ba", x"b3", x"b5", x"be", x"ca", x"d9", x"e6", x"f0", x"f3", x"f4", x"f2", x"ef", x"f0", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f2", x"f1", x"f2", x"f2", x"f0", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"ef", x"f0", x"ed", x"f2", x"f2", x"f3", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", 
        x"f2", x"f3", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"ef", 
        x"ee", x"98", x"8a", x"d7", x"c4", x"b3", x"c0", x"b7", x"b0", x"a5", x"7e", x"73", x"7d", x"8b", x"97", 
        x"9d", x"93", x"82", x"6a", x"67", x"6e", x"6a", x"5c", x"3c", x"61", x"79", x"78", x"80", x"89", x"91", 
        x"9e", x"b0", x"c3", x"d2", x"dd", x"e5", x"e4", x"e0", x"df", x"df", x"df", x"dd", x"de", x"de", x"c8", 
        x"b9", x"b9", x"b7", x"b7", x"b6", x"b5", x"b5", x"b6", x"b7", x"b7", x"b2", x"b5", x"b1", x"ac", x"d0", 
        x"e6", x"df", x"e0", x"e2", x"de", x"dd", x"df", x"de", x"e0", x"dd", x"dc", x"df", x"e1", x"e1", x"df", 
        x"dd", x"de", x"df", x"de", x"de", x"e0", x"e1", x"e1", x"e2", x"e2", x"d9", x"ce", x"c5", x"bd", x"b2", 
        x"a6", x"9e", x"9d", x"9e", x"a2", x"aa", x"b2", x"b2", x"b1", x"a7", x"9f", x"8b", x"77", x"5c", x"43", 
        x"30", x"1d", x"0d", x"0b", x"0d", x"13", x"1d", x"27", x"2c", x"31", x"3d", x"4b", x"53", x"5a", x"5f", 
        x"68", x"78", x"83", x"84", x"82", x"7f", x"7b", x"7e", x"7f", x"79", x"75", x"72", x"6b", x"57", x"32", 
        x"3f", x"50", x"68", x"9c", x"b4", x"bf", x"d0", x"e0", x"e8", x"e8", x"e7", x"e8", x"e6", x"e6", x"e6", 
        x"99", x"99", x"98", x"98", x"97", x"96", x"96", x"96", x"96", x"96", x"95", x"94", x"94", x"95", x"94", 
        x"96", x"97", x"95", x"96", x"96", x"97", x"96", x"95", x"95", x"95", x"97", x"96", x"95", x"97", x"96", 
        x"96", x"96", x"95", x"95", x"93", x"93", x"94", x"95", x"96", x"97", x"97", x"96", x"96", x"97", x"97", 
        x"99", x"96", x"95", x"94", x"97", x"97", x"98", x"97", x"95", x"97", x"99", x"97", x"97", x"97", x"95", 
        x"96", x"97", x"96", x"96", x"98", x"97", x"96", x"96", x"96", x"96", x"97", x"98", x"98", x"99", x"99", 
        x"97", x"97", x"98", x"99", x"9a", x"98", x"97", x"98", x"98", x"98", x"9a", x"99", x"99", x"98", x"98", 
        x"97", x"96", x"96", x"97", x"98", x"97", x"98", x"99", x"98", x"98", x"99", x"9a", x"9a", x"98", x"9b", 
        x"9a", x"99", x"6c", x"24", x"25", x"2f", x"3c", x"44", x"50", x"53", x"51", x"50", x"50", x"50", x"4e", 
        x"4c", x"4c", x"49", x"40", x"3e", x"3e", x"32", x"44", x"57", x"48", x"46", x"43", x"44", x"47", x"43", 
        x"41", x"44", x"46", x"46", x"46", x"48", x"4a", x"4a", x"48", x"47", x"47", x"47", x"46", x"46", x"47", 
        x"41", x"59", x"cc", x"df", x"d7", x"d8", x"d8", x"db", x"df", x"d1", x"d0", x"d1", x"d3", x"d3", x"d3", 
        x"d2", x"d2", x"d2", x"d3", x"d4", x"d3", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d4", 
        x"d4", x"d5", x"d5", x"d2", x"d4", x"d7", x"d3", x"d3", x"d2", x"d2", x"d3", x"d1", x"d1", x"d2", x"d3", 
        x"d3", x"d2", x"d2", x"d3", x"d3", x"d2", x"d2", x"d1", x"d0", x"db", x"d2", x"d3", x"d3", x"d2", x"d3", 
        x"d2", x"d6", x"f0", x"ef", x"f0", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"ee", x"ef", 
        x"f1", x"f2", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"eb", x"f0", x"ef", 
        x"ef", x"ef", x"f3", x"f1", x"ee", x"ef", x"f1", x"f1", x"f0", x"f0", x"f3", x"f0", x"f1", x"f2", x"ef", 
        x"f1", x"f1", x"ee", x"f2", x"f5", x"f4", x"f3", x"eb", x"db", x"c5", x"ac", x"92", x"78", x"61", x"4f", 
        x"44", x"3f", x"42", x"4d", x"51", x"53", x"58", x"58", x"56", x"56", x"59", x"5a", x"59", x"56", x"53", 
        x"51", x"51", x"52", x"55", x"51", x"50", x"4d", x"4f", x"50", x"52", x"56", x"5d", x"64", x"68", x"5f", 
        x"58", x"52", x"49", x"3b", x"28", x"1d", x"15", x"0d", x"04", x"04", x"0b", x"1a", x"2e", x"43", x"57", 
        x"6e", x"7e", x"86", x"82", x"78", x"71", x"6a", x"74", x"83", x"93", x"ab", x"c7", x"e0", x"f0", x"f4", 
        x"f5", x"f5", x"f5", x"f4", x"f1", x"f3", x"f4", x"f3", x"f2", x"f3", x"f4", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"ef", x"ed", x"f2", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f4", x"f4", x"f3", x"f2", 
        x"f3", x"f4", x"f2", x"f1", x"f2", x"f4", x"f5", x"f4", x"f2", x"f2", x"f3", x"f3", x"f3", x"f6", x"f7", 
        x"f3", x"e0", x"d0", x"c1", x"b3", x"b0", x"b6", x"c0", x"d3", x"e5", x"f1", x"f4", x"f4", x"f3", x"f3", 
        x"f4", x"f4", x"f2", x"f0", x"f0", x"f3", x"f3", x"f0", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"ef", x"f1", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"ef", x"f0", x"ed", x"f2", x"f2", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", 
        x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"ef", 
        x"ef", x"99", x"6a", x"a5", x"9a", x"8e", x"90", x"ad", x"bd", x"d3", x"c4", x"9d", x"a0", x"9a", x"89", 
        x"7c", x"75", x"76", x"6d", x"65", x"65", x"5d", x"58", x"4b", x"7a", x"97", x"a1", x"b2", x"c5", x"d6", 
        x"e1", x"e4", x"e5", x"e4", x"e3", x"e1", x"df", x"df", x"e2", x"e1", x"e0", x"df", x"dd", x"de", x"c9", 
        x"b9", x"bb", x"ba", x"bb", x"b9", x"b7", x"b6", x"b6", x"b6", x"b6", x"b6", x"b7", x"b1", x"a9", x"cc", 
        x"e5", x"e4", x"e0", x"e1", x"df", x"de", x"e0", x"de", x"df", x"e0", x"df", x"df", x"e0", x"e0", x"e0", 
        x"df", x"e0", x"e2", x"e5", x"e6", x"e4", x"da", x"cf", x"c6", x"bd", x"b2", x"a7", x"9f", x"9e", x"9f", 
        x"a2", x"aa", x"b1", x"b7", x"b3", x"ac", x"a2", x"8d", x"72", x"5a", x"41", x"28", x"13", x"06", x"03", 
        x"0d", x"13", x"1b", x"1f", x"23", x"30", x"3e", x"4b", x"54", x"5b", x"65", x"6f", x"79", x"7f", x"81", 
        x"81", x"81", x"7f", x"7c", x"7b", x"7a", x"77", x"71", x"6d", x"62", x"61", x"69", x"78", x"83", x"8f", 
        x"ae", x"c9", x"db", x"e5", x"e7", x"ec", x"e9", x"e8", x"e7", x"e4", x"e3", x"e6", x"e5", x"e5", x"e7", 
        x"99", x"99", x"9a", x"9a", x"98", x"98", x"97", x"98", x"98", x"96", x"95", x"94", x"94", x"95", x"94", 
        x"97", x"97", x"95", x"95", x"96", x"96", x"97", x"98", x"97", x"94", x"96", x"95", x"94", x"96", x"96", 
        x"96", x"96", x"95", x"96", x"95", x"96", x"95", x"96", x"98", x"9a", x"9a", x"99", x"99", x"98", x"98", 
        x"99", x"97", x"97", x"95", x"96", x"95", x"98", x"99", x"95", x"96", x"99", x"98", x"95", x"93", x"93", 
        x"96", x"97", x"97", x"98", x"99", x"96", x"96", x"97", x"96", x"96", x"95", x"96", x"98", x"9b", x"99", 
        x"97", x"98", x"99", x"99", x"9a", x"99", x"98", x"99", x"98", x"97", x"99", x"99", x"99", x"99", x"99", 
        x"98", x"98", x"98", x"99", x"99", x"98", x"9a", x"9a", x"98", x"98", x"99", x"99", x"97", x"9a", x"9a", 
        x"9a", x"9a", x"8a", x"6a", x"6f", x"63", x"5e", x"4f", x"48", x"40", x"3d", x"40", x"45", x"4c", x"52", 
        x"53", x"50", x"4e", x"4b", x"44", x"42", x"31", x"43", x"5a", x"48", x"44", x"44", x"44", x"47", x"46", 
        x"43", x"47", x"4c", x"4a", x"46", x"47", x"4a", x"4a", x"47", x"47", x"48", x"49", x"49", x"4a", x"4a", 
        x"45", x"5f", x"cf", x"e1", x"d7", x"d7", x"d6", x"d9", x"e0", x"d1", x"cf", x"d1", x"d3", x"d3", x"d2", 
        x"d2", x"d2", x"d3", x"d4", x"d3", x"d3", x"d2", x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d4", 
        x"d4", x"d5", x"d5", x"d2", x"d4", x"d7", x"d3", x"d3", x"d1", x"d2", x"d3", x"d1", x"d1", x"d3", x"d3", 
        x"d2", x"d1", x"d3", x"d4", x"d4", x"d2", x"d2", x"d2", x"d1", x"dc", x"d2", x"d4", x"d3", x"d2", x"d2", 
        x"d1", x"d6", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"f0", x"ef", 
        x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", 
        x"f1", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"ea", x"f0", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ee", x"f0", x"f3", x"f0", x"ee", x"ef", x"ef", 
        x"f1", x"f1", x"ef", x"f1", x"f1", x"ef", x"f2", x"f3", x"f3", x"f5", x"f5", x"f0", x"e7", x"d6", x"c3", 
        x"ab", x"8f", x"73", x"58", x"45", x"40", x"3f", x"42", x"4d", x"56", x"5b", x"58", x"55", x"54", x"56", 
        x"5a", x"55", x"52", x"56", x"53", x"55", x"54", x"55", x"54", x"54", x"54", x"52", x"54", x"5b", x"62", 
        x"62", x"5d", x"54", x"50", x"4a", x"49", x"4a", x"46", x"37", x"21", x"13", x"0f", x"07", x"08", x"0c", 
        x"15", x"22", x"34", x"4a", x"64", x"77", x"7f", x"83", x"81", x"7a", x"73", x"73", x"79", x"88", x"a0", 
        x"bc", x"d8", x"e9", x"f2", x"f4", x"f4", x"f5", x"f4", x"f2", x"f3", x"f4", x"f1", x"f0", x"f1", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f0", x"ed", x"f3", x"f4", x"f2", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f4", x"f4", x"f3", x"f3", 
        x"f4", x"f5", x"f3", x"f4", x"f3", x"f2", x"f2", x"f3", x"f4", x"f3", x"f4", x"f4", x"f0", x"ee", x"f0", 
        x"f2", x"f4", x"f2", x"f0", x"eb", x"df", x"d1", x"c1", x"b4", x"ad", x"ad", x"bc", x"d5", x"eb", x"f5", 
        x"f3", x"f1", x"f3", x"f2", x"f1", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"ee", x"f1", x"f2", x"f0", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"ef", x"f0", x"ed", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"f2", x"f2", x"f2", x"f4", 
        x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ec", x"ef", 
        x"f1", x"a3", x"55", x"aa", x"be", x"ba", x"b9", x"e2", x"e8", x"da", x"be", x"7f", x"6b", x"6a", x"75", 
        x"79", x"79", x"74", x"71", x"78", x"8e", x"9f", x"b0", x"bd", x"ce", x"dc", x"e0", x"e5", x"e5", x"e3", 
        x"e1", x"de", x"de", x"df", x"df", x"e0", x"df", x"de", x"de", x"e0", x"e0", x"de", x"dd", x"e0", x"cc", 
        x"b8", x"bb", x"ba", x"b9", x"b8", x"b8", x"b7", x"b7", x"b8", x"b6", x"b0", x"af", x"ae", x"a0", x"c2", 
        x"e5", x"e2", x"df", x"e1", x"df", x"df", x"e0", x"de", x"de", x"e0", x"dd", x"dd", x"df", x"e4", x"e7", 
        x"e8", x"e5", x"dc", x"cd", x"bf", x"b4", x"ab", x"a4", x"a3", x"a5", x"a7", x"a8", x"ae", x"b7", x"bc", 
        x"b9", x"ad", x"99", x"7c", x"58", x"40", x"31", x"21", x"15", x"1b", x"11", x"09", x"0a", x"1f", x"30", 
        x"32", x"30", x"3e", x"4a", x"54", x"66", x"6f", x"76", x"7a", x"7c", x"7d", x"7d", x"7c", x"78", x"79", 
        x"7c", x"79", x"76", x"6d", x"63", x"5d", x"60", x"6f", x"83", x"9a", x"b1", x"c6", x"d6", x"e2", x"e8", 
        x"ef", x"ec", x"eb", x"e6", x"e4", x"e8", x"e7", x"e4", x"e6", x"e8", x"eb", x"ef", x"ee", x"e7", x"d9", 
        x"97", x"98", x"98", x"98", x"97", x"96", x"95", x"98", x"99", x"97", x"96", x"96", x"96", x"96", x"94", 
        x"97", x"98", x"94", x"95", x"96", x"96", x"98", x"99", x"98", x"96", x"98", x"96", x"94", x"95", x"94", 
        x"95", x"96", x"95", x"97", x"96", x"98", x"96", x"97", x"98", x"98", x"98", x"96", x"96", x"99", x"97", 
        x"97", x"97", x"99", x"97", x"95", x"94", x"98", x"99", x"96", x"95", x"98", x"98", x"97", x"96", x"96", 
        x"99", x"99", x"97", x"98", x"98", x"96", x"97", x"98", x"98", x"97", x"95", x"94", x"98", x"9a", x"99", 
        x"96", x"97", x"99", x"98", x"98", x"97", x"98", x"9a", x"99", x"98", x"9a", x"9a", x"9a", x"9a", x"9a", 
        x"9a", x"9a", x"9a", x"9b", x"9b", x"9a", x"9b", x"9b", x"98", x"98", x"99", x"97", x"98", x"9c", x"9a", 
        x"9e", x"99", x"8c", x"84", x"89", x"7e", x"89", x"85", x"7e", x"73", x"68", x"5e", x"57", x"50", x"46", 
        x"41", x"41", x"44", x"4a", x"48", x"45", x"32", x"44", x"5e", x"47", x"48", x"48", x"44", x"47", x"4a", 
        x"49", x"48", x"49", x"4a", x"49", x"4a", x"4c", x"4a", x"48", x"48", x"49", x"4a", x"4b", x"4c", x"4c", 
        x"46", x"5e", x"cf", x"e1", x"d6", x"d7", x"d7", x"da", x"df", x"cf", x"ce", x"d0", x"d2", x"d3", x"d4", 
        x"d3", x"d3", x"d4", x"d4", x"d3", x"d2", x"d1", x"d2", x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d4", 
        x"d4", x"d5", x"d5", x"d2", x"d4", x"d6", x"d4", x"d4", x"d2", x"d3", x"d4", x"d2", x"d1", x"d3", x"d3", 
        x"d1", x"d1", x"d3", x"d4", x"d4", x"d2", x"d2", x"d2", x"d2", x"dc", x"d2", x"d5", x"d4", x"d2", x"d2", 
        x"d1", x"d5", x"ee", x"ee", x"ef", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"ef", x"ee", x"ee", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"e9", x"f0", x"ef", 
        x"f1", x"f0", x"ef", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"ee", x"f0", x"f0", x"ee", x"ef", x"f0", 
        x"ef", x"f1", x"f0", x"f3", x"f1", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"ee", x"e4", x"d9", x"c6", x"b0", x"99", x"7d", x"62", x"51", x"46", x"44", x"4a", x"4f", x"53", x"55", 
        x"57", x"54", x"54", x"5a", x"56", x"57", x"54", x"51", x"51", x"51", x"52", x"52", x"4f", x"49", x"51", 
        x"55", x"5a", x"66", x"77", x"6f", x"5a", x"58", x"60", x"5c", x"53", x"57", x"59", x"38", x"22", x"1a", 
        x"0d", x"09", x"0b", x"10", x"19", x"24", x"31", x"49", x"61", x"73", x"7d", x"80", x"7e", x"77", x"74", 
        x"75", x"7c", x"8e", x"a5", x"bb", x"d2", x"e2", x"ee", x"f1", x"f3", x"f4", x"f3", x"f1", x"f2", x"f3", 
        x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f4", x"f3", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f0", x"ec", x"f3", x"f4", x"f2", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", 
        x"f3", x"f4", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f4", x"f3", x"f1", x"f0", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"ef", x"ed", x"e4", x"d8", x"cb", x"bc", x"b2", x"b3", x"be", 
        x"cf", x"e2", x"ed", x"f2", x"f3", x"f2", x"f3", x"f3", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"ee", x"f2", x"f3", x"f1", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"ef", x"f0", x"ee", x"f2", x"f1", x"f1", x"f1", x"f1", x"f3", x"f2", x"f1", x"f1", x"f5", 
        x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ef", x"f0", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ef", x"b1", x"70", x"cc", x"d4", x"c0", x"a9", x"a4", x"ad", x"a7", x"ae", x"a7", x"80", x"75", x"7c", 
        x"81", x"90", x"a1", x"af", x"c0", x"d1", x"da", x"e2", x"e5", x"e5", x"e4", x"e1", x"e2", x"e0", x"df", 
        x"e0", x"df", x"df", x"e1", x"df", x"dd", x"df", x"e0", x"de", x"df", x"e0", x"dd", x"dc", x"e1", x"ce", 
        x"b9", x"ba", x"b8", x"b8", x"b8", x"b6", x"b4", x"b1", x"ae", x"aa", x"a0", x"95", x"87", x"6d", x"a1", 
        x"e3", x"e4", x"e0", x"e0", x"de", x"de", x"e0", x"df", x"e0", x"e2", x"e3", x"e0", x"df", x"d9", x"cd", 
        x"bf", x"b5", x"ae", x"a8", x"a6", x"a8", x"ab", x"ac", x"af", x"b7", x"b6", x"b0", x"a7", x"98", x"7d", 
        x"5e", x"43", x"36", x"29", x"25", x"30", x"42", x"4b", x"42", x"49", x"23", x"09", x"18", x"4c", x"62", 
        x"61", x"58", x"6a", x"7b", x"7d", x"7d", x"7e", x"7e", x"7d", x"7a", x"77", x"76", x"75", x"72", x"6d", 
        x"66", x"62", x"69", x"7a", x"8c", x"a1", x"b4", x"c6", x"d4", x"df", x"e7", x"ec", x"e7", x"e8", x"e7", 
        x"e9", x"e5", x"e5", x"e8", x"e6", x"e8", x"e9", x"e8", x"e6", x"dd", x"cd", x"b7", x"9a", x"77", x"57", 
        x"98", x"99", x"9b", x"9a", x"98", x"95", x"94", x"98", x"98", x"97", x"97", x"98", x"98", x"97", x"95", 
        x"95", x"97", x"96", x"96", x"95", x"95", x"97", x"99", x"9a", x"99", x"98", x"96", x"96", x"97", x"98", 
        x"97", x"98", x"98", x"97", x"95", x"96", x"95", x"98", x"98", x"95", x"96", x"98", x"98", x"98", x"97", 
        x"95", x"95", x"96", x"97", x"97", x"96", x"97", x"97", x"96", x"96", x"97", x"98", x"98", x"98", x"97", 
        x"95", x"95", x"97", x"98", x"98", x"99", x"9a", x"99", x"98", x"99", x"98", x"96", x"99", x"9a", x"99", 
        x"98", x"99", x"99", x"99", x"99", x"98", x"98", x"99", x"99", x"99", x"9b", x"98", x"99", x"9b", x"9a", 
        x"9a", x"99", x"9a", x"9b", x"9b", x"9a", x"9b", x"9b", x"9a", x"9a", x"9b", x"9b", x"9b", x"9b", x"99", 
        x"9c", x"9c", x"8b", x"7d", x"83", x"7d", x"89", x"8b", x"8b", x"8c", x"90", x"91", x"8c", x"84", x"7b", 
        x"71", x"69", x"59", x"4b", x"48", x"46", x"35", x"46", x"59", x"47", x"4d", x"49", x"47", x"49", x"4c", 
        x"4a", x"49", x"45", x"49", x"4e", x"4d", x"4b", x"49", x"4b", x"4b", x"4a", x"49", x"48", x"47", x"44", 
        x"3c", x"57", x"ce", x"e3", x"d8", x"d9", x"d8", x"dc", x"df", x"d1", x"d0", x"d0", x"d3", x"d2", x"d3", 
        x"d2", x"d2", x"d3", x"d4", x"d4", x"d4", x"d3", x"d2", x"d0", x"d3", x"d5", x"d4", x"d3", x"d2", x"d2", 
        x"d4", x"d4", x"d3", x"d3", x"d4", x"d6", x"d6", x"d4", x"d2", x"d1", x"d3", x"d3", x"d3", x"d4", x"d4", 
        x"d4", x"d5", x"d4", x"d3", x"d3", x"d3", x"d3", x"d0", x"d2", x"db", x"d1", x"d2", x"d4", x"d4", x"d3", 
        x"d0", x"d3", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ed", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ed", x"ee", x"f0", x"ef", x"ee", 
        x"ed", x"ee", x"ed", x"ee", x"ee", x"ef", x"f0", x"f1", x"f2", x"f1", x"f0", x"f1", x"e5", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f3", x"f3", x"f1", x"ec", x"e3", x"d6", x"c2", x"a7", x"83", x"65", x"50", x"42", x"3f", 
        x"4c", x"61", x"65", x"68", x"66", x"64", x"6c", x"73", x"70", x"6c", x"69", x"6a", x"67", x"64", x"6b", 
        x"74", x"86", x"90", x"7f", x"5b", x"4f", x"56", x"5b", x"64", x"79", x"7a", x"6a", x"64", x"60", x"56", 
        x"46", x"35", x"26", x"18", x"0d", x"09", x"09", x"0c", x"13", x"1b", x"2c", x"46", x"5f", x"77", x"81", 
        x"88", x"87", x"82", x"73", x"6c", x"70", x"81", x"9c", x"bc", x"d8", x"eb", x"f1", x"f2", x"f6", x"f6", 
        x"f4", x"f5", x"f4", x"f2", x"f2", x"f2", x"f1", x"f2", x"f5", x"f4", x"f2", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f4", x"f1", x"f1", x"f3", x"f3", x"f1", x"ef", x"ec", x"f4", x"f4", x"f3", 
        x"f3", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f5", x"f4", x"f0", x"ec", x"e5", x"d6", x"c1", 
        x"ae", x"a1", x"ae", x"c5", x"de", x"ee", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f3", x"f4", x"f5", 
        x"f1", x"f2", x"f1", x"ef", x"ef", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", x"f3", x"f3", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"ef", x"f1", x"f1", x"f0", x"f1", x"f3", x"f4", x"f3", x"f2", x"f2", x"f4", 
        x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f0", x"f0", x"ef", x"f0", x"f1", x"f2", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f0", 
        x"f1", x"b8", x"65", x"9f", x"93", x"91", x"99", x"9a", x"c7", x"de", x"e3", x"dd", x"a6", x"96", x"b6", 
        x"c8", x"d4", x"de", x"e4", x"e5", x"e5", x"e3", x"e2", x"e0", x"e1", x"e2", x"e4", x"e2", x"df", x"df", 
        x"df", x"dd", x"de", x"df", x"e0", x"de", x"df", x"e3", x"df", x"dc", x"dc", x"da", x"dc", x"e1", x"d4", 
        x"bf", x"bb", x"b6", x"b1", x"b0", x"a8", x"9d", x"93", x"86", x"73", x"53", x"38", x"25", x"1a", x"7f", 
        x"e3", x"e4", x"df", x"dc", x"e0", x"e5", x"e7", x"e7", x"e2", x"da", x"cd", x"b8", x"ab", x"a5", x"a3", 
        x"a7", x"a9", x"ac", x"b1", x"b3", x"b8", x"bd", x"ba", x"af", x"9b", x"79", x"53", x"36", x"29", x"20", 
        x"1f", x"33", x"47", x"52", x"5c", x"63", x"60", x"5a", x"45", x"58", x"31", x"17", x"37", x"8a", x"93", 
        x"8a", x"7b", x"69", x"69", x"76", x"7c", x"78", x"79", x"78", x"74", x"6b", x"5f", x"5c", x"64", x"75", 
        x"8f", x"a9", x"c5", x"d7", x"e1", x"e6", x"e8", x"e8", x"e8", x"e5", x"e5", x"e8", x"e5", x"e8", x"e3", 
        x"e6", x"e8", x"e9", x"ee", x"eb", x"e3", x"cf", x"af", x"8e", x"69", x"42", x"2b", x"1f", x"15", x"0f", 
        x"99", x"9a", x"9a", x"9a", x"98", x"97", x"97", x"97", x"97", x"97", x"98", x"99", x"99", x"96", x"96", 
        x"97", x"98", x"98", x"98", x"97", x"97", x"98", x"99", x"9a", x"98", x"97", x"96", x"96", x"97", x"98", 
        x"97", x"98", x"99", x"96", x"94", x"95", x"95", x"98", x"97", x"95", x"96", x"98", x"99", x"98", x"98", 
        x"96", x"96", x"96", x"97", x"98", x"97", x"98", x"98", x"98", x"98", x"98", x"99", x"98", x"98", x"98", 
        x"97", x"98", x"9a", x"99", x"97", x"99", x"9a", x"99", x"98", x"99", x"99", x"98", x"9a", x"9a", x"99", 
        x"99", x"99", x"9a", x"9a", x"99", x"9a", x"9a", x"9a", x"99", x"99", x"99", x"98", x"9a", x"9a", x"9a", 
        x"99", x"99", x"9a", x"9b", x"9a", x"9a", x"9a", x"9b", x"9c", x"9b", x"9b", x"9b", x"9a", x"9a", x"9a", 
        x"9c", x"9d", x"8a", x"7c", x"83", x"7d", x"86", x"86", x"87", x"88", x"87", x"89", x"89", x"89", x"8c", 
        x"8f", x"8f", x"92", x"88", x"76", x"50", x"39", x"43", x"57", x"46", x"4a", x"47", x"49", x"4a", x"4e", 
        x"4c", x"4e", x"4c", x"4d", x"4d", x"4d", x"4f", x"4e", x"50", x"4c", x"49", x"4a", x"48", x"40", x"40", 
        x"39", x"55", x"cd", x"e1", x"d7", x"d8", x"d6", x"da", x"df", x"d1", x"d2", x"d0", x"d3", x"d2", x"d2", 
        x"d1", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d2", x"d1", x"d3", x"d5", x"d3", x"d4", x"d3", x"d1", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d4", x"d2", x"d1", x"d2", x"d3", x"d4", x"d3", x"d4", 
        x"d6", x"d5", x"d4", x"d3", x"d3", x"d4", x"d3", x"d0", x"d2", x"dc", x"d1", x"d2", x"d4", x"d4", x"d2", 
        x"d0", x"d4", x"ed", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f0", x"f0", x"f0", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f1", x"f2", x"f2", x"f2", x"f0", x"f1", x"e4", x"ee", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f2", x"ee", x"ea", x"e3", x"d4", x"b7", x"9c", 
        x"80", x"66", x"4a", x"49", x"5c", x"68", x"6a", x"67", x"6c", x"74", x"76", x"76", x"76", x"77", x"78", 
        x"6c", x"5e", x"53", x"51", x"48", x"53", x"59", x"6c", x"75", x"64", x"5c", x"64", x"70", x"6c", x"67", 
        x"67", x"68", x"69", x"62", x"55", x"44", x"30", x"24", x"1b", x"10", x"0c", x"0e", x"11", x"17", x"25", 
        x"3c", x"57", x"6a", x"75", x"84", x"89", x"80", x"72", x"6a", x"6e", x"7e", x"96", x"ad", x"c8", x"df", 
        x"e9", x"f1", x"f6", x"f4", x"f2", x"f3", x"f2", x"f1", x"f3", x"f5", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f3", x"f3", x"f5", x"f5", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"eb", x"f4", x"f3", x"f3", 
        x"f3", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f4", x"f4", x"ef", 
        x"ea", x"e1", x"cc", x"b6", x"a9", x"ad", x"bd", x"d0", x"e3", x"ea", x"f0", x"f4", x"f5", x"f3", x"f1", 
        x"ef", x"f2", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f2", x"f3", x"f2", x"ef", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f0", x"f1", x"f1", x"f1", x"f3", x"f2", x"f2", x"f1", 
        x"f2", x"b4", x"49", x"9d", x"c8", x"cb", x"c9", x"b4", x"cf", x"e4", x"e6", x"e5", x"e0", x"da", x"e3", 
        x"e5", x"e5", x"e0", x"df", x"e3", x"e3", x"e2", x"e2", x"e2", x"e3", x"e3", x"e3", x"e2", x"e2", x"e1", 
        x"e0", x"e0", x"e2", x"e0", x"de", x"dd", x"de", x"e0", x"e0", x"e0", x"e1", x"dd", x"d8", x"ce", x"bb", 
        x"a8", x"9d", x"93", x"87", x"74", x"5c", x"3f", x"29", x"1f", x"1b", x"25", x"26", x"27", x"2a", x"86", 
        x"e0", x"e5", x"e2", x"e3", x"df", x"d2", x"c6", x"b6", x"ac", x"a7", x"a9", x"ad", x"af", x"ae", x"b1", 
        x"b6", x"ba", x"b9", x"af", x"a2", x"8e", x"69", x"44", x"2d", x"27", x"28", x"2e", x"3e", x"50", x"5c", 
        x"62", x"65", x"61", x"57", x"52", x"4f", x"4f", x"56", x"5a", x"78", x"4e", x"21", x"3b", x"8f", x"96", 
        x"8c", x"8b", x"7c", x"6c", x"67", x"63", x"63", x"63", x"68", x"75", x"86", x"9e", x"b8", x"cf", x"e1", 
        x"e8", x"e8", x"ea", x"e9", x"e7", x"e7", x"e8", x"e5", x"e5", x"e6", x"e6", x"e6", x"ea", x"e8", x"e6", 
        x"de", x"cc", x"b4", x"99", x"74", x"4f", x"2e", x"1c", x"19", x"18", x"16", x"1f", x"31", x"4f", x"61", 
        x"99", x"9a", x"99", x"98", x"98", x"98", x"9a", x"98", x"97", x"98", x"99", x"9a", x"98", x"96", x"95", 
        x"96", x"97", x"97", x"97", x"96", x"96", x"97", x"97", x"98", x"97", x"96", x"95", x"95", x"96", x"97", 
        x"96", x"97", x"97", x"96", x"94", x"95", x"95", x"97", x"97", x"95", x"96", x"97", x"98", x"97", x"97", 
        x"96", x"97", x"96", x"97", x"97", x"98", x"99", x"98", x"98", x"97", x"98", x"98", x"97", x"98", x"99", 
        x"98", x"99", x"9b", x"99", x"96", x"97", x"99", x"98", x"98", x"9a", x"99", x"98", x"9b", x"9a", x"98", 
        x"98", x"98", x"9a", x"9b", x"99", x"9a", x"9a", x"9a", x"99", x"98", x"97", x"99", x"9a", x"9a", x"9a", 
        x"99", x"99", x"9a", x"9a", x"99", x"99", x"9a", x"9b", x"9b", x"9a", x"9b", x"9b", x"98", x"9a", x"9b", 
        x"9c", x"9c", x"89", x"7c", x"84", x"7d", x"87", x"88", x"88", x"88", x"87", x"88", x"88", x"87", x"88", 
        x"88", x"87", x"88", x"8a", x"79", x"4e", x"3c", x"41", x"58", x"48", x"48", x"48", x"4c", x"4a", x"4c", 
        x"4c", x"4d", x"4f", x"50", x"4e", x"50", x"51", x"4d", x"4d", x"4d", x"4c", x"51", x"51", x"4c", x"4f", 
        x"43", x"59", x"cd", x"e0", x"d8", x"d9", x"d6", x"d8", x"dd", x"d1", x"d3", x"d2", x"d4", x"d1", x"d2", 
        x"d2", x"d2", x"d2", x"d1", x"d2", x"d2", x"d3", x"d2", x"d1", x"d2", x"d3", x"d2", x"d3", x"d3", x"d1", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d5", x"d4", x"d4", x"d3", x"d1", x"d2", x"d2", x"d2", x"d2", x"d4", 
        x"d5", x"d4", x"d3", x"d3", x"d4", x"d5", x"d3", x"d1", x"d3", x"dd", x"d3", x"d2", x"d3", x"d5", x"d1", 
        x"d0", x"d5", x"ec", x"ef", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"e4", x"ee", x"ef", 
        x"ef", x"ef", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f1", 
        x"ea", x"dc", x"c5", x"aa", x"8f", x"6b", x"48", x"43", x"44", x"44", x"42", x"43", x"48", x"4e", x"49", 
        x"50", x"5a", x"57", x"5b", x"51", x"53", x"5f", x"67", x"6b", x"6d", x"6b", x"69", x"6d", x"6a", x"68", 
        x"69", x"68", x"67", x"6a", x"6d", x"6f", x"6c", x"5e", x"55", x"43", x"37", x"2c", x"23", x"12", x"0f", 
        x"0d", x"0c", x"11", x"1e", x"39", x"5e", x"6f", x"7d", x"87", x"87", x"7c", x"6a", x"5f", x"69", x"7f", 
        x"97", x"b3", x"cd", x"dd", x"e9", x"f3", x"f5", x"f1", x"f1", x"f5", x"f3", x"f1", x"f3", x"f2", x"f3", 
        x"f2", x"f0", x"f2", x"f4", x"f1", x"f1", x"f2", x"f2", x"f0", x"f1", x"f1", x"eb", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"f3", x"f2", x"f0", x"f1", x"f4", 
        x"f5", x"f4", x"f4", x"f1", x"ea", x"d7", x"bf", x"ae", x"a8", x"b6", x"c8", x"da", x"e6", x"ec", x"ef", 
        x"f2", x"f3", x"f1", x"ed", x"ee", x"f1", x"f3", x"f3", x"f2", x"f0", x"f2", x"f4", x"f4", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f1", x"ef", x"f1", x"f3", x"f3", x"f1", x"f0", x"f0", x"f1", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"be", x"60", x"b4", x"de", x"d3", x"dc", x"d8", x"de", x"e4", x"e0", x"df", x"e2", x"e7", x"e3", 
        x"e2", x"e3", x"de", x"e3", x"e2", x"e3", x"e4", x"e4", x"e3", x"e1", x"df", x"e2", x"e3", x"e2", x"de", 
        x"dd", x"dd", x"df", x"e0", x"de", x"dd", x"df", x"de", x"db", x"d1", x"be", x"a7", x"95", x"88", x"7d", 
        x"6d", x"53", x"3f", x"28", x"1a", x"19", x"1e", x"25", x"2d", x"32", x"40", x"5b", x"76", x"87", x"b1", 
        x"d6", x"d0", x"c1", x"b6", x"a5", x"a0", x"a3", x"a9", x"ab", x"af", x"b4", x"b8", x"b7", x"b6", x"b2", 
        x"a4", x"8d", x"6a", x"41", x"2a", x"23", x"24", x"2d", x"3f", x"59", x"64", x"6b", x"68", x"60", x"5b", 
        x"57", x"50", x"51", x"5b", x"6a", x"73", x"7c", x"83", x"7d", x"92", x"59", x"1f", x"38", x"86", x"8e", 
        x"81", x"7e", x"77", x"71", x"6c", x"70", x"84", x"a2", x"be", x"d7", x"e8", x"ed", x"eb", x"e9", x"eb", 
        x"ed", x"e9", x"e6", x"e5", x"e4", x"e7", x"ea", x"ea", x"e9", x"e7", x"e1", x"d3", x"c4", x"aa", x"8b", 
        x"69", x"3d", x"1f", x"12", x"15", x"15", x"1a", x"21", x"35", x"50", x"68", x"7a", x"8b", x"8e", x"8a", 
        x"99", x"99", x"99", x"98", x"97", x"98", x"99", x"98", x"98", x"98", x"98", x"99", x"98", x"97", x"97", 
        x"98", x"99", x"99", x"98", x"98", x"99", x"99", x"99", x"99", x"99", x"98", x"98", x"97", x"97", x"97", 
        x"97", x"97", x"97", x"96", x"96", x"96", x"97", x"97", x"97", x"97", x"97", x"98", x"98", x"97", x"97", 
        x"97", x"97", x"97", x"97", x"96", x"98", x"99", x"98", x"97", x"96", x"97", x"97", x"97", x"99", x"99", 
        x"97", x"98", x"9a", x"9a", x"97", x"97", x"9a", x"9a", x"9a", x"9b", x"9a", x"98", x"9a", x"9a", x"99", 
        x"99", x"99", x"9a", x"9a", x"99", x"99", x"99", x"99", x"99", x"98", x"99", x"9b", x"9b", x"9b", x"9a", 
        x"99", x"9a", x"9b", x"9b", x"9a", x"99", x"9a", x"9a", x"9a", x"99", x"9b", x"9c", x"99", x"9a", x"9b", 
        x"9c", x"9a", x"88", x"7c", x"85", x"7d", x"87", x"89", x"88", x"88", x"86", x"87", x"87", x"88", x"87", 
        x"88", x"87", x"89", x"87", x"7b", x"65", x"4a", x"41", x"57", x"48", x"47", x"4f", x"5a", x"53", x"50", 
        x"4d", x"4b", x"4d", x"4a", x"48", x"4d", x"4d", x"4f", x"53", x"4f", x"4d", x"51", x"51", x"50", x"51", 
        x"46", x"5e", x"cf", x"e0", x"da", x"db", x"d8", x"d8", x"dc", x"d1", x"d4", x"d2", x"d4", x"d1", x"d2", 
        x"d2", x"d2", x"d2", x"d1", x"d1", x"d2", x"d3", x"d1", x"d0", x"d1", x"d3", x"d3", x"d2", x"d2", x"d2", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d4", x"d4", x"d2", x"d2", x"d1", x"d2", x"d2", x"d2", 
        x"d4", x"d5", x"d5", x"d4", x"d4", x"d5", x"d3", x"d2", x"d3", x"dd", x"d4", x"d2", x"d4", x"d5", x"d0", 
        x"d0", x"d6", x"eb", x"ef", x"f0", x"ee", x"f0", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", 
        x"ef", x"f0", x"f0", x"f1", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"e4", x"ee", x"ef", 
        x"ef", x"ef", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f1", x"f2", x"f2", 
        x"f1", x"f2", x"f1", x"ee", x"e9", x"db", x"c6", x"a8", x"8f", x"74", x"5f", x"54", x"53", x"54", x"52", 
        x"54", x"5a", x"5a", x"5f", x"53", x"56", x"5f", x"65", x"69", x"6a", x"6a", x"68", x"68", x"65", x"64", 
        x"65", x"66", x"68", x"67", x"65", x"65", x"68", x"61", x"63", x"59", x"5c", x"61", x"64", x"4c", x"3c", 
        x"2a", x"1c", x"16", x"12", x"10", x"12", x"17", x"26", x"3d", x"51", x"65", x"77", x"7f", x"83", x"7e", 
        x"73", x"6f", x"75", x"86", x"9a", x"b2", x"c8", x"d6", x"e4", x"f1", x"f5", x"f4", x"f2", x"f2", x"f1", 
        x"f3", x"f4", x"f4", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"eb", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f3", x"f4", x"f0", x"ea", x"e0", x"cf", x"bc", x"b1", x"b7", x"c4", x"d0", 
        x"de", x"e6", x"ec", x"f0", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f1", x"f0", x"f1", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f3", x"f2", x"f1", x"ef", x"ef", x"f1", x"f3", x"f4", x"f2", 
        x"f1", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f4", x"f3", x"f4", x"f2", x"f4", x"f2", x"ee", x"ee", x"ee", 
        x"eb", x"d8", x"b3", x"da", x"e3", x"e1", x"e1", x"e6", x"e5", x"e6", x"e4", x"e4", x"e2", x"e6", x"e3", 
        x"e5", x"e4", x"df", x"e6", x"e3", x"e2", x"e2", x"e2", x"e1", x"e1", x"e0", x"e0", x"e1", x"e1", x"e1", 
        x"e2", x"e1", x"db", x"d8", x"d1", x"c9", x"ba", x"a6", x"9a", x"8a", x"74", x"5e", x"4e", x"3e", x"2d", 
        x"21", x"19", x"20", x"27", x"2c", x"3b", x"4a", x"5d", x"78", x"8e", x"a1", x"a7", x"ab", x"ac", x"a6", 
        x"a3", x"9d", x"9e", x"a4", x"a9", x"b2", x"b1", x"b7", x"bc", x"b7", x"a9", x"97", x"81", x"69", x"4a", 
        x"2f", x"29", x"2c", x"34", x"47", x"58", x"5e", x"62", x"63", x"5e", x"5a", x"54", x"53", x"58", x"62", 
        x"6d", x"7a", x"7a", x"80", x"84", x"84", x"84", x"7e", x"7b", x"91", x"5c", x"23", x"36", x"72", x"85", 
        x"83", x"87", x"96", x"af", x"c6", x"d5", x"e1", x"e6", x"e8", x"ea", x"e8", x"e7", x"e8", x"e7", x"e6", 
        x"e8", x"ea", x"e9", x"e9", x"e8", x"e2", x"d8", x"ca", x"b9", x"a3", x"91", x"7d", x"44", x"1e", x"13", 
        x"0e", x"12", x"21", x"2c", x"43", x"56", x"6e", x"7c", x"87", x"8d", x"8c", x"89", x"85", x"81", x"7f", 
        x"97", x"99", x"9a", x"99", x"97", x"96", x"96", x"98", x"99", x"98", x"97", x"97", x"98", x"99", x"98", 
        x"96", x"98", x"98", x"98", x"98", x"98", x"9a", x"9a", x"99", x"99", x"9a", x"9a", x"99", x"98", x"99", 
        x"99", x"98", x"98", x"98", x"99", x"98", x"9a", x"99", x"98", x"99", x"99", x"98", x"98", x"96", x"97", 
        x"98", x"99", x"98", x"97", x"96", x"97", x"98", x"97", x"96", x"96", x"96", x"97", x"96", x"97", x"99", 
        x"97", x"98", x"9a", x"99", x"97", x"99", x"9b", x"9b", x"9b", x"9c", x"9b", x"99", x"99", x"9a", x"9a", 
        x"9a", x"9a", x"9a", x"99", x"99", x"99", x"99", x"99", x"99", x"9a", x"9c", x"9d", x"9c", x"9b", x"9a", 
        x"9a", x"9a", x"9a", x"9c", x"9b", x"9a", x"9a", x"9a", x"99", x"98", x"9b", x"9e", x"9b", x"9b", x"9b", 
        x"9c", x"9a", x"86", x"7c", x"87", x"7d", x"87", x"8a", x"88", x"88", x"89", x"88", x"87", x"86", x"86", 
        x"86", x"87", x"89", x"84", x"83", x"8f", x"61", x"43", x"58", x"43", x"45", x"6e", x"92", x"8b", x"7f", 
        x"6f", x"63", x"5b", x"53", x"51", x"4f", x"48", x"4b", x"4c", x"4f", x"51", x"53", x"51", x"50", x"52", 
        x"4a", x"5f", x"ce", x"de", x"d9", x"dc", x"d7", x"d8", x"dc", x"d1", x"d5", x"d2", x"d3", x"d1", x"d2", 
        x"d4", x"d3", x"d2", x"d2", x"d2", x"d2", x"d3", x"d0", x"d0", x"d2", x"d3", x"d5", x"d3", x"d1", x"d2", 
        x"d4", x"d4", x"d3", x"d3", x"d3", x"d5", x"d6", x"d3", x"d3", x"d2", x"d1", x"d0", x"d2", x"d2", x"d1", 
        x"d4", x"d6", x"d6", x"d5", x"d4", x"d3", x"d3", x"d4", x"d3", x"dd", x"d5", x"d2", x"d3", x"d5", x"d0", 
        x"d1", x"d6", x"ec", x"f0", x"f0", x"ee", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"f0", x"f1", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"e4", x"ee", x"ef", 
        x"ef", x"ef", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f3", x"f4", x"f3", x"f2", 
        x"f1", x"ee", x"eb", x"ef", x"f2", x"ef", x"f2", x"f7", x"f2", x"e8", x"d8", x"ba", x"99", x"7c", x"66", 
        x"54", x"4f", x"51", x"54", x"4a", x"4f", x"61", x"6a", x"6b", x"65", x"67", x"6a", x"67", x"67", x"6a", 
        x"6a", x"6b", x"6c", x"6b", x"68", x"66", x"67", x"5f", x"5b", x"54", x"5c", x"5f", x"60", x"56", x"4e", 
        x"46", x"3f", x"36", x"2d", x"23", x"20", x"1b", x"14", x"0e", x"0c", x"10", x"1d", x"33", x"4e", x"68", 
        x"7a", x"87", x"87", x"7b", x"6d", x"66", x"6c", x"77", x"8e", x"ae", x"c5", x"d7", x"e8", x"f3", x"f4", 
        x"f2", x"f3", x"f4", x"f2", x"f3", x"f3", x"f2", x"f3", x"f5", x"f4", x"f0", x"eb", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f4", x"f5", x"f5", x"f3", 
        x"f2", x"f2", x"f3", x"f2", x"f0", x"f1", x"f1", x"f1", x"f4", x"f7", x"f7", x"ee", x"d9", x"c4", x"b5", 
        x"b3", x"be", x"ca", x"d6", x"e1", x"ec", x"f3", x"f5", x"f4", x"f1", x"ef", x"ef", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f0", x"ef", x"f1", x"f3", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f4", x"f1", x"f4", x"f0", x"e8", x"e7", x"e4", 
        x"e2", x"e7", x"e9", x"ea", x"e1", x"e0", x"df", x"e5", x"e1", x"e2", x"e1", x"e3", x"e4", x"e2", x"e0", 
        x"e2", x"e1", x"e2", x"e4", x"e4", x"e2", x"e1", x"e1", x"e2", x"e3", x"e4", x"e3", x"e0", x"dd", x"da", 
        x"d4", x"c6", x"b2", x"a1", x"93", x"82", x"6c", x"56", x"47", x"37", x"23", x"16", x"16", x"1b", x"25", 
        x"33", x"3b", x"48", x"58", x"74", x"94", x"ab", x"b4", x"b4", x"b0", x"a8", x"a3", x"a1", x"a6", x"a4", 
        x"a2", x"aa", x"af", x"ad", x"af", x"ab", x"b6", x"b2", x"a5", x"6e", x"40", x"21", x"0c", x"1a", x"28", 
        x"3d", x"56", x"64", x"65", x"63", x"5e", x"55", x"4d", x"47", x"49", x"5a", x"6d", x"7c", x"86", x"8a", 
        x"8b", x"88", x"80", x"80", x"7d", x"75", x"72", x"6e", x"6d", x"81", x"64", x"4c", x"6a", x"9e", x"bc", 
        x"d4", x"e6", x"ef", x"ed", x"eb", x"e8", x"e5", x"e6", x"e7", x"e6", x"e4", x"e8", x"ec", x"eb", x"eb", 
        x"e9", x"e0", x"d4", x"c6", x"b2", x"97", x"80", x"72", x"68", x"67", x"76", x"8a", x"36", x"05", x"05", 
        x"0a", x"30", x"6a", x"84", x"8d", x"8f", x"8d", x"8e", x"89", x"83", x"7f", x"82", x"82", x"7e", x"7d", 
        x"97", x"99", x"9a", x"9a", x"99", x"97", x"97", x"99", x"99", x"99", x"97", x"97", x"97", x"9a", x"97", 
        x"96", x"98", x"99", x"98", x"98", x"99", x"99", x"97", x"96", x"96", x"97", x"97", x"96", x"96", x"99", 
        x"99", x"98", x"97", x"98", x"9a", x"99", x"9b", x"98", x"97", x"98", x"98", x"97", x"97", x"97", x"97", 
        x"98", x"99", x"99", x"98", x"97", x"97", x"98", x"98", x"98", x"97", x"98", x"99", x"98", x"98", x"9a", 
        x"99", x"9a", x"9b", x"9a", x"98", x"9a", x"9b", x"9b", x"9a", x"9c", x"9c", x"99", x"99", x"9a", x"9a", 
        x"9a", x"9a", x"9a", x"99", x"9a", x"9a", x"9a", x"99", x"99", x"9b", x"9c", x"9c", x"9c", x"9b", x"9a", 
        x"9b", x"9a", x"99", x"9b", x"9b", x"9a", x"9a", x"9a", x"9a", x"99", x"9a", x"9d", x"9e", x"9c", x"9b", 
        x"9e", x"9d", x"86", x"7b", x"87", x"7c", x"86", x"8a", x"87", x"87", x"89", x"89", x"8a", x"8c", x"8a", 
        x"88", x"88", x"88", x"82", x"81", x"95", x"5c", x"3c", x"57", x"45", x"41", x"67", x"8f", x"8c", x"8c", 
        x"8d", x"8e", x"8e", x"86", x"81", x"76", x"6f", x"65", x"4b", x"49", x"4c", x"4b", x"4d", x"49", x"4f", 
        x"47", x"5d", x"cc", x"dd", x"d8", x"db", x"d6", x"d8", x"dd", x"d1", x"d4", x"d1", x"d2", x"d1", x"d3", 
        x"d5", x"d4", x"d4", x"d4", x"d3", x"d3", x"d2", x"d0", x"d2", x"d3", x"d3", x"d6", x"d3", x"d1", x"d2", 
        x"d4", x"d4", x"d3", x"d3", x"d4", x"d6", x"d6", x"d3", x"d3", x"d2", x"d1", x"d0", x"d2", x"d2", x"d2", 
        x"d5", x"d7", x"d6", x"d5", x"d3", x"d2", x"d3", x"d4", x"d2", x"dc", x"d5", x"d1", x"d4", x"d5", x"d1", 
        x"d1", x"d6", x"ee", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"ee", x"ee", x"ef", 
        x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"e4", x"ee", x"ef", 
        x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f3", x"f3", x"f1", x"f0", 
        x"f0", x"f0", x"ed", x"f1", x"f2", x"ed", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"ef", x"eb", x"dc", 
        x"c6", x"af", x"9a", x"7f", x"64", x"58", x"58", x"5c", x"63", x"67", x"6b", x"6d", x"6b", x"69", x"65", 
        x"64", x"65", x"68", x"6c", x"6d", x"6c", x"6d", x"63", x"59", x"54", x"51", x"43", x"38", x"31", x"33", 
        x"3a", x"40", x"3e", x"3d", x"38", x"36", x"2e", x"29", x"25", x"1d", x"14", x"10", x"11", x"13", x"16", 
        x"1f", x"30", x"45", x"58", x"6b", x"7a", x"83", x"86", x"7f", x"77", x"7a", x"81", x"90", x"a6", x"bc", 
        x"d2", x"e5", x"f2", x"f6", x"f8", x"f8", x"f5", x"f2", x"f1", x"f2", x"f0", x"eb", x"f3", x"f2", x"f3", 
        x"f3", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f4", x"f5", x"f3", x"f1", x"f1", 
        x"f1", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", 
        x"e2", x"d8", x"ca", x"bf", x"c0", x"c5", x"c9", x"d8", x"e4", x"ef", x"f5", x"f5", x"f2", x"f0", x"f2", 
        x"f2", x"f1", x"f1", x"f0", x"ee", x"f1", x"f3", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f4", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f3", x"ef", x"f3", x"ed", x"e2", x"e2", x"e2", 
        x"e5", x"e7", x"e5", x"e1", x"e7", x"e5", x"e4", x"e3", x"e2", x"e6", x"e5", x"e5", x"e5", x"e5", x"e1", 
        x"e2", x"e2", x"e4", x"e0", x"e2", x"e4", x"e6", x"e6", x"e2", x"d8", x"cf", x"c9", x"bd", x"b0", x"a2", 
        x"92", x"79", x"60", x"4c", x"41", x"37", x"28", x"1e", x"1e", x"24", x"2a", x"38", x"4b", x"59", x"6b", 
        x"84", x"94", x"9e", x"a5", x"a7", x"a6", x"a2", x"a1", x"a4", x"a4", x"a9", x"ab", x"a9", x"aa", x"ab", 
        x"ab", x"ad", x"b0", x"ad", x"a8", x"74", x"7f", x"90", x"7e", x"2f", x"0f", x"0c", x"14", x"4d", x"62", 
        x"51", x"48", x"46", x"4a", x"4f", x"59", x"68", x"72", x"7b", x"84", x"85", x"86", x"86", x"85", x"84", 
        x"80", x"73", x"67", x"65", x"69", x"6b", x"77", x"89", x"9b", x"ba", x"c9", x"d1", x"df", x"e7", x"ea", 
        x"eb", x"e9", x"e7", x"e8", x"e8", x"e9", x"e9", x"eb", x"ed", x"ec", x"eb", x"e4", x"d6", x"c5", x"b1", 
        x"9a", x"87", x"7a", x"78", x"7b", x"80", x"87", x"91", x"9a", x"a0", x"a7", x"b2", x"4e", x"12", x"08", 
        x"14", x"3b", x"70", x"78", x"7b", x"80", x"81", x"81", x"7f", x"7f", x"7f", x"81", x"81", x"82", x"81", 
        x"98", x"9a", x"9b", x"9b", x"9a", x"9a", x"9b", x"99", x"99", x"9a", x"99", x"97", x"98", x"99", x"97", 
        x"96", x"98", x"99", x"98", x"98", x"99", x"99", x"98", x"97", x"97", x"99", x"99", x"98", x"97", x"98", 
        x"99", x"97", x"95", x"98", x"9a", x"99", x"9a", x"96", x"95", x"97", x"97", x"95", x"96", x"97", x"98", 
        x"98", x"98", x"98", x"98", x"98", x"98", x"99", x"99", x"99", x"99", x"9a", x"9b", x"9b", x"9b", x"9b", 
        x"99", x"99", x"9c", x"9c", x"9a", x"9b", x"9b", x"9a", x"99", x"9a", x"9a", x"99", x"9a", x"9a", x"99", 
        x"99", x"99", x"9a", x"9a", x"9b", x"9b", x"9b", x"9b", x"9a", x"9a", x"9a", x"9c", x"9b", x"9b", x"9b", 
        x"9c", x"9b", x"98", x"9a", x"9a", x"99", x"9a", x"9b", x"9c", x"9c", x"99", x"9b", x"9f", x"9c", x"9b", 
        x"9f", x"a0", x"87", x"7a", x"87", x"7c", x"86", x"8a", x"86", x"86", x"87", x"87", x"89", x"8c", x"8a", 
        x"88", x"88", x"89", x"88", x"82", x"91", x"5c", x"3d", x"56", x"48", x"41", x"68", x"8f", x"89", x"86", 
        x"86", x"87", x"8a", x"8d", x"8d", x"8b", x"94", x"81", x"4b", x"3b", x"3d", x"4f", x"6b", x"55", x"55", 
        x"4c", x"5e", x"cc", x"de", x"da", x"dc", x"d7", x"d9", x"dd", x"d2", x"d4", x"d0", x"d1", x"d1", x"d4", 
        x"d5", x"d4", x"d5", x"d5", x"d4", x"d3", x"d2", x"d0", x"d3", x"d3", x"d2", x"d5", x"d3", x"d1", x"d3", 
        x"d4", x"d4", x"d4", x"d4", x"d4", x"d5", x"d4", x"d2", x"d2", x"d1", x"d0", x"d0", x"d2", x"d4", x"d3", 
        x"d5", x"d6", x"d5", x"d4", x"d3", x"d2", x"d3", x"d4", x"d1", x"db", x"d4", x"d1", x"d3", x"d4", x"d1", 
        x"d0", x"d5", x"ef", x"ef", x"ed", x"ee", x"ef", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"f1", x"f0", x"f0", x"ef", x"f1", x"f1", x"f1", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ee", x"f0", x"f1", 
        x"f0", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"e4", x"ee", x"ef", 
        x"ef", x"ef", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"ee", x"f0", x"ee", x"f0", x"f2", x"f1", x"f3", x"f2", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"f3", 
        x"f4", x"f4", x"f2", x"e1", x"cb", x"b6", x"a0", x"8d", x"7c", x"6e", x"68", x"5f", x"5c", x"5e", x"5e", 
        x"62", x"64", x"62", x"62", x"64", x"66", x"68", x"61", x"5b", x"59", x"47", x"33", x"30", x"34", x"39", 
        x"3d", x"3c", x"39", x"37", x"2b", x"27", x"1f", x"1c", x"1d", x"18", x"12", x"15", x"1a", x"1b", x"16", 
        x"13", x"13", x"12", x"15", x"22", x"32", x"46", x"5f", x"74", x"7c", x"80", x"81", x"7a", x"7a", x"7c", 
        x"85", x"96", x"ac", x"c1", x"d6", x"e6", x"f1", x"f2", x"f3", x"f4", x"f2", x"ec", x"f4", x"f3", x"f3", 
        x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f4", x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f4", 
        x"f4", x"f4", x"f3", x"f4", x"f4", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", 
        x"f3", x"f5", x"f2", x"e9", x"dd", x"cf", x"c4", x"c1", x"c2", x"c7", x"d4", x"e2", x"ed", x"f0", x"f2", 
        x"f2", x"f1", x"f1", x"f0", x"ef", x"f2", x"f4", x"f2", x"f2", x"f2", x"f3", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f3", x"f4", x"f4", x"f3", x"f0", x"f1", x"f2", x"f3", x"f2", x"f1", x"f0", x"ef", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"ef", x"f3", x"ed", x"e3", x"e3", x"e5", 
        x"e7", x"e4", x"e1", x"e5", x"e5", x"e3", x"e1", x"e0", x"e4", x"e6", x"e3", x"e5", x"e4", x"e5", x"e1", 
        x"e3", x"e3", x"e6", x"e5", x"e4", x"dc", x"d2", x"c8", x"bc", x"ad", x"a0", x"90", x"79", x"5f", x"4a", 
        x"3c", x"30", x"26", x"21", x"20", x"21", x"27", x"34", x"43", x"59", x"6b", x"7f", x"95", x"a0", x"a8", 
        x"ab", x"ac", x"a7", x"9f", x"9c", x"9d", x"9e", x"a4", x"a6", x"a4", x"a9", x"aa", x"ab", x"ac", x"af", 
        x"b0", x"af", x"ae", x"af", x"ab", x"51", x"51", x"9e", x"a0", x"43", x"1f", x"17", x"17", x"58", x"6c", 
        x"5a", x"5a", x"60", x"71", x"7e", x"83", x"86", x"88", x"89", x"85", x"81", x"7a", x"74", x"6f", x"6c", 
        x"6d", x"71", x"79", x"8a", x"9e", x"b1", x"c6", x"da", x"e6", x"ed", x"ef", x"ee", x"e9", x"e6", x"e5", 
        x"e7", x"e5", x"e7", x"ea", x"eb", x"eb", x"e9", x"e2", x"d4", x"c3", x"ae", x"95", x"82", x"79", x"76", 
        x"78", x"7e", x"89", x"96", x"a2", x"aa", x"ae", x"ae", x"b3", x"b2", x"b6", x"c0", x"63", x"1c", x"0a", 
        x"11", x"33", x"69", x"76", x"7b", x"7d", x"7c", x"7f", x"7f", x"81", x"81", x"82", x"81", x"7f", x"7f", 
        x"9a", x"9a", x"9a", x"99", x"99", x"9a", x"9a", x"9a", x"9a", x"9b", x"9a", x"97", x"96", x"96", x"97", 
        x"99", x"9a", x"99", x"98", x"97", x"99", x"99", x"97", x"97", x"98", x"99", x"98", x"98", x"97", x"99", 
        x"99", x"9a", x"99", x"98", x"98", x"99", x"99", x"98", x"98", x"99", x"98", x"98", x"98", x"98", x"99", 
        x"9a", x"9b", x"9a", x"99", x"98", x"99", x"97", x"97", x"98", x"98", x"9b", x"9b", x"99", x"99", x"99", 
        x"97", x"99", x"9b", x"9c", x"9b", x"9a", x"9a", x"99", x"99", x"99", x"99", x"99", x"9b", x"9a", x"9a", 
        x"9a", x"9a", x"9a", x"9b", x"9b", x"9b", x"9b", x"9b", x"9a", x"9a", x"9a", x"99", x"9a", x"9b", x"9d", 
        x"9e", x"9d", x"99", x"9b", x"9b", x"9a", x"9c", x"9e", x"9d", x"9d", x"9c", x"9d", x"9d", x"9c", x"9b", 
        x"9d", x"9f", x"88", x"77", x"86", x"7d", x"87", x"8b", x"89", x"87", x"88", x"89", x"89", x"8b", x"8b", 
        x"88", x"87", x"89", x"8a", x"83", x"8f", x"5d", x"3d", x"57", x"49", x"40", x"69", x"90", x"8a", x"8a", 
        x"89", x"86", x"88", x"8b", x"89", x"88", x"90", x"82", x"47", x"39", x"38", x"5b", x"86", x"62", x"5e", 
        x"55", x"63", x"cd", x"df", x"db", x"dd", x"d9", x"db", x"dd", x"d1", x"d3", x"d1", x"d0", x"d2", x"d2", 
        x"d2", x"d2", x"d4", x"d5", x"d5", x"d4", x"d3", x"d2", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d3", 
        x"d3", x"d3", x"d5", x"d6", x"d5", x"d4", x"d3", x"d3", x"d2", x"d2", x"d1", x"d1", x"d2", x"d3", x"d5", 
        x"d7", x"d7", x"d5", x"d3", x"d2", x"d2", x"d4", x"d4", x"cf", x"da", x"d5", x"d2", x"d3", x"d0", x"d0", 
        x"d1", x"d4", x"ed", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", 
        x"ed", x"ed", x"ed", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ef", x"f0", x"f1", 
        x"f0", x"ef", x"ee", x"ed", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"ef", x"f0", x"ef", x"ef", x"ee", x"ef", x"f1", x"f1", x"f0", 
        x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"e6", x"ee", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"ef", 
        x"f0", x"f0", x"f2", x"f2", x"f4", x"f3", x"f1", x"ec", x"de", x"cb", x"b6", x"9c", x"81", x"67", x"50", 
        x"4b", x"54", x"5e", x"61", x"65", x"66", x"5c", x"54", x"56", x"5e", x"4e", x"3a", x"3e", x"3c", x"35", 
        x"2b", x"1b", x"14", x"17", x"11", x"0c", x"0e", x"15", x"1a", x"1c", x"1b", x"1a", x"19", x"18", x"21", 
        x"30", x"28", x"12", x"10", x"12", x"0c", x"09", x"0c", x"18", x"26", x"35", x"4f", x"6b", x"7a", x"86", 
        x"8b", x"88", x"81", x"7c", x"7d", x"88", x"a0", x"b6", x"d9", x"ed", x"f3", x"ed", x"f4", x"f2", x"f3", 
        x"f4", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f4", x"f5", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f3", x"f4", x"f3", x"ef", x"e6", x"dd", x"d0", x"c2", x"bb", x"be", x"c8", x"dc", 
        x"ec", x"f5", x"f6", x"f2", x"ee", x"f0", x"f2", x"f1", x"f3", x"f4", x"f4", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f1", x"f4", x"f6", x"f4", x"f2", x"f0", x"f1", x"f2", x"f2", x"f0", x"f0", x"f2", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f3", x"f2", x"ef", x"f4", x"ee", x"e5", x"e7", x"e6", 
        x"e4", x"e1", x"e3", x"e8", x"e3", x"e5", x"e3", x"e3", x"e4", x"e2", x"e0", x"e2", x"e6", x"eb", x"eb", 
        x"e7", x"dd", x"cf", x"c5", x"bb", x"ae", x"a3", x"94", x"77", x"53", x"3a", x"2c", x"25", x"24", x"25", 
        x"25", x"22", x"21", x"32", x"24", x"2e", x"64", x"82", x"93", x"9c", x"a2", x"a6", x"a8", x"a4", x"a2", 
        x"a0", x"a2", x"a4", x"a4", x"a3", x"a6", x"a8", x"a9", x"a9", x"a7", x"a8", x"a9", x"a6", x"a6", x"ab", 
        x"ae", x"b2", x"af", x"b0", x"b5", x"61", x"53", x"b9", x"b9", x"58", x"36", x"2f", x"27", x"78", x"98", 
        x"90", x"91", x"8f", x"8b", x"87", x"88", x"83", x"79", x"70", x"64", x"5d", x"5f", x"6e", x"86", x"9f", 
        x"b5", x"ca", x"d7", x"e2", x"e8", x"e9", x"e9", x"ec", x"eb", x"e5", x"e5", x"e5", x"e4", x"e8", x"ea", 
        x"ef", x"ef", x"ec", x"e3", x"d0", x"b2", x"96", x"7a", x"6d", x"72", x"78", x"82", x"8e", x"97", x"a4", 
        x"aa", x"a7", x"a4", x"ab", x"b6", x"bf", x"c2", x"c6", x"c4", x"c5", x"cd", x"d5", x"76", x"1b", x"0b", 
        x"13", x"3c", x"6a", x"75", x"7e", x"7b", x"7d", x"7e", x"7d", x"7f", x"80", x"81", x"80", x"81", x"80", 
        x"9b", x"9a", x"99", x"99", x"99", x"99", x"99", x"9a", x"9b", x"9b", x"9a", x"99", x"97", x"97", x"98", 
        x"9a", x"9a", x"9a", x"99", x"99", x"9a", x"9a", x"98", x"99", x"9a", x"9a", x"99", x"98", x"98", x"97", 
        x"98", x"9a", x"9a", x"97", x"97", x"99", x"99", x"9a", x"9a", x"9b", x"9a", x"9a", x"99", x"99", x"9a", 
        x"9b", x"9b", x"9b", x"9a", x"9a", x"9b", x"98", x"98", x"99", x"9a", x"9d", x"9d", x"9a", x"9a", x"9a", 
        x"99", x"99", x"99", x"99", x"99", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9b", x"9b", x"9b", 
        x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9c", x"9b", x"9c", 
        x"9c", x"9b", x"9b", x"9d", x"9c", x"9b", x"9d", x"9e", x"9d", x"9d", x"9e", x"9e", x"9c", x"9c", x"9b", 
        x"9c", x"9e", x"88", x"77", x"86", x"7e", x"88", x"8b", x"8b", x"88", x"89", x"8b", x"8a", x"8b", x"8c", 
        x"89", x"89", x"89", x"8a", x"84", x"92", x"5e", x"3c", x"58", x"49", x"3e", x"66", x"8e", x"89", x"8b", 
        x"8a", x"88", x"89", x"8a", x"88", x"88", x"8d", x"84", x"4a", x"3a", x"38", x"5a", x"85", x"62", x"60", 
        x"57", x"64", x"c9", x"dc", x"d9", x"d9", x"d6", x"d9", x"de", x"d0", x"d4", x"d3", x"d1", x"d4", x"d2", 
        x"d2", x"d2", x"d3", x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d3", x"d3", x"d3", x"d4", x"d5", x"d5", 
        x"d4", x"d3", x"d3", x"d4", x"d5", x"d4", x"d4", x"d3", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", 
        x"d6", x"d6", x"d5", x"d4", x"d3", x"d3", x"d5", x"d4", x"ce", x"da", x"d5", x"d3", x"d3", x"d2", x"d3", 
        x"d4", x"d6", x"ed", x"f0", x"ee", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"ef", x"ee", x"f0", x"f0", 
        x"f0", x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f2", x"f1", x"ef", 
        x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"e7", x"ed", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f3", x"f2", x"f3", x"f2", x"ed", x"e1", x"d4", x"c2", 
        x"ab", x"93", x"79", x"60", x"57", x"5a", x"5f", x"5d", x"5c", x"5d", x"4d", x"38", x"32", x"21", x"19", 
        x"19", x"15", x"15", x"1b", x"18", x"1a", x"1b", x"1c", x"1d", x"1e", x"21", x"22", x"2a", x"34", x"3b", 
        x"42", x"3c", x"37", x"43", x"4c", x"4d", x"44", x"34", x"26", x"19", x"0f", x"12", x"1c", x"24", x"2e", 
        x"47", x"67", x"7c", x"81", x"8a", x"8c", x"8c", x"8f", x"8b", x"8f", x"b3", x"e4", x"f4", x"f1", x"f3", 
        x"f5", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f4", x"f5", x"f5", x"f4", x"f4", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f1", x"ee", x"eb", x"e3", x"d8", x"ce", x"c7", 
        x"c4", x"cc", x"d6", x"e3", x"ee", x"f1", x"f2", x"f1", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", 
        x"f1", x"f2", x"f5", x"f4", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f3", x"f0", x"f1", x"f1", x"ef", x"f4", x"ee", x"e3", x"e5", x"e4", 
        x"e4", x"e4", x"e3", x"e4", x"e3", x"e2", x"e2", x"e5", x"e6", x"e3", x"e4", x"e4", x"db", x"cf", x"bd", 
        x"b2", x"aa", x"97", x"83", x"6f", x"54", x"3b", x"2d", x"25", x"24", x"27", x"26", x"26", x"2f", x"3d", 
        x"51", x"6c", x"8a", x"67", x"26", x"30", x"80", x"9e", x"af", x"aa", x"a6", x"a7", x"a8", x"a8", x"a7", 
        x"a7", x"a7", x"aa", x"ac", x"ac", x"ab", x"ab", x"ab", x"ab", x"aa", x"a8", x"a8", x"a8", x"ab", x"ac", 
        x"aa", x"a9", x"ad", x"b0", x"b5", x"69", x"51", x"b4", x"b9", x"5f", x"3b", x"3c", x"30", x"81", x"a3", 
        x"95", x"8e", x"88", x"7d", x"74", x"6e", x"67", x"6f", x"83", x"97", x"a9", x"be", x"d1", x"dd", x"e5", 
        x"ea", x"eb", x"ed", x"eb", x"e8", x"e6", x"e5", x"e8", x"e6", x"e7", x"ed", x"ed", x"e9", x"e1", x"d4", 
        x"c0", x"a9", x"8f", x"7b", x"74", x"78", x"7e", x"85", x"90", x"a1", x"a8", x"a9", x"aa", x"a9", x"b0", 
        x"b9", x"c1", x"c4", x"c4", x"c4", x"c4", x"c8", x"d4", x"d2", x"ce", x"cc", x"ce", x"78", x"1e", x"11", 
        x"1d", x"46", x"67", x"73", x"85", x"82", x"80", x"7f", x"7f", x"7f", x"80", x"7f", x"7d", x"7b", x"7d", 
        x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"99", 
        x"98", x"99", x"9a", x"99", x"9a", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9a", x"99", 
        x"9a", x"9b", x"9b", x"99", x"99", x"9b", x"9a", x"9a", x"9b", x"9b", x"9b", x"9a", x"9a", x"9a", x"9b", 
        x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"98", x"98", x"99", x"99", x"9c", x"9c", x"99", x"99", x"9b", 
        x"9b", x"99", x"98", x"98", x"99", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9b", x"9b", x"9b", 
        x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9c", x"9b", x"9b", x"9b", x"9b", 
        x"9a", x"9a", x"9b", x"9d", x"9b", x"9a", x"9c", x"9e", x"9c", x"9c", x"9d", x"9d", x"9c", x"9d", x"9c", 
        x"9d", x"9e", x"88", x"77", x"86", x"7e", x"87", x"8a", x"8b", x"89", x"89", x"8b", x"8a", x"8b", x"8c", 
        x"8a", x"8b", x"8b", x"8b", x"87", x"93", x"5f", x"3c", x"58", x"4b", x"40", x"67", x"8e", x"88", x"89", 
        x"88", x"88", x"8a", x"88", x"88", x"8a", x"8e", x"86", x"4d", x"3a", x"39", x"59", x"86", x"64", x"61", 
        x"58", x"66", x"c9", x"dd", x"da", x"d9", x"d6", x"da", x"df", x"d2", x"d5", x"d4", x"d3", x"d5", x"d4", 
        x"d3", x"d3", x"d3", x"d3", x"d3", x"d4", x"d5", x"d4", x"d4", x"d3", x"d3", x"d3", x"d4", x"d5", x"d6", 
        x"d4", x"d3", x"d2", x"d3", x"d4", x"d5", x"d4", x"d3", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d1", 
        x"d3", x"d4", x"d4", x"d3", x"d3", x"d4", x"d5", x"d3", x"cf", x"da", x"d6", x"d4", x"d4", x"d4", x"d4", 
        x"d5", x"d6", x"ed", x"ef", x"ed", x"ef", x"ef", x"ee", x"ed", x"ee", x"ef", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"ef", x"f0", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"e7", x"ed", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f2", x"f4", x"f3", x"f3", x"f3", 
        x"ee", x"e8", x"de", x"ca", x"b3", x"9b", x"7c", x"63", x"57", x"59", x"44", x"22", x"12", x"12", x"17", 
        x"21", x"22", x"1f", x"21", x"20", x"1e", x"1f", x"22", x"2b", x"35", x"40", x"47", x"48", x"48", x"4d", 
        x"5c", x"6a", x"71", x"73", x"73", x"78", x"80", x"7e", x"71", x"60", x"4b", x"39", x"24", x"18", x"14", 
        x"11", x"19", x"1f", x"2c", x"51", x"70", x"7e", x"80", x"62", x"4f", x"9b", x"e0", x"f3", x"f1", x"f3", 
        x"f5", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f4", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f0", x"f0", x"f4", x"f7", x"f6", x"f1", x"ee", x"eb", 
        x"e4", x"d7", x"c9", x"c5", x"c6", x"c8", x"d7", x"e9", x"ee", x"f3", x"f6", x"f4", x"f1", x"ef", x"ef", 
        x"f4", x"f6", x"f8", x"f6", x"f2", x"f1", x"f3", x"f2", x"f1", x"f2", x"f1", x"ef", x"ee", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"ef", x"f0", x"f0", x"ef", x"f4", x"ef", x"e7", x"e8", x"e4", 
        x"e3", x"e5", x"e3", x"e3", x"e5", x"e7", x"e4", x"e3", x"dc", x"ce", x"bf", x"b6", x"ac", x"9d", x"84", 
        x"6c", x"56", x"3a", x"26", x"23", x"2a", x"31", x"32", x"2f", x"31", x"39", x"55", x"6e", x"8a", x"a0", 
        x"a8", x"ae", x"ba", x"81", x"36", x"2f", x"7a", x"93", x"ab", x"ac", x"aa", x"ac", x"af", x"af", x"af", 
        x"af", x"b1", x"b0", x"ad", x"ad", x"ac", x"ac", x"ac", x"ac", x"ad", x"b1", x"ad", x"ac", x"ab", x"a9", 
        x"ab", x"ae", x"aa", x"a9", x"ae", x"69", x"4f", x"b1", x"bf", x"69", x"3d", x"3f", x"34", x"79", x"99", 
        x"86", x"78", x"6f", x"75", x"84", x"9c", x"b4", x"cb", x"de", x"e7", x"ea", x"ec", x"ec", x"ec", x"ec", 
        x"ea", x"e9", x"e9", x"eb", x"e9", x"e7", x"e8", x"e9", x"e7", x"df", x"d0", x"b9", x"a0", x"87", x"6f", 
        x"6b", x"71", x"7d", x"8e", x"a0", x"ac", x"ae", x"aa", x"a7", x"ab", x"b2", x"bd", x"c6", x"c8", x"c6", 
        x"c1", x"c3", x"c7", x"ce", x"d4", x"d1", x"cb", x"c6", x"c3", x"c6", x"cf", x"da", x"8a", x"24", x"12", 
        x"1c", x"42", x"61", x"6f", x"86", x"86", x"82", x"80", x"7f", x"7e", x"80", x"80", x"7f", x"7e", x"7f", 
        x"9a", x"9b", x"9b", x"9c", x"9b", x"9a", x"99", x"9a", x"9a", x"98", x"98", x"9a", x"9a", x"9a", x"99", 
        x"98", x"99", x"9a", x"9a", x"9a", x"99", x"99", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"99", 
        x"99", x"9a", x"99", x"98", x"98", x"9a", x"9a", x"9a", x"9b", x"9b", x"9b", x"9a", x"9a", x"9a", x"9b", 
        x"9a", x"9a", x"9a", x"9b", x"9b", x"9b", x"99", x"9a", x"9b", x"9a", x"9c", x"9c", x"98", x"97", x"9a", 
        x"9d", x"9b", x"99", x"9a", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", 
        x"9b", x"9b", x"9b", x"9b", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"98", x"99", x"9b", x"9c", 
        x"9c", x"9b", x"9c", x"9d", x"9b", x"9a", x"9c", x"9d", x"9c", x"9c", x"9c", x"9c", x"9d", x"9e", x"9d", 
        x"9d", x"9e", x"88", x"78", x"87", x"7f", x"87", x"8a", x"8b", x"8a", x"8a", x"8b", x"8b", x"8b", x"8a", 
        x"8b", x"8d", x"8b", x"8c", x"89", x"93", x"5f", x"3c", x"58", x"4a", x"3f", x"65", x"8f", x"8a", x"8c", 
        x"8c", x"8b", x"8a", x"89", x"8c", x"8e", x"8f", x"84", x"4b", x"3a", x"3a", x"58", x"85", x"67", x"63", 
        x"5d", x"6c", x"cc", x"df", x"d9", x"d4", x"d0", x"d4", x"df", x"d2", x"d4", x"d3", x"d2", x"d5", x"d4", 
        x"d3", x"d4", x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d3", x"d2", x"d2", x"d3", x"d5", x"d6", 
        x"d5", x"d3", x"d3", x"d4", x"d5", x"d5", x"d4", x"d3", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d1", 
        x"d2", x"d4", x"d3", x"d3", x"d3", x"d5", x"d6", x"d2", x"cf", x"d9", x"d7", x"d5", x"d5", x"d3", x"d2", 
        x"d3", x"d5", x"ec", x"ef", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"e7", x"ed", x"f1", 
        x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f2", x"f3", x"f3", x"f0", x"ef", 
        x"f2", x"f4", x"f5", x"f4", x"f0", x"eb", x"e2", x"d1", x"bb", x"a5", x"82", x"58", x"3b", x"23", x"1f", 
        x"24", x"2a", x"2e", x"37", x"3b", x"41", x"45", x"49", x"4b", x"4e", x"51", x"55", x"59", x"6a", x"7c", 
        x"7f", x"7b", x"7c", x"7f", x"7d", x"78", x"7b", x"7d", x"79", x"7c", x"84", x"84", x"78", x"69", x"59", 
        x"41", x"39", x"2f", x"29", x"18", x"16", x"1b", x"49", x"6e", x"9d", x"d4", x"e4", x"f2", x"f2", x"f4", 
        x"f5", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f4", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f0", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"ef", x"ef", x"ef", x"f0", x"f1", x"f5", x"f4", 
        x"f1", x"ef", x"ed", x"ec", x"db", x"c0", x"b3", x"b3", x"bf", x"ce", x"de", x"e9", x"ef", x"f2", x"f3", 
        x"f4", x"f4", x"f6", x"f5", x"f1", x"ef", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f3", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"ef", x"ef", x"ef", x"ef", x"f2", x"ef", x"e5", x"e6", x"e6", 
        x"e5", x"e7", x"e8", x"e4", x"db", x"cf", x"c1", x"b4", x"a6", x"93", x"7c", x"6a", x"51", x"39", x"28", 
        x"26", x"27", x"2b", x"2f", x"33", x"37", x"40", x"54", x"74", x"8f", x"9e", x"a9", x"af", x"b2", x"ad", 
        x"a6", x"a7", x"b4", x"88", x"49", x"35", x"79", x"93", x"b1", x"b1", x"b1", x"b2", x"b3", x"b2", x"b0", 
        x"af", x"b0", x"ae", x"ac", x"ad", x"ad", x"ae", x"ae", x"ae", x"ae", x"af", x"ab", x"ae", x"b0", x"b1", 
        x"b1", x"ad", x"ad", x"ae", x"b2", x"6f", x"4f", x"ae", x"c3", x"69", x"35", x"34", x"32", x"6e", x"98", 
        x"a1", x"ad", x"c2", x"d7", x"e1", x"e7", x"eb", x"eb", x"eb", x"eb", x"eb", x"eb", x"e8", x"ea", x"ec", 
        x"ea", x"eb", x"e9", x"ea", x"e5", x"d8", x"c7", x"b0", x"96", x"83", x"75", x"70", x"74", x"86", x"95", 
        x"a5", x"af", x"b0", x"ac", x"a9", x"b0", x"b9", x"c4", x"c9", x"c8", x"c4", x"c2", x"c5", x"cb", x"d2", 
        x"d6", x"d2", x"ca", x"c4", x"c6", x"cc", x"d1", x"d6", x"d4", x"cc", x"c7", x"cc", x"8d", x"28", x"19", 
        x"1a", x"3a", x"58", x"62", x"79", x"81", x"81", x"80", x"7e", x"7e", x"7f", x"80", x"7f", x"7f", x"7f", 
        x"9b", x"9b", x"9c", x"9c", x"9b", x"9a", x"99", x"9a", x"9a", x"98", x"97", x"98", x"98", x"97", x"98", 
        x"99", x"99", x"9a", x"9a", x"98", x"97", x"97", x"99", x"99", x"99", x"99", x"99", x"99", x"99", x"9b", 
        x"9c", x"9b", x"98", x"98", x"98", x"99", x"9a", x"9b", x"9b", x"9b", x"9b", x"9a", x"9a", x"9a", x"9b", 
        x"9a", x"9a", x"9a", x"9b", x"9b", x"9b", x"99", x"9a", x"9b", x"99", x"9a", x"9b", x"99", x"98", x"9b", 
        x"9e", x"9c", x"99", x"9a", x"9c", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", 
        x"9b", x"9b", x"9b", x"9c", x"9c", x"9d", x"9c", x"9c", x"9c", x"9c", x"9c", x"99", x"9a", x"9b", x"9c", 
        x"9c", x"9b", x"9d", x"9d", x"9b", x"9a", x"9c", x"9d", x"9d", x"9c", x"9c", x"9c", x"9c", x"9e", x"9d", 
        x"9e", x"9f", x"89", x"77", x"87", x"7f", x"88", x"8a", x"8b", x"8b", x"8c", x"8c", x"8c", x"8a", x"89", 
        x"8a", x"8b", x"8a", x"8a", x"89", x"93", x"60", x"3c", x"56", x"4b", x"41", x"65", x"8f", x"89", x"89", 
        x"88", x"8a", x"8d", x"8a", x"8d", x"8e", x"8d", x"82", x"4b", x"3a", x"3c", x"57", x"86", x"6b", x"67", 
        x"5f", x"67", x"c8", x"de", x"da", x"d7", x"d8", x"dc", x"e0", x"d1", x"d4", x"d2", x"d1", x"d4", x"d4", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d3", x"d3", x"d3", x"d5", x"d6", x"d5", x"d3", x"d4", x"d7", x"d7", 
        x"d5", x"d5", x"d5", x"d7", x"d7", x"d6", x"d4", x"d3", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d2", 
        x"d3", x"d4", x"d3", x"d2", x"d2", x"d2", x"d5", x"d1", x"d0", x"d9", x"d7", x"d5", x"d4", x"d4", x"d3", 
        x"d3", x"d6", x"ed", x"ef", x"ed", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"ef", x"ef", 
        x"ef", x"ef", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"e7", x"ed", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f2", x"f2", 
        x"f0", x"f1", x"f2", x"f0", x"f0", x"ef", x"f1", x"f5", x"f5", x"f4", x"ef", x"e5", x"d9", x"b8", x"91", 
        x"6a", x"4b", x"43", x"49", x"51", x"5a", x"5e", x"62", x"64", x"66", x"6e", x"76", x"78", x"78", x"76", 
        x"76", x"7b", x"80", x"7b", x"7c", x"7d", x"7e", x"82", x"7e", x"7e", x"83", x"84", x"84", x"8b", x"94", 
        x"8d", x"80", x"67", x"60", x"3a", x"20", x"17", x"67", x"b9", x"e0", x"dd", x"e1", x"f1", x"f3", x"f3", 
        x"f5", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", x"f2", x"f2", x"f2", x"f1", x"f3", 
        x"f2", x"f1", x"f0", x"f2", x"f2", x"ef", x"ee", x"e3", x"cb", x"b6", x"ad", x"b4", x"c2", x"d0", x"e1", 
        x"ec", x"f3", x"f4", x"f2", x"f1", x"f4", x"f1", x"f0", x"f1", x"f1", x"f2", x"f0", x"ee", x"ef", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"ee", x"ef", x"ef", x"f0", x"f1", x"ef", x"e7", x"e6", x"e6", 
        x"db", x"cd", x"c2", x"b2", x"9d", x"8b", x"77", x"5f", x"48", x"31", x"1f", x"1a", x"24", x"32", x"3f", 
        x"3e", x"37", x"41", x"57", x"77", x"90", x"a5", x"b3", x"ba", x"b5", x"ab", x"a7", x"a9", x"aa", x"a9", 
        x"aa", x"ac", x"b7", x"89", x"53", x"38", x"75", x"95", x"b7", x"b2", x"b3", x"b3", x"b4", x"b2", x"b0", 
        x"ae", x"ae", x"ad", x"ac", x"ac", x"ac", x"ac", x"ae", x"b0", x"b1", x"b1", x"b1", x"b4", x"b3", x"b1", 
        x"b0", x"aa", x"9f", x"9c", x"9e", x"66", x"4a", x"a2", x"bc", x"7d", x"6b", x"91", x"b0", x"d4", x"e6", 
        x"ee", x"ee", x"ed", x"ee", x"ef", x"eb", x"e8", x"e7", x"e8", x"eb", x"ec", x"ee", x"ea", x"e7", x"e4", 
        x"da", x"cb", x"b8", x"a1", x"85", x"74", x"70", x"6e", x"79", x"89", x"a5", x"b6", x"b8", x"b6", x"b1", 
        x"af", x"b4", x"bd", x"c7", x"cf", x"cf", x"c6", x"c6", x"ca", x"cb", x"d0", x"d6", x"d3", x"cb", x"c6", 
        x"c9", x"ce", x"d4", x"d9", x"d6", x"cb", x"c2", x"c6", x"cd", x"d3", x"d3", x"d7", x"9d", x"29", x"18", 
        x"1b", x"44", x"68", x"71", x"80", x"82", x"7b", x"79", x"79", x"7b", x"7d", x"7e", x"7d", x"7d", x"7e", 
        x"9c", x"9c", x"9b", x"9b", x"9b", x"9a", x"9a", x"9b", x"9b", x"9a", x"99", x"98", x"98", x"98", x"99", 
        x"9a", x"9a", x"9a", x"9b", x"9a", x"97", x"97", x"9a", x"9a", x"9b", x"9b", x"9a", x"9a", x"99", x"9b", 
        x"9c", x"9b", x"98", x"99", x"9b", x"9a", x"9b", x"9b", x"9c", x"9c", x"9b", x"9b", x"9b", x"9a", x"9b", 
        x"9b", x"9b", x"9b", x"9b", x"9a", x"9b", x"99", x"9b", x"9a", x"97", x"99", x"9a", x"9b", x"9a", x"9b", 
        x"9e", x"9c", x"98", x"99", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9b", x"9c", x"9c", 
        x"9c", x"9c", x"9c", x"9b", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9d", x"9e", x"9e", x"9c", x"9b", 
        x"9a", x"9b", x"9e", x"9e", x"9c", x"9a", x"9c", x"9e", x"9d", x"9c", x"9c", x"9c", x"9b", x"9d", x"9d", 
        x"9e", x"a0", x"89", x"76", x"88", x"82", x"89", x"8b", x"8a", x"8a", x"8c", x"8b", x"8c", x"8b", x"89", 
        x"8a", x"89", x"8a", x"89", x"88", x"93", x"62", x"3e", x"56", x"48", x"3f", x"61", x"8d", x"89", x"8a", 
        x"89", x"8c", x"90", x"8b", x"8a", x"8b", x"8b", x"83", x"4c", x"3b", x"3d", x"57", x"87", x"6f", x"6c", 
        x"63", x"68", x"c9", x"df", x"d9", x"d8", x"d9", x"db", x"df", x"d1", x"d3", x"d1", x"d0", x"d4", x"d4", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d3", x"d2", x"d2", x"d3", x"d4", x"d3", x"d1", x"d1", x"d5", x"d6", 
        x"d5", x"d4", x"d5", x"d6", x"d6", x"d5", x"d4", x"d3", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", 
        x"d5", x"d5", x"d4", x"d2", x"d2", x"d2", x"d5", x"d0", x"d1", x"d9", x"d7", x"d4", x"d2", x"d6", x"d7", 
        x"d7", x"d7", x"ee", x"ef", x"ed", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", 
        x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", 
        x"ee", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"e7", x"ed", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f3", x"f3", x"f1", x"f2", x"f3", x"f2", 
        x"f2", x"f3", x"f2", x"f0", x"f1", x"f3", x"f1", x"f4", x"f3", x"f3", x"f0", x"f3", x"f4", x"f2", x"ec", 
        x"e2", x"cf", x"b4", x"95", x"7d", x"70", x"6f", x"6e", x"6d", x"6d", x"6e", x"72", x"78", x"7a", x"7c", 
        x"7a", x"75", x"6e", x"6a", x"65", x"5c", x"54", x"52", x"54", x"56", x"58", x"59", x"5f", x"59", x"53", 
        x"45", x"3b", x"3c", x"70", x"62", x"4d", x"4c", x"9e", x"dd", x"dd", x"dc", x"df", x"f1", x"f4", x"f3", 
        x"f4", x"f4", x"f4", x"f4", x"f5", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f5", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f3", x"f4", 
        x"f4", x"f3", x"f0", x"f2", x"f3", x"f3", x"f6", x"f5", x"f2", x"ef", x"e4", x"d3", x"c3", x"b7", x"b3", 
        x"be", x"cb", x"d8", x"e2", x"ea", x"f2", x"f4", x"f2", x"ef", x"f0", x"f2", x"f3", x"f2", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"c8", x"9f", x"9e", 
        x"97", x"7a", x"65", x"58", x"4b", x"38", x"2b", x"23", x"26", x"2d", x"36", x"3f", x"4a", x"52", x"60", 
        x"73", x"8b", x"a1", x"ad", x"b2", x"b1", x"ad", x"a9", x"aa", x"ad", x"ae", x"ac", x"ad", x"ad", x"ae", 
        x"b1", x"b0", x"b8", x"8b", x"54", x"38", x"70", x"92", x"b6", x"b0", x"b2", x"b3", x"b4", x"b3", x"b1", 
        x"b0", x"b0", x"b0", x"ae", x"af", x"b0", x"b1", x"b2", x"b2", x"b2", x"b0", x"ab", x"a7", x"a5", x"9f", 
        x"99", x"93", x"90", x"91", x"96", x"86", x"86", x"c6", x"da", x"d6", x"db", x"e6", x"ec", x"ee", x"e9", 
        x"ec", x"ec", x"eb", x"e9", x"eb", x"ec", x"ee", x"ed", x"e9", x"e3", x"da", x"d0", x"ba", x"a7", x"99", 
        x"8a", x"80", x"7a", x"7b", x"89", x"99", x"a6", x"ab", x"b0", x"b2", x"b6", x"b6", x"b9", x"c4", x"c7", 
        x"c9", x"ce", x"ce", x"ca", x"ca", x"cf", x"cf", x"d2", x"d6", x"d1", x"ce", x"cb", x"cd", x"d3", x"d3", 
        x"d1", x"d1", x"cd", x"ca", x"cc", x"cf", x"d2", x"d3", x"cf", x"cd", x"ce", x"d5", x"a8", x"31", x"1d", 
        x"19", x"3e", x"66", x"75", x"8a", x"8d", x"83", x"7d", x"79", x"77", x"77", x"78", x"78", x"7d", x"7c", 
        x"9c", x"9c", x"9b", x"9a", x"9a", x"9b", x"9b", x"9b", x"9c", x"9c", x"9c", x"9a", x"99", x"99", x"99", 
        x"99", x"9a", x"9b", x"9c", x"9c", x"99", x"98", x"99", x"9b", x"9c", x"9c", x"9b", x"9a", x"98", x"98", 
        x"9a", x"99", x"97", x"9a", x"9c", x"9c", x"9b", x"9b", x"9c", x"9c", x"9c", x"9b", x"9a", x"99", x"9a", 
        x"9b", x"9c", x"9b", x"9a", x"9a", x"9c", x"9c", x"9c", x"9c", x"99", x"9b", x"9d", x"9d", x"9a", x"9a", 
        x"9d", x"9d", x"9a", x"9b", x"9e", x"9d", x"9d", x"9d", x"9d", x"9d", x"9d", x"9c", x"9c", x"9c", x"9c", 
        x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9d", x"9e", x"9d", x"9b", x"9b", 
        x"9c", x"9d", x"9e", x"9e", x"9c", x"9b", x"9d", x"9f", x"9d", x"9d", x"9d", x"9c", x"9b", x"9c", x"9c", 
        x"9e", x"a1", x"89", x"76", x"89", x"83", x"8b", x"8b", x"8a", x"89", x"8a", x"88", x"8b", x"8b", x"8a", 
        x"8b", x"88", x"8b", x"89", x"88", x"94", x"65", x"41", x"57", x"4c", x"43", x"64", x"90", x"8b", x"8a", 
        x"8a", x"8a", x"8e", x"8b", x"8a", x"8a", x"8b", x"84", x"4d", x"3b", x"3e", x"56", x"88", x"73", x"70", 
        x"65", x"66", x"c6", x"dd", x"d5", x"d6", x"da", x"da", x"df", x"d1", x"d3", x"d1", x"d0", x"d4", x"d5", 
        x"d5", x"d5", x"d4", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", x"d3", x"d2", x"d0", x"d0", x"d4", x"d6", 
        x"d4", x"d3", x"d2", x"d4", x"d5", x"d4", x"d3", x"d3", x"d2", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", 
        x"d5", x"d6", x"d5", x"d3", x"d2", x"d3", x"d4", x"cf", x"d2", x"d9", x"d8", x"d3", x"cf", x"d4", x"d6", 
        x"d6", x"d7", x"ee", x"f0", x"ed", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ed", x"ed", x"ee", 
        x"ef", x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ed", x"ef", x"f0", x"f0", x"ed", x"ec", 
        x"ee", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"e7", x"ed", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"f2", x"ef", x"ef", x"f0", x"ef", x"f1", x"f3", x"f4", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f2", x"f1", x"f2", x"f4", x"f5", x"f2", x"f3", x"f2", 
        x"f2", x"f5", x"f6", x"f0", x"e6", x"d3", x"bc", x"9e", x"83", x"74", x"6a", x"65", x"63", x"58", x"53", 
        x"56", x"53", x"3f", x"28", x"1c", x"14", x"0f", x"16", x"1b", x"14", x"10", x"10", x"14", x"13", x"13", 
        x"1c", x"22", x"3a", x"91", x"74", x"4d", x"56", x"ad", x"e0", x"dd", x"de", x"df", x"f2", x"f6", x"f3", 
        x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f5", x"f4", x"f3", x"f3", x"f3", x"f5", x"f4", x"f5", x"f5", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f4", x"f1", x"ee", x"f1", x"f2", x"f2", x"f4", x"f2", 
        x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f4", x"f4", x"f2", x"f3", x"f5", x"f5", x"f4", x"ef", x"de", 
        x"ca", x"b5", x"b1", x"b9", x"c3", x"cf", x"db", x"e6", x"ef", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f0", x"ee", x"c1", x"64", x"35", 
        x"2b", x"24", x"1e", x"1d", x"23", x"2d", x"38", x"43", x"4a", x"50", x"5f", x"72", x"8b", x"a1", x"b3", 
        x"b6", x"b0", x"ab", x"a9", x"a9", x"a9", x"a9", x"aa", x"ad", x"b1", x"b3", x"b0", x"b1", x"b1", x"b2", 
        x"b6", x"b4", x"bb", x"96", x"58", x"3a", x"71", x"8f", x"b6", x"b3", x"b3", x"b6", x"b6", x"b5", x"b3", 
        x"b2", x"b2", x"b3", x"b3", x"b2", x"af", x"ad", x"aa", x"a8", x"a6", x"a2", x"9c", x"9b", x"9e", x"9b", 
        x"97", x"9d", x"a8", x"b8", x"cc", x"e0", x"e7", x"f1", x"ee", x"ef", x"ee", x"ed", x"eb", x"e9", x"eb", 
        x"ef", x"ee", x"ed", x"ee", x"ec", x"e4", x"da", x"cb", x"b6", x"9f", x"8d", x"80", x"73", x"75", x"81", 
        x"8b", x"a1", x"aa", x"b1", x"b7", x"b7", x"b3", x"b5", x"bf", x"c1", x"c6", x"ca", x"cd", x"cf", x"cb", 
        x"cd", x"d2", x"d2", x"d2", x"d5", x"d6", x"cd", x"cc", x"d2", x"d1", x"d2", x"d1", x"cd", x"cb", x"ca", 
        x"d0", x"d1", x"d1", x"d0", x"d0", x"cb", x"c9", x"d0", x"d1", x"d4", x"d2", x"d6", x"b3", x"3c", x"25", 
        x"16", x"39", x"63", x"73", x"84", x"8a", x"8a", x"87", x"81", x"7d", x"79", x"75", x"73", x"77", x"79", 
        x"9d", x"9c", x"9c", x"9b", x"9b", x"9b", x"9a", x"9b", x"9b", x"9c", x"9c", x"9b", x"9b", x"9b", x"9b", 
        x"99", x"9a", x"9b", x"9b", x"9a", x"99", x"99", x"9b", x"9b", x"9b", x"9b", x"9c", x"9b", x"9a", x"99", 
        x"9a", x"9a", x"9a", x"9c", x"9c", x"9b", x"9b", x"9b", x"9b", x"9b", x"9b", x"9a", x"99", x"9a", x"9a", 
        x"9a", x"9a", x"9a", x"9a", x"9a", x"9c", x"9c", x"9c", x"9c", x"9b", x"9b", x"9a", x"99", x"9a", x"9a", 
        x"9d", x"9d", x"9b", x"9b", x"9d", x"9c", x"9c", x"9c", x"9c", x"9c", x"9b", x"9b", x"9c", x"9d", x"9b", 
        x"9c", x"9c", x"9b", x"9d", x"9f", x"9f", x"9e", x"9c", x"9b", x"9c", x"9c", x"9c", x"9c", x"9c", x"9b", 
        x"9d", x"9f", x"9e", x"9e", x"9d", x"9b", x"9e", x"9e", x"9c", x"9d", x"9e", x"9d", x"9d", x"9e", x"9d", 
        x"9e", x"a1", x"8a", x"74", x"89", x"81", x"8a", x"8b", x"89", x"88", x"89", x"88", x"8a", x"8a", x"8a", 
        x"8a", x"8b", x"8c", x"8b", x"87", x"92", x"65", x"41", x"58", x"4a", x"44", x"65", x"8f", x"8d", x"8e", 
        x"8e", x"8d", x"8c", x"8a", x"8b", x"8d", x"8c", x"84", x"4e", x"3b", x"3e", x"54", x"89", x"74", x"70", 
        x"6a", x"6d", x"c7", x"de", x"d6", x"d6", x"d8", x"da", x"df", x"d2", x"d3", x"d3", x"d2", x"d5", x"d4", 
        x"d5", x"d6", x"d4", x"d3", x"d3", x"d3", x"d5", x"d3", x"d4", x"d4", x"d3", x"d1", x"d2", x"d6", x"d6", 
        x"d4", x"d3", x"d2", x"d1", x"d1", x"d3", x"d4", x"d3", x"d3", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", 
        x"d3", x"d4", x"d3", x"d2", x"d3", x"d5", x"d4", x"d0", x"d2", x"d7", x"d5", x"d2", x"d1", x"d3", x"d4", 
        x"d5", x"d5", x"ee", x"ef", x"ed", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"ef", x"f0", x"e9", x"ec", x"f2", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f0", x"f1", x"f2", x"f2", x"f3", x"f4", x"f3", x"f4", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f5", x"f5", x"f3", x"ee", x"e2", x"cd", x"b7", x"9c", x"7e", x"66", 
        x"51", x"34", x"13", x"08", x"0e", x"15", x"1b", x"26", x"2c", x"23", x"1d", x"1d", x"23", x"2d", x"38", 
        x"34", x"40", x"78", x"c0", x"81", x"49", x"4f", x"a1", x"df", x"da", x"de", x"e0", x"f1", x"f4", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", 
        x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f2", x"f0", x"f0", x"f5", x"f5", x"f3", x"f2", x"f3", x"f3", x"f2", x"f1", x"f5", 
        x"f9", x"f6", x"eb", x"dc", x"cb", x"bd", x"b4", x"b0", x"b5", x"c6", x"da", x"eb", x"f2", x"f5", x"f3", 
        x"f1", x"f0", x"f2", x"f3", x"f2", x"f3", x"f1", x"f0", x"f3", x"f4", x"f2", x"f0", x"f0", x"a5", x"2c", 
        x"11", x"27", x"2f", x"3a", x"4d", x"5c", x"68", x"7d", x"92", x"a2", x"ad", x"b0", x"ab", x"a8", x"a6", 
        x"a5", x"a4", x"a4", x"a5", x"a9", x"ab", x"ac", x"af", x"b1", x"b2", x"b3", x"b4", x"b3", x"b1", x"b0", 
        x"b1", x"b1", x"ba", x"9b", x"5b", x"3d", x"6a", x"89", x"b3", x"b7", x"b7", x"b7", x"b8", x"b8", x"b7", 
        x"b3", x"ae", x"ab", x"a7", x"a4", x"a1", x"9e", x"9c", x"9d", x"9e", x"9e", x"9f", x"9e", x"9f", x"98", 
        x"b0", x"df", x"ef", x"f2", x"ee", x"ed", x"ee", x"eb", x"eb", x"ec", x"ed", x"f1", x"f1", x"f1", x"ef", 
        x"e5", x"d7", x"c6", x"b2", x"9c", x"8b", x"85", x"83", x"80", x"83", x"8f", x"9f", x"ab", x"b0", x"b3", 
        x"b4", x"bc", x"bd", x"bc", x"be", x"c3", x"c8", x"cf", x"d3", x"d2", x"ce", x"cc", x"cb", x"cf", x"d4", 
        x"d7", x"d8", x"d4", x"cf", x"cd", x"ce", x"d0", x"d2", x"d5", x"d1", x"cc", x"cb", x"cc", x"d0", x"d1", 
        x"d2", x"d1", x"ce", x"cc", x"cc", x"ce", x"d1", x"d5", x"d0", x"ce", x"cd", x"d1", x"b7", x"43", x"25", 
        x"16", x"37", x"64", x"73", x"81", x"8d", x"8b", x"87", x"86", x"86", x"84", x"7e", x"7a", x"78", x"74", 
        x"9c", x"9d", x"9d", x"9d", x"9d", x"9c", x"9b", x"9b", x"9b", x"9b", x"9a", x"9a", x"9a", x"9a", x"9a", 
        x"9b", x"9b", x"9b", x"9a", x"99", x"99", x"99", x"9b", x"9c", x"9b", x"9b", x"9c", x"9b", x"9a", x"99", 
        x"9a", x"9b", x"9c", x"9c", x"9a", x"99", x"9b", x"9b", x"9b", x"9a", x"99", x"99", x"9a", x"9b", x"9b", 
        x"9a", x"9a", x"9a", x"9b", x"9b", x"9c", x"9b", x"9a", x"9b", x"9c", x"9c", x"9a", x"99", x"9b", x"9d", 
        x"9d", x"9d", x"9c", x"9b", x"9c", x"9d", x"9c", x"9b", x"9a", x"9b", x"9c", x"9c", x"9d", x"9f", x"9c", 
        x"9d", x"9d", x"9c", x"9e", x"9d", x"9d", x"9e", x"9d", x"9b", x"9c", x"9d", x"9c", x"9e", x"9d", x"9b", 
        x"9c", x"9e", x"9e", x"9e", x"9d", x"9c", x"9d", x"9d", x"9c", x"9c", x"9e", x"9e", x"9f", x"9f", x"9d", 
        x"a0", x"a2", x"8b", x"72", x"88", x"7f", x"89", x"8e", x"8b", x"8b", x"8b", x"8c", x"8c", x"8a", x"8b", 
        x"8b", x"8e", x"8e", x"8d", x"89", x"92", x"63", x"3b", x"53", x"48", x"45", x"65", x"90", x"8e", x"8d", 
        x"89", x"8d", x"8e", x"88", x"8b", x"8f", x"8d", x"83", x"4e", x"3c", x"3d", x"53", x"8c", x"7a", x"77", 
        x"71", x"75", x"cc", x"df", x"d6", x"d8", x"d8", x"d9", x"df", x"d2", x"d3", x"d3", x"d4", x"d4", x"d4", 
        x"d5", x"d6", x"d4", x"d4", x"d3", x"d4", x"d6", x"d4", x"d4", x"d3", x"d3", x"d2", x"d3", x"d5", x"d5", 
        x"d4", x"d5", x"d4", x"d1", x"d1", x"d4", x"d4", x"d2", x"d3", x"d4", x"d2", x"d1", x"d1", x"d2", x"d2", 
        x"d2", x"d3", x"d2", x"d1", x"d3", x"d5", x"d4", x"d1", x"d1", x"d7", x"d5", x"d2", x"d5", x"d4", x"d4", 
        x"d4", x"d3", x"ed", x"ef", x"ef", x"ee", x"ed", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"f2", x"ef", x"f0", x"ea", x"eb", x"f3", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f4", x"f4", x"f4", x"f3", x"ee", x"e3", x"d0", 
        x"bc", x"a3", x"82", x"66", x"50", x"3b", x"31", x"36", x"40", x"44", x"48", x"4c", x"4e", x"56", x"59", 
        x"62", x"88", x"b3", x"c2", x"81", x"4b", x"4e", x"9e", x"e0", x"dc", x"de", x"e1", x"f2", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f4", x"f5", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f2", x"f3", x"f4", x"f3", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", 
        x"f1", x"f1", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f5", x"f2", x"f2", x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f4", 
        x"f7", x"f7", x"f6", x"f7", x"f4", x"eb", x"df", x"d1", x"c1", x"b5", x"b0", x"b5", x"c0", x"d2", x"e3", 
        x"ef", x"f1", x"f2", x"f3", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"ef", x"ef", x"f4", x"d2", x"5a", 
        x"25", x"22", x"45", x"6b", x"80", x"91", x"9c", x"a2", x"a1", x"a1", x"a1", x"a0", x"9d", x"a0", x"a3", 
        x"a4", x"a5", x"a6", x"a8", x"aa", x"ad", x"ad", x"af", x"b1", x"b2", x"b4", x"b5", x"b3", x"b3", x"b2", 
        x"b3", x"b4", x"bc", x"9d", x"5e", x"3e", x"65", x"8d", x"b8", x"b8", x"ba", x"ba", x"b4", x"ae", x"a9", 
        x"a6", x"a3", x"a0", x"9d", x"9d", x"9d", x"9c", x"9d", x"9e", x"9f", x"9b", x"9c", x"9c", x"a1", x"95", 
        x"af", x"eb", x"f0", x"ed", x"ea", x"ec", x"ef", x"eb", x"ed", x"ed", x"eb", x"e1", x"d3", x"c3", x"af", 
        x"98", x"8c", x"88", x"84", x"84", x"8e", x"a0", x"aa", x"ae", x"b2", x"b5", x"b9", x"c0", x"c3", x"c1", 
        x"c1", x"c5", x"c7", x"cb", x"d2", x"d5", x"d1", x"cc", x"ce", x"d2", x"d3", x"d4", x"d6", x"d3", x"d1", 
        x"d0", x"cf", x"d2", x"d8", x"d8", x"d4", x"d0", x"d0", x"d4", x"d2", x"d0", x"d4", x"d1", x"cd", x"cb", 
        x"d0", x"d1", x"d3", x"d3", x"d0", x"d0", x"cd", x"cf", x"ce", x"cf", x"d2", x"d6", x"bd", x"48", x"1e", 
        x"13", x"31", x"60", x"74", x"81", x"90", x"90", x"8b", x"88", x"87", x"84", x"81", x"81", x"81", x"7a", 
        x"99", x"9c", x"9d", x"9e", x"9c", x"9c", x"9c", x"9b", x"9a", x"9a", x"9a", x"99", x"99", x"9a", x"9a", 
        x"9a", x"9a", x"9b", x"9b", x"9b", x"9b", x"98", x"99", x"9c", x"9c", x"9b", x"9c", x"9a", x"97", x"99", 
        x"9b", x"9c", x"9c", x"9b", x"9a", x"99", x"9a", x"9c", x"9b", x"9a", x"99", x"99", x"9a", x"9b", x"9b", 
        x"9b", x"9a", x"9a", x"9b", x"9b", x"9c", x"9a", x"99", x"99", x"9a", x"9c", x"9c", x"9b", x"9b", x"9c", 
        x"9d", x"9c", x"9b", x"9c", x"9c", x"9c", x"9c", x"9b", x"9b", x"9c", x"9c", x"9d", x"9e", x"9f", x"9d", 
        x"9e", x"a0", x"9e", x"9e", x"9a", x"9a", x"9d", x"9d", x"9d", x"9d", x"9e", x"9e", x"9f", x"9f", x"9d", 
        x"9d", x"9f", x"9f", x"9e", x"9d", x"9c", x"9d", x"9d", x"9c", x"9d", x"9e", x"9d", x"9e", x"9e", x"9c", 
        x"9f", x"a2", x"8b", x"73", x"87", x"7e", x"88", x"8c", x"89", x"8a", x"8b", x"8c", x"8d", x"8b", x"8c", 
        x"8d", x"8f", x"8c", x"8b", x"8b", x"95", x"62", x"3a", x"55", x"4c", x"44", x"63", x"91", x"8f", x"90", 
        x"8c", x"8c", x"8f", x"8a", x"8b", x"8c", x"90", x"86", x"4e", x"3b", x"3f", x"57", x"92", x"84", x"76", 
        x"5c", x"53", x"c0", x"de", x"d7", x"d8", x"d5", x"d8", x"df", x"d3", x"d3", x"d2", x"d3", x"d4", x"d5", 
        x"d4", x"d6", x"d4", x"d4", x"d3", x"d4", x"d7", x"d4", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", 
        x"d4", x"d4", x"d4", x"d4", x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", x"d1", x"d1", x"d1", x"d2", x"d3", 
        x"d3", x"d3", x"d2", x"d2", x"d3", x"d4", x"d3", x"d0", x"d1", x"d9", x"d7", x"d2", x"d5", x"d4", x"d4", 
        x"d6", x"d5", x"ea", x"ec", x"ee", x"ef", x"ed", x"ee", x"ed", x"ec", x"ed", x"ee", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ed", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"f2", x"f0", x"f0", x"ea", x"ea", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f5", x"f5", x"f3", 
        x"f4", x"f5", x"ed", x"dd", x"cc", x"b3", x"94", x"79", x"62", x"4f", x"4c", x"52", x"63", x"6e", x"78", 
        x"a2", x"ba", x"bc", x"c1", x"86", x"4e", x"4d", x"9a", x"df", x"e0", x"e1", x"df", x"f1", x"f3", x"f2", 
        x"f4", x"f3", x"f2", x"f5", x"f5", x"f5", x"f4", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f1", x"f2", x"f6", x"f3", x"f1", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f6", 
        x"f7", x"f6", x"f6", x"f6", x"f5", x"f2", x"f3", x"f2", x"ef", x"e7", x"d8", x"c6", x"ba", x"ac", x"ab", 
        x"b6", x"cc", x"e3", x"f2", x"f5", x"f1", x"f0", x"f0", x"f1", x"f3", x"f3", x"ee", x"ef", x"ea", x"8c", 
        x"3e", x"1e", x"60", x"94", x"8a", x"8f", x"91", x"91", x"92", x"96", x"98", x"98", x"9b", x"9b", x"9e", 
        x"a2", x"a6", x"a8", x"a9", x"ab", x"ae", x"ad", x"ae", x"b1", x"b2", x"b6", x"b7", x"b4", x"b2", x"b1", 
        x"b4", x"b5", x"bd", x"a4", x"63", x"3f", x"64", x"8f", x"b3", x"ad", x"a9", x"a7", x"a3", x"a0", x"9f", 
        x"a0", x"a1", x"a1", x"9f", x"9f", x"9e", x"9d", x"9c", x"9d", x"9f", x"9e", x"9d", x"9b", x"9f", x"92", 
        x"a5", x"e7", x"f1", x"f0", x"f3", x"f3", x"ed", x"e1", x"c9", x"b0", x"a0", x"92", x"86", x"82", x"85", 
        x"8c", x"9a", x"a8", x"ae", x"af", x"b0", x"b6", x"bd", x"c1", x"c7", x"c8", x"c6", x"c7", x"ca", x"cf", 
        x"d6", x"d7", x"d2", x"cb", x"c8", x"cc", x"d2", x"d7", x"d9", x"d7", x"ce", x"ca", x"cf", x"d3", x"d7", 
        x"d7", x"d3", x"d1", x"d2", x"d3", x"d6", x"da", x"da", x"d8", x"ce", x"c8", x"cd", x"d1", x"d4", x"d6", 
        x"d7", x"d1", x"cd", x"cd", x"cf", x"d3", x"d4", x"d6", x"d0", x"cb", x"cc", x"d1", x"be", x"4f", x"20", 
        x"15", x"2e", x"5c", x"74", x"83", x"92", x"92", x"8d", x"88", x"87", x"85", x"82", x"82", x"80", x"81", 
        x"98", x"9c", x"9f", x"9e", x"9c", x"9b", x"9b", x"9a", x"9a", x"9a", x"9a", x"9a", x"9b", x"9c", x"9b", 
        x"9a", x"9b", x"9b", x"9c", x"9c", x"9c", x"9b", x"9b", x"9c", x"9a", x"9a", x"9c", x"9c", x"99", x"99", 
        x"9b", x"9c", x"9c", x"9a", x"9a", x"9a", x"9b", x"9d", x"9e", x"9d", x"9b", x"9b", x"9b", x"9c", x"9c", 
        x"9b", x"9b", x"9b", x"9c", x"9c", x"9c", x"9b", x"9a", x"99", x"9a", x"9c", x"9e", x"9c", x"9b", x"9c", 
        x"9d", x"9c", x"9c", x"9e", x"9d", x"9a", x"9c", x"9e", x"9e", x"9e", x"9c", x"9b", x"9e", x"9e", x"9d", 
        x"9e", x"a0", x"9f", x"9e", x"9c", x"9c", x"9d", x"9e", x"9d", x"9d", x"9d", x"9f", x"a0", x"9f", x"9e", 
        x"9e", x"9e", x"9e", x"9e", x"9e", x"9d", x"9d", x"9d", x"9d", x"9e", x"9e", x"9d", x"9e", x"9e", x"9d", 
        x"a0", x"a1", x"89", x"6e", x"85", x"7e", x"88", x"8b", x"8a", x"8c", x"8b", x"8b", x"8c", x"8b", x"8c", 
        x"8c", x"8d", x"8a", x"88", x"8a", x"94", x"64", x"3c", x"56", x"4b", x"40", x"62", x"94", x"91", x"92", 
        x"90", x"8d", x"8d", x"89", x"8d", x"8c", x"8d", x"86", x"52", x"3a", x"42", x"5a", x"79", x"51", x"32", 
        x"1f", x"3b", x"c1", x"e5", x"d9", x"d8", x"d5", x"da", x"e0", x"d3", x"d3", x"d1", x"d2", x"d4", x"d5", 
        x"d4", x"d6", x"d4", x"d4", x"d3", x"d4", x"d6", x"d4", x"d3", x"d3", x"d3", x"d5", x"d5", x"d4", x"d4", 
        x"d5", x"d4", x"d4", x"d5", x"d5", x"d4", x"d1", x"d2", x"d2", x"d1", x"d1", x"d1", x"d1", x"d2", x"d4", 
        x"d4", x"d3", x"d2", x"d2", x"d1", x"d2", x"d2", x"cd", x"ce", x"d8", x"d6", x"d1", x"d5", x"d7", x"d4", 
        x"d4", x"d6", x"ed", x"f0", x"ed", x"ee", x"ef", x"ef", x"ee", x"ed", x"ec", x"ed", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f1", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ee", 
        x"ee", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f2", x"f1", x"f0", x"e9", x"ea", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f0", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f4", 
        x"f1", x"f0", x"f3", x"f4", x"f5", x"f5", x"ee", x"e1", x"d4", x"c2", x"a6", x"8c", x"72", x"68", x"83", 
        x"ad", x"b5", x"be", x"c8", x"92", x"50", x"4e", x"9c", x"e2", x"e1", x"df", x"e0", x"f3", x"f5", x"f2", 
        x"f5", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f4", x"f2", x"f2", x"f6", x"f4", x"f1", x"f2", x"f3", x"f1", x"f1", x"f2", x"f4", x"f4", x"f4", x"f6", 
        x"f6", x"f7", x"f7", x"f5", x"f4", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"ee", x"eb", x"e2", x"d4", 
        x"c4", x"b6", x"ad", x"b3", x"c4", x"d8", x"e7", x"ef", x"f2", x"f0", x"ee", x"ed", x"ed", x"f1", x"a8", 
        x"51", x"2e", x"5a", x"92", x"8b", x"8b", x"8a", x"87", x"88", x"8e", x"91", x"92", x"97", x"9a", x"9e", 
        x"a3", x"a7", x"a8", x"a9", x"ab", x"af", x"ae", x"af", x"b1", x"b0", x"b4", x"b7", x"b7", x"b7", x"b8", 
        x"ba", x"b9", x"bd", x"a5", x"65", x"40", x"5f", x"86", x"a0", x"9e", x"9f", x"a2", x"a2", x"a1", x"a1", 
        x"a0", x"9f", x"9f", x"9e", x"9f", x"9f", x"9e", x"9d", x"9e", x"9f", x"9d", x"9c", x"9b", x"9c", x"95", 
        x"a6", x"dc", x"e1", x"d0", x"b6", x"92", x"82", x"87", x"81", x"80", x"89", x"9a", x"a9", x"b1", x"b2", 
        x"b1", x"b4", x"ba", x"c4", x"c8", x"c9", x"ca", x"ca", x"cb", x"d1", x"d4", x"d5", x"d6", x"d3", x"cf", 
        x"ce", x"cd", x"d3", x"d7", x"d6", x"d1", x"cd", x"ca", x"ce", x"d6", x"d9", x"d8", x"d6", x"d1", x"d0", 
        x"d4", x"d7", x"da", x"d9", x"d4", x"ce", x"ca", x"ca", x"d4", x"d5", x"d6", x"d7", x"d2", x"cd", x"cd", 
        x"d5", x"d6", x"d9", x"d8", x"d2", x"cb", x"c7", x"d1", x"d5", x"d8", x"d9", x"d9", x"c2", x"53", x"22", 
        x"18", x"2d", x"59", x"73", x"7f", x"91", x"91", x"8c", x"89", x"88", x"86", x"84", x"82", x"82", x"7f", 
        x"9a", x"9e", x"9f", x"9e", x"9b", x"9a", x"9b", x"9c", x"9c", x"9c", x"9b", x"9b", x"9b", x"9b", x"9a", 
        x"9a", x"9b", x"9c", x"9d", x"9d", x"9d", x"9d", x"9d", x"9c", x"99", x"98", x"9b", x"9d", x"9b", x"9a", 
        x"9c", x"9c", x"9c", x"9b", x"9b", x"9b", x"9d", x"9d", x"9e", x"9d", x"9b", x"9b", x"9c", x"9d", x"9c", 
        x"9c", x"9b", x"9b", x"9c", x"9d", x"9d", x"9d", x"9c", x"9b", x"9b", x"9b", x"9c", x"9b", x"9b", x"9c", 
        x"9c", x"9c", x"9c", x"9e", x"9e", x"9c", x"9c", x"9c", x"9c", x"9d", x"9d", x"9d", x"9d", x"9c", x"9c", 
        x"9d", x"9e", x"9e", x"9d", x"9f", x"9f", x"9e", x"9e", x"9e", x"9e", x"9d", x"9f", x"9f", x"9e", x"9e", 
        x"9d", x"9d", x"9d", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9f", x"9e", x"9d", x"9e", x"9e", x"9d", 
        x"a0", x"a2", x"86", x"66", x"7f", x"78", x"80", x"84", x"87", x"8b", x"88", x"88", x"89", x"8a", x"8c", 
        x"8c", x"8d", x"8d", x"89", x"89", x"90", x"63", x"3d", x"54", x"48", x"3d", x"61", x"94", x"90", x"91", 
        x"92", x"92", x"92", x"8b", x"8d", x"8f", x"94", x"86", x"51", x"3c", x"3d", x"34", x"31", x"22", x"1c", 
        x"11", x"38", x"be", x"dd", x"d5", x"da", x"d8", x"d9", x"df", x"d3", x"d3", x"d1", x"d0", x"d3", x"d5", 
        x"d4", x"d5", x"d4", x"d5", x"d3", x"d3", x"d5", x"d4", x"d3", x"d3", x"d3", x"d5", x"d5", x"d4", x"d4", 
        x"d6", x"d4", x"d3", x"d4", x"d5", x"d4", x"d2", x"d3", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d4", 
        x"d4", x"d3", x"d3", x"d2", x"d1", x"d0", x"d3", x"ce", x"ce", x"d7", x"d6", x"d1", x"d6", x"d6", x"d3", 
        x"d3", x"d5", x"e8", x"ef", x"ee", x"ed", x"ed", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"ee", x"ed", x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", 
        x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f0", x"e9", x"ea", x"f1", 
        x"f3", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f3", x"f0", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f5", x"f5", x"f4", x"f1", x"f0", 
        x"f2", x"f4", x"f3", x"f2", x"f1", x"f3", x"f4", x"f3", x"f3", x"f3", x"ed", x"e4", x"d8", x"cb", x"ba", 
        x"9f", x"93", x"96", x"a2", x"7b", x"4d", x"47", x"96", x"e2", x"e6", x"e6", x"e3", x"f0", x"f0", x"ee", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f5", x"f3", x"f3", x"f7", x"f5", x"f1", x"f1", x"f2", x"f1", x"f1", x"f3", x"f5", x"f6", x"f6", x"f6", 
        x"f7", x"f8", x"f7", x"f4", x"f2", x"f2", x"f3", x"f2", x"f1", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", 
        x"ee", x"e8", x"e1", x"cf", x"b9", x"a8", x"ab", x"b9", x"cd", x"df", x"ea", x"ef", x"f2", x"f2", x"b3", 
        x"56", x"4b", x"5a", x"96", x"92", x"91", x"91", x"8e", x"8b", x"8e", x"92", x"95", x"97", x"9d", x"a2", 
        x"a4", x"a5", x"a8", x"ab", x"ad", x"b1", x"b1", x"b3", x"b5", x"b5", x"b8", x"bd", x"bd", x"ba", x"b3", 
        x"b0", x"aa", x"a9", x"9c", x"65", x"41", x"5c", x"84", x"99", x"9f", x"a0", x"a0", x"a0", x"9f", x"9f", 
        x"9f", x"9e", x"9f", x"9f", x"9f", x"9e", x"9c", x"9b", x"9c", x"9c", x"9d", x"9a", x"9c", x"9a", x"98", 
        x"9c", x"a9", x"95", x"7a", x"5f", x"39", x"46", x"8e", x"b0", x"b5", x"b7", x"b9", x"bb", x"bf", x"c3", 
        x"c4", x"c9", x"cf", x"ce", x"cc", x"cf", x"d6", x"d8", x"d7", x"d6", x"d1", x"ce", x"d3", x"d7", x"d6", 
        x"d5", x"d2", x"d1", x"d0", x"d3", x"d7", x"da", x"d9", x"d6", x"d7", x"d3", x"d3", x"d8", x"d9", x"da", 
        x"d5", x"ce", x"ca", x"cd", x"d3", x"d9", x"d9", x"d4", x"d3", x"cf", x"cf", x"d5", x"d7", x"d4", x"d4", 
        x"d6", x"d3", x"d2", x"d3", x"d3", x"d3", x"d1", x"d3", x"d2", x"cf", x"d1", x"d5", x"c9", x"64", x"23", 
        x"18", x"29", x"59", x"78", x"80", x"91", x"94", x"92", x"8f", x"8d", x"8b", x"89", x"87", x"86", x"82", 
        x"9d", x"9e", x"9f", x"9d", x"9b", x"9b", x"9b", x"9c", x"9c", x"9c", x"9b", x"9c", x"9c", x"9c", x"9b", 
        x"99", x"9a", x"9b", x"9c", x"9c", x"9c", x"9c", x"9a", x"9a", x"9a", x"9a", x"9a", x"9a", x"9b", x"9b", 
        x"9b", x"9c", x"9b", x"9b", x"9b", x"9c", x"9f", x"9e", x"9b", x"9a", x"9b", x"9c", x"9d", x"9d", x"9d", 
        x"9c", x"9c", x"9c", x"9d", x"9d", x"9d", x"9d", x"9e", x"9d", x"9c", x"9c", x"9c", x"9b", x"9b", x"9d", 
        x"9d", x"9d", x"9d", x"9e", x"9e", x"9c", x"9d", x"9d", x"9d", x"9d", x"9d", x"9d", x"9c", x"9b", x"9d", 
        x"9d", x"9c", x"9e", x"9c", x"9f", x"9e", x"9d", x"9d", x"9f", x"a0", x"a0", x"a0", x"9e", x"9d", x"9e", 
        x"9d", x"9d", x"9e", x"9e", x"9f", x"a0", x"9f", x"9f", x"a0", x"9f", x"9e", x"9d", x"9e", x"9f", x"9d", 
        x"a0", x"a2", x"89", x"70", x"97", x"97", x"9f", x"9f", x"9b", x"99", x"93", x"91", x"91", x"8f", x"8f", 
        x"8d", x"8b", x"8c", x"8a", x"89", x"91", x"63", x"36", x"4c", x"46", x"41", x"66", x"99", x"99", x"99", 
        x"96", x"91", x"8e", x"8a", x"8f", x"95", x"96", x"7b", x"46", x"26", x"22", x"1c", x"19", x"0f", x"09", 
        x"06", x"37", x"c1", x"e1", x"d9", x"da", x"d6", x"d7", x"de", x"d3", x"d3", x"d1", x"d0", x"d3", x"d5", 
        x"d3", x"d5", x"d4", x"d5", x"d3", x"d2", x"d4", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"d5", 
        x"d6", x"d4", x"d4", x"d5", x"d5", x"d4", x"d3", x"d4", x"d2", x"d0", x"d0", x"d1", x"d2", x"d2", x"d4", 
        x"d4", x"d3", x"d3", x"d3", x"d1", x"d0", x"d5", x"cf", x"cf", x"d7", x"d7", x"d3", x"d6", x"d3", x"d1", 
        x"d3", x"d5", x"e7", x"ef", x"ee", x"ec", x"ec", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ed", x"ec", x"ec", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f2", x"ef", x"ea", x"eb", x"f1", 
        x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f0", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f0", x"ef", 
        x"f2", x"f4", x"f3", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f4", x"f4", x"f5", x"f1", x"f1", x"ee", 
        x"e4", x"de", x"d2", x"ba", x"9c", x"7c", x"5d", x"97", x"e0", x"e6", x"e3", x"e1", x"ea", x"f2", x"f3", 
        x"f6", x"f3", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f5", x"f5", x"f4", x"f7", x"f5", x"f1", x"f1", x"f3", x"f2", x"f2", x"f4", x"f6", x"f6", x"f6", x"f6", 
        x"f8", x"f9", x"f6", x"f4", x"f2", x"f1", x"f2", x"f1", x"ef", x"f0", x"f2", x"f2", x"ef", x"ee", x"f3", 
        x"f5", x"f0", x"ee", x"ef", x"ed", x"e4", x"d3", x"bc", x"ab", x"a6", x"b2", x"c7", x"da", x"e4", x"b6", 
        x"55", x"58", x"5c", x"9d", x"95", x"93", x"96", x"92", x"8e", x"90", x"96", x"99", x"9c", x"a0", x"a5", 
        x"a5", x"a5", x"aa", x"af", x"b0", x"b4", x"b5", x"b8", x"b9", x"b4", x"b1", x"af", x"ad", x"a8", x"a0", 
        x"9f", x"9f", x"a2", x"9c", x"66", x"41", x"58", x"84", x"97", x"9f", x"9d", x"9c", x"9e", x"9f", x"9e", 
        x"9c", x"9a", x"99", x"9a", x"9b", x"9b", x"9a", x"9a", x"9a", x"9b", x"99", x"98", x"9a", x"97", x"98", 
        x"95", x"8d", x"91", x"95", x"82", x"52", x"64", x"b0", x"c2", x"c1", x"c5", x"ca", x"d0", x"d3", x"d4", 
        x"d1", x"d1", x"d6", x"d8", x"d8", x"d7", x"d5", x"d1", x"cf", x"d7", x"db", x"da", x"d6", x"d2", x"d1", 
        x"d5", x"d7", x"d9", x"d9", x"d6", x"d3", x"d2", x"d4", x"dc", x"df", x"d8", x"d3", x"d1", x"ce", x"ce", 
        x"d4", x"d7", x"d6", x"d3", x"d2", x"d2", x"d3", x"d5", x"da", x"d6", x"d1", x"d1", x"cf", x"cd", x"d1", 
        x"dc", x"da", x"d7", x"d4", x"cf", x"cd", x"cc", x"d7", x"d9", x"d7", x"d7", x"d7", x"cc", x"6a", x"24", 
        x"16", x"25", x"5a", x"7d", x"83", x"95", x"94", x"91", x"8e", x"8c", x"8b", x"8a", x"87", x"89", x"89", 
        x"9f", x"9e", x"9e", x"9d", x"9c", x"9c", x"9d", x"9c", x"9b", x"9b", x"9b", x"9b", x"9c", x"9d", x"9b", 
        x"9a", x"9b", x"9b", x"9c", x"9c", x"9c", x"9c", x"9a", x"99", x"9c", x"9d", x"99", x"99", x"9c", x"9c", 
        x"9b", x"9b", x"9b", x"9c", x"9c", x"9c", x"9f", x"9d", x"9b", x"9c", x"9d", x"9c", x"9b", x"9d", x"9e", 
        x"9d", x"9d", x"9d", x"9d", x"9d", x"9c", x"9c", x"9d", x"9d", x"9c", x"9c", x"9d", x"9c", x"9c", x"9e", 
        x"9f", x"9e", x"9d", x"9c", x"9d", x"9d", x"9e", x"9e", x"9e", x"9d", x"9c", x"9c", x"9c", x"9c", x"9f", 
        x"9d", x"9c", x"9f", x"9d", x"9c", x"9c", x"9c", x"9e", x"a0", x"a0", x"9f", x"9f", x"9d", x"9d", x"9f", 
        x"9f", x"9e", x"9f", x"9e", x"9f", x"a1", x"a0", x"a0", x"a1", x"9f", x"9e", x"9e", x"a0", x"a0", x"9e", 
        x"a1", x"a3", x"8b", x"77", x"a4", x"a3", x"a9", x"ac", x"ad", x"ae", x"ab", x"a7", x"a6", x"a2", x"a0", 
        x"9b", x"98", x"97", x"92", x"8c", x"93", x"66", x"3d", x"66", x"70", x"6a", x"7c", x"9f", x"9c", x"9b", 
        x"92", x"92", x"92", x"93", x"8f", x"7a", x"56", x"33", x"20", x"1a", x"13", x"0c", x"07", x"05", x"06", 
        x"07", x"36", x"bf", x"e2", x"d8", x"d5", x"d5", x"da", x"dd", x"d2", x"d4", x"d2", x"d0", x"d2", x"d4", 
        x"d2", x"d4", x"d4", x"d5", x"d3", x"d3", x"d4", x"d3", x"d4", x"d3", x"d3", x"d2", x"d3", x"d5", x"d6", 
        x"d5", x"d5", x"d6", x"d6", x"d5", x"d4", x"d3", x"d5", x"d2", x"d0", x"d0", x"d2", x"d3", x"d3", x"d3", 
        x"d2", x"d3", x"d3", x"d4", x"d2", x"d0", x"d3", x"cf", x"ce", x"d5", x"d6", x"d2", x"d3", x"d2", x"d5", 
        x"d6", x"d0", x"db", x"e9", x"ec", x"ee", x"f0", x"f1", x"f0", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ee", x"ed", x"ee", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ee", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"ef", x"eb", x"ec", x"f1", 
        x"f3", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f4", x"f3", x"f3", x"f4", x"f3", x"ef", x"f1", x"f1", x"f2", 
        x"f5", x"f0", x"f1", x"f2", x"ee", x"e9", x"d6", x"dd", x"e9", x"e7", x"e6", x"d6", x"d3", x"de", x"e5", 
        x"eb", x"f1", x"f4", x"f5", x"f5", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f2", x"f2", x"f3", x"f4", x"f4", x"f5", x"f5", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f6", x"f6", x"f4", x"f6", x"f5", x"f1", x"f2", x"f4", x"f4", x"f5", x"f6", x"f7", x"f6", x"f6", x"f7", 
        x"fa", x"f7", x"f3", x"f3", x"f3", x"f1", x"f2", x"f2", x"f0", x"ef", x"f1", x"f3", x"f1", x"f3", x"ef", 
        x"ee", x"f0", x"f1", x"ef", x"f1", x"f2", x"f2", x"f2", x"ed", x"df", x"c6", x"ae", x"a2", x"ac", x"93", 
        x"4f", x"66", x"5f", x"9c", x"9e", x"9b", x"9b", x"96", x"91", x"92", x"95", x"99", x"9f", x"a2", x"a6", 
        x"a8", x"ab", x"b0", x"b2", x"b1", x"b1", x"ae", x"ad", x"ac", x"a3", x"9e", x"9d", x"a1", x"a2", x"9e", 
        x"9e", x"9d", x"9e", x"9b", x"67", x"42", x"55", x"86", x"97", x"9f", x"9b", x"9b", x"9b", x"9a", x"99", 
        x"99", x"9b", x"9a", x"96", x"97", x"98", x"97", x"97", x"98", x"9a", x"9a", x"9b", x"99", x"9a", x"99", 
        x"95", x"93", x"99", x"99", x"a2", x"6f", x"62", x"ba", x"d5", x"d4", x"d8", x"d9", x"d9", x"d7", x"d6", 
        x"dc", x"db", x"d6", x"d4", x"d3", x"d6", x"dc", x"db", x"d7", x"d6", x"d6", x"d5", x"d9", x"d9", x"d8", 
        x"d7", x"d2", x"d0", x"d1", x"d5", x"d9", x"d7", x"d2", x"ce", x"d2", x"d1", x"d2", x"d6", x"d7", x"d7", 
        x"d0", x"d2", x"d6", x"d7", x"d7", x"d8", x"d6", x"d2", x"d6", x"d3", x"d2", x"d7", x"d8", x"d7", x"d3", 
        x"d2", x"d1", x"d3", x"d6", x"d7", x"d8", x"d4", x"d3", x"d1", x"ce", x"d2", x"d8", x"d4", x"77", x"27", 
        x"17", x"23", x"56", x"7b", x"89", x"a6", x"99", x"94", x"94", x"92", x"90", x"8b", x"84", x"78", x"66", 
        x"9f", x"9d", x"9c", x"9c", x"9c", x"9d", x"9e", x"9d", x"9c", x"9b", x"9a", x"9a", x"9b", x"9b", x"9c", 
        x"9c", x"9c", x"9c", x"9d", x"9d", x"9c", x"9c", x"9c", x"9b", x"9d", x"9d", x"9a", x"9b", x"9e", x"9d", 
        x"9b", x"9c", x"9d", x"9d", x"9d", x"9c", x"9d", x"9c", x"9d", x"9e", x"9f", x"9e", x"9a", x"9c", x"9d", 
        x"9c", x"9c", x"9d", x"9d", x"9e", x"9e", x"9d", x"9d", x"9c", x"9c", x"9d", x"9e", x"9e", x"9e", x"9f", 
        x"9f", x"9e", x"9d", x"9c", x"9e", x"9f", x"9e", x"9c", x"9c", x"9d", x"9d", x"9d", x"9d", x"9d", x"a0", 
        x"9f", x"9d", x"9f", x"9e", x"9d", x"9d", x"9d", x"9e", x"a0", x"9f", x"9f", x"9f", x"9e", x"9e", x"9f", 
        x"9f", x"9e", x"9e", x"9d", x"9e", x"a0", x"a0", x"a0", x"a0", x"9e", x"9d", x"9f", x"9f", x"9f", x"9f", 
        x"a2", x"a3", x"8a", x"73", x"a4", x"a5", x"a9", x"a9", x"a8", x"a8", x"ab", x"aa", x"ab", x"ad", x"ae", 
        x"ac", x"ad", x"ad", x"a9", x"a9", x"b0", x"7a", x"44", x"6e", x"7b", x"75", x"87", x"ab", x"ab", x"a9", 
        x"97", x"90", x"85", x"6a", x"48", x"2a", x"1c", x"17", x"15", x"09", x"05", x"05", x"03", x"03", x"03", 
        x"08", x"39", x"bc", x"e1", x"d9", x"d9", x"d9", x"dc", x"dd", x"d2", x"d4", x"d2", x"d1", x"d2", x"d4", 
        x"d2", x"d3", x"d3", x"d4", x"d3", x"d3", x"d4", x"d4", x"d4", x"d4", x"d3", x"d2", x"d3", x"d5", x"d6", 
        x"d4", x"d5", x"d5", x"d7", x"d4", x"d2", x"d4", x"d5", x"d2", x"d1", x"d1", x"d2", x"d2", x"d1", x"d2", 
        x"d4", x"d3", x"d4", x"d4", x"d3", x"d2", x"cf", x"ce", x"cd", x"d5", x"d5", x"d2", x"d7", x"d4", x"cd", 
        x"c1", x"b2", x"b5", x"bd", x"c5", x"cf", x"d7", x"de", x"e6", x"eb", x"ef", x"f2", x"f2", x"f0", x"f0", 
        x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ed", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"f0", x"f1", 
        x"f0", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", x"ef", x"ec", x"eb", x"f0", 
        x"f1", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f0", x"f0", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f4", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f2", x"f1", 
        x"f0", x"f1", x"f3", x"f2", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f1", x"f0", x"f2", 
        x"f0", x"f3", x"f4", x"f5", x"f3", x"ee", x"f1", x"f4", x"f1", x"f3", x"ef", x"d9", x"ca", x"c5", x"c2", 
        x"c2", x"cd", x"d5", x"dc", x"e3", x"ed", x"f4", x"f6", x"f5", x"f4", x"f3", x"f2", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f2", 
        x"f3", x"f4", x"f3", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f5", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", 
        x"f4", x"f6", x"f4", x"f5", x"f4", x"f0", x"f0", x"f4", x"f4", x"f6", x"f7", x"f7", x"f5", x"f5", x"f8", 
        x"f9", x"f6", x"f2", x"f1", x"f2", x"f1", x"f0", x"f2", x"f2", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", 
        x"f2", x"f1", x"ef", x"ef", x"f1", x"f1", x"f2", x"f3", x"f1", x"f2", x"f2", x"ef", x"e6", x"d8", x"a0", 
        x"46", x"65", x"53", x"80", x"8a", x"91", x"98", x"9b", x"98", x"9a", x"9e", x"a0", x"a2", x"a5", x"a7", 
        x"a8", x"aa", x"a9", x"a6", x"a0", x"9f", x"9d", x"9d", x"9f", x"a1", x"9d", x"9b", x"9e", x"a1", x"9e", 
        x"9c", x"9b", x"9c", x"9d", x"6c", x"46", x"53", x"86", x"95", x"9d", x"99", x"99", x"9a", x"98", x"97", 
        x"97", x"98", x"99", x"97", x"97", x"96", x"95", x"95", x"95", x"96", x"97", x"98", x"95", x"98", x"97", 
        x"93", x"96", x"94", x"95", x"aa", x"77", x"5a", x"bb", x"df", x"da", x"dd", x"e0", x"e1", x"dd", x"d8", 
        x"d9", x"da", x"d9", x"da", x"d8", x"d6", x"d6", x"d5", x"d6", x"db", x"dd", x"dc", x"d8", x"d5", x"d0", 
        x"d2", x"d5", x"d7", x"d6", x"d3", x"d0", x"d0", x"d3", x"d4", x"da", x"db", x"d8", x"d6", x"d4", x"d6", 
        x"d5", x"d6", x"d7", x"d5", x"d5", x"d6", x"d5", x"d6", x"dd", x"da", x"d5", x"d4", x"d2", x"d1", x"d4", 
        x"d9", x"d9", x"d8", x"d3", x"cf", x"d1", x"d3", x"d7", x"da", x"d7", x"d5", x"d3", x"d1", x"7d", x"27", 
        x"18", x"21", x"52", x"7b", x"8d", x"ae", x"97", x"86", x"7a", x"67", x"54", x"47", x"3e", x"37", x"35", 
        x"9d", x"9d", x"9c", x"9b", x"9c", x"9c", x"9d", x"9d", x"9c", x"9b", x"9b", x"9c", x"9d", x"9c", x"9e", 
        x"9e", x"9c", x"9d", x"9e", x"9f", x"9d", x"9b", x"9b", x"9d", x"9d", x"9c", x"9b", x"9c", x"9d", x"9d", 
        x"9b", x"9d", x"9f", x"9e", x"9c", x"9c", x"9c", x"9c", x"9e", x"9b", x"9c", x"a0", x"9d", x"9c", x"9c", 
        x"9c", x"9c", x"9d", x"9e", x"9e", x"9f", x"9f", x"9e", x"9d", x"9c", x"9d", x"9e", x"9f", x"9f", x"9f", 
        x"9e", x"9d", x"9d", x"9d", x"9d", x"9d", x"9e", x"9d", x"9e", x"9d", x"9d", x"9d", x"9e", x"9e", x"9f", 
        x"9f", x"9f", x"9f", x"9e", x"9f", x"9f", x"9f", x"9e", x"9e", x"9f", x"a0", x"9f", x"9e", x"9e", x"9e", 
        x"9d", x"9c", x"9b", x"9c", x"9d", x"9e", x"a0", x"9f", x"9f", x"9d", x"9e", x"a0", x"a0", x"9e", x"a1", 
        x"a1", x"a1", x"8d", x"75", x"a4", x"a5", x"a7", x"a8", x"a8", x"a8", x"aa", x"aa", x"a8", x"aa", x"aa", 
        x"a6", x"a9", x"a9", x"a5", x"a7", x"b0", x"78", x"3e", x"68", x"72", x"6e", x"87", x"b0", x"ac", x"a0", 
        x"7c", x"5f", x"44", x"2f", x"20", x"19", x"11", x"08", x"06", x"05", x"04", x"05", x"0a", x"15", x"2e", 
        x"3f", x"49", x"c0", x"e4", x"d7", x"da", x"d8", x"da", x"df", x"d2", x"d3", x"d2", x"d2", x"d3", x"d4", 
        x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d5", x"d5", x"d4", x"d3", x"d3", x"d4", x"d5", x"d4", 
        x"d4", x"d4", x"d2", x"d6", x"d2", x"d0", x"d7", x"d5", x"d2", x"d2", x"d1", x"d0", x"d3", x"d3", x"d2", 
        x"d3", x"d3", x"d5", x"d5", x"d2", x"d2", x"cf", x"d1", x"cd", x"d6", x"db", x"d3", x"c7", x"b2", x"a7", 
        x"a0", x"aa", x"c7", x"c3", x"ba", x"b5", x"b4", x"b6", x"ba", x"c0", x"c9", x"d2", x"d9", x"e0", x"e7", 
        x"eb", x"ed", x"ef", x"f0", x"ef", x"ee", x"ed", x"ec", x"ed", x"ec", x"ec", x"eb", x"ee", x"ee", x"ee", 
        x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"ee", x"ee", x"f0", x"f1", x"f1", 
        x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"e8", x"f1", 
        x"f1", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"ef", x"ef", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f0", x"ef", x"ef", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f2", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f0", x"ed", x"ec", x"e4", 
        x"d7", x"cc", x"c4", x"be", x"c3", x"cc", x"d3", x"da", x"e4", x"ed", x"f3", x"f4", x"f3", x"f3", x"f4", 
        x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f3", x"f4", x"f3", x"f2", x"f1", 
        x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f4", x"f5", x"f4", x"f4", x"f0", x"ef", x"f4", x"f5", x"f6", x"f8", x"f8", x"f5", x"f5", x"f8", 
        x"f8", x"f5", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"ef", x"ef", x"f3", x"ce", 
        x"56", x"6e", x"57", x"78", x"73", x"76", x"7b", x"83", x"88", x"94", x"a0", x"a6", x"a2", x"a3", x"9f", 
        x"9b", x"9c", x"9b", x"97", x"96", x"99", x"9a", x"98", x"9c", x"a3", x"9a", x"98", x"98", x"9c", x"9d", 
        x"98", x"99", x"9a", x"9d", x"6c", x"47", x"4c", x"83", x"91", x"99", x"96", x"97", x"97", x"97", x"96", 
        x"95", x"96", x"96", x"94", x"93", x"94", x"95", x"96", x"95", x"94", x"94", x"95", x"94", x"93", x"92", 
        x"92", x"95", x"91", x"91", x"a7", x"89", x"5e", x"b5", x"e8", x"e0", x"dd", x"dc", x"dc", x"df", x"e1", 
        x"de", x"d9", x"d6", x"d6", x"d8", x"dc", x"dd", x"db", x"d9", x"d6", x"d7", x"d9", x"d9", x"dc", x"d6", 
        x"d4", x"d0", x"d2", x"d4", x"d7", x"d8", x"d7", x"d5", x"d4", x"d5", x"d7", x"d7", x"d7", x"d7", x"d8", 
        x"d5", x"d4", x"d8", x"d9", x"db", x"dc", x"dc", x"d8", x"d7", x"d7", x"d5", x"d8", x"d7", x"d2", x"d3", 
        x"d4", x"d4", x"d7", x"db", x"db", x"d7", x"d3", x"d5", x"d4", x"d1", x"d5", x"d6", x"d2", x"87", x"2a", 
        x"1f", x"24", x"4d", x"6a", x"63", x"66", x"4e", x"40", x"3c", x"34", x"35", x"43", x"57", x"6b", x"84", 
        x"9d", x"9d", x"9e", x"9f", x"9f", x"9e", x"9e", x"9c", x"9b", x"9a", x"9b", x"9c", x"9b", x"9a", x"9b", 
        x"9c", x"9e", x"9d", x"9c", x"9c", x"9d", x"9d", x"9c", x"9c", x"9c", x"9b", x"9b", x"9b", x"9d", x"9c", 
        x"9c", x"9d", x"9e", x"9e", x"9d", x"9c", x"9c", x"9d", x"9e", x"9c", x"9d", x"a0", x"9d", x"9d", x"9d", 
        x"9d", x"9d", x"9d", x"9d", x"9e", x"9c", x"9c", x"9c", x"9d", x"9d", x"9e", x"9f", x"9e", x"9e", x"9f", 
        x"9f", x"9f", x"9e", x"9d", x"9d", x"9e", x"9e", x"9f", x"9f", x"9e", x"9d", x"9d", x"9e", x"9e", x"9e", 
        x"9e", x"9e", x"9e", x"9e", x"9f", x"a0", x"9f", x"9e", x"9e", x"9f", x"a0", x"9e", x"9e", x"9e", x"9f", 
        x"9f", x"9f", x"9f", x"9e", x"9d", x"9e", x"a0", x"9f", x"9e", x"9d", x"9e", x"a0", x"a1", x"a2", x"a1", 
        x"a1", x"a0", x"8a", x"75", x"a3", x"a4", x"a6", x"a8", x"ab", x"ab", x"a7", x"ab", x"a9", x"a9", x"ab", 
        x"a8", x"a6", x"a9", x"a7", x"a5", x"ae", x"79", x"3f", x"66", x"79", x"7d", x"8d", x"9a", x"78", x"55", 
        x"38", x"2e", x"25", x"1e", x"12", x"09", x"03", x"02", x"03", x"04", x"05", x"18", x"46", x"63", x"7e", 
        x"80", x"56", x"c1", x"e2", x"d7", x"dd", x"d9", x"d6", x"df", x"d3", x"d3", x"d1", x"d2", x"d2", x"d3", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d4", x"d3", x"d3", x"d4", x"d5", x"d4", 
        x"d3", x"d3", x"d0", x"d3", x"d0", x"ce", x"d5", x"d3", x"d1", x"d5", x"d3", x"d1", x"d2", x"d4", x"d4", 
        x"ce", x"d1", x"d4", x"d4", x"d3", x"d1", x"ce", x"d8", x"d9", x"d5", x"bc", x"a3", x"9c", x"a1", x"bb", 
        x"d1", x"da", x"ef", x"f1", x"f0", x"eb", x"e3", x"d7", x"c8", x"bd", x"b6", x"b3", x"b1", x"b1", x"b6", 
        x"bc", x"c6", x"d3", x"de", x"e4", x"eb", x"f0", x"f3", x"f3", x"f0", x"ee", x"ec", x"ea", x"ec", x"ee", 
        x"ef", x"ed", x"ee", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"ef", x"ed", x"e8", x"f2", 
        x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"ef", x"ec", x"f1", x"f5", 
        x"f6", x"f5", x"f0", x"e5", x"dc", x"d3", x"c8", x"bf", x"be", x"c1", x"ca", x"d5", x"e1", x"ec", x"f3", 
        x"f4", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f0", x"f4", x"f6", x"f5", x"f2", 
        x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f5", x"f5", x"f4", x"f5", x"ef", x"ee", x"f4", x"f6", x"f8", x"f9", x"f7", x"f6", x"f5", x"f7", 
        x"f7", x"f5", x"f3", x"f2", x"f1", x"f1", x"f4", x"f4", x"f4", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f5", x"d3", 
        x"56", x"6d", x"66", x"a3", x"a2", x"95", x"85", x"74", x"6c", x"6d", x"77", x"80", x"89", x"96", x"9d", 
        x"9a", x"95", x"96", x"97", x"96", x"94", x"94", x"94", x"9a", x"a3", x"9d", x"96", x"96", x"9a", x"99", 
        x"93", x"93", x"96", x"9b", x"6e", x"4a", x"4a", x"82", x"8e", x"95", x"93", x"93", x"93", x"93", x"93", 
        x"94", x"94", x"93", x"91", x"90", x"91", x"93", x"93", x"93", x"91", x"92", x"93", x"93", x"91", x"90", 
        x"91", x"93", x"8f", x"89", x"a0", x"89", x"5a", x"b0", x"e4", x"e1", x"e2", x"de", x"db", x"dc", x"dc", 
        x"d8", x"da", x"df", x"dc", x"da", x"d7", x"d7", x"d7", x"d9", x"d8", x"d9", x"d8", x"d3", x"d6", x"d6", 
        x"da", x"db", x"d8", x"d6", x"d4", x"d4", x"d5", x"d7", x"da", x"db", x"d9", x"d8", x"d8", x"da", x"dd", 
        x"df", x"dd", x"db", x"d7", x"d6", x"d5", x"d5", x"d8", x"db", x"d7", x"d2", x"d4", x"d5", x"d6", x"dc", 
        x"df", x"da", x"d7", x"d7", x"d5", x"d0", x"cf", x"d8", x"da", x"d5", x"d3", x"d0", x"cd", x"88", x"2b", 
        x"25", x"22", x"32", x"35", x"2c", x"31", x"43", x"56", x"71", x"86", x"9c", x"af", x"bf", x"cd", x"d9", 
        x"9e", x"9e", x"9f", x"a0", x"a0", x"9f", x"9e", x"9c", x"9b", x"9b", x"9c", x"9d", x"9c", x"9a", x"9d", 
        x"a0", x"a1", x"a0", x"9c", x"9b", x"9c", x"9d", x"9c", x"9d", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", 
        x"9d", x"9c", x"9c", x"9e", x"9e", x"9c", x"9c", x"9d", x"9e", x"9d", x"9d", x"9f", x"9d", x"9c", x"9c", 
        x"9c", x"9c", x"9d", x"9f", x"9f", x"9e", x"9c", x"9d", x"9d", x"9d", x"9d", x"9d", x"9e", x"9e", x"9f", 
        x"a0", x"9f", x"9f", x"9e", x"9e", x"9e", x"9f", x"9f", x"9f", x"9e", x"9d", x"9d", x"9e", x"9e", x"9d", 
        x"9d", x"9d", x"9e", x"9e", x"9f", x"a0", x"a0", x"9f", x"9e", x"9f", x"a0", x"9f", x"9e", x"9f", x"9f", 
        x"9f", x"a0", x"a2", x"9f", x"9e", x"9f", x"a0", x"9f", x"9e", x"9e", x"9e", x"9e", x"a0", x"a3", x"a2", 
        x"a2", x"a2", x"89", x"72", x"a2", x"a5", x"a8", x"a9", x"ab", x"aa", x"a7", x"aa", x"a7", x"a5", x"a8", 
        x"a9", x"a7", x"ab", x"a9", x"a6", x"b2", x"7a", x"42", x"70", x"73", x"61", x"50", x"4a", x"35", x"25", 
        x"1c", x"17", x"0e", x"05", x"03", x"04", x"05", x"0a", x"0b", x"1b", x"30", x"54", x"8f", x"89", x"84", 
        x"77", x"51", x"bc", x"de", x"d4", x"d9", x"d8", x"d8", x"df", x"d3", x"d3", x"d1", x"d1", x"d2", x"d3", 
        x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d4", x"d3", x"d3", x"d4", x"d5", x"d4", 
        x"d3", x"d3", x"d1", x"d3", x"d0", x"ce", x"d5", x"d6", x"d2", x"d4", x"d2", x"cf", x"d0", x"d1", x"d4", 
        x"d2", x"d4", x"d2", x"cf", x"d6", x"d9", x"d3", x"bc", x"99", x"8c", x"9b", x"b7", x"cb", x"d9", x"de", 
        x"da", x"d4", x"e9", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"ef", x"eb", x"e6", x"dd", x"d4", x"ce", 
        x"c5", x"bd", x"b7", x"b2", x"af", x"b3", x"bb", x"c5", x"d0", x"dc", x"e7", x"ed", x"ee", x"ef", x"f0", 
        x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f0", x"ee", x"e8", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"eb", x"ef", x"f1", 
        x"f4", x"f4", x"f1", x"f3", x"f5", x"f4", x"f1", x"e9", x"de", x"d7", x"cd", x"c2", x"b9", x"b7", x"be", 
        x"ca", x"d4", x"e1", x"ee", x"f3", x"f5", x"f3", x"f1", x"f2", x"f5", x"f5", x"f5", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f5", x"f4", x"f2", x"f0", x"f0", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f5", x"f5", x"f3", x"f4", x"f0", x"ef", x"f6", x"f8", x"f9", x"f8", x"f6", x"f6", x"f6", x"f6", 
        x"f5", x"f4", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"f6", x"d9", 
        x"5d", x"6a", x"62", x"a5", x"a6", x"a3", x"a3", x"9e", x"95", x"87", x"7c", x"73", x"66", x"67", x"71", 
        x"7d", x"8a", x"95", x"99", x"90", x"8f", x"92", x"92", x"93", x"9a", x"99", x"95", x"94", x"98", x"98", 
        x"92", x"91", x"93", x"99", x"71", x"4c", x"46", x"80", x"8b", x"92", x"91", x"90", x"8f", x"8f", x"91", 
        x"92", x"92", x"90", x"91", x"90", x"90", x"91", x"92", x"92", x"91", x"91", x"91", x"91", x"91", x"90", 
        x"90", x"90", x"8d", x"87", x"a3", x"95", x"5f", x"aa", x"e1", x"d7", x"da", x"dd", x"e0", x"e0", x"de", 
        x"d8", x"d5", x"d7", x"da", x"db", x"da", x"d8", x"d6", x"d5", x"d4", x"da", x"de", x"da", x"d8", x"d5", 
        x"d5", x"d2", x"d5", x"d9", x"da", x"d8", x"d5", x"d4", x"da", x"df", x"e2", x"e2", x"df", x"db", x"d8", 
        x"d5", x"d4", x"d8", x"d7", x"d7", x"d5", x"d3", x"d4", x"d9", x"dc", x"db", x"dc", x"da", x"d9", x"d8", 
        x"d5", x"d6", x"d8", x"db", x"da", x"d6", x"d0", x"d1", x"d8", x"d6", x"d7", x"dc", x"da", x"98", x"37", 
        x"41", x"53", x"6b", x"7d", x"8f", x"9f", x"ad", x"bc", x"ca", x"d0", x"d3", x"d4", x"d5", x"d4", x"d7", 
        x"a0", x"9f", x"9f", x"9e", x"9e", x"9e", x"9e", x"9d", x"9c", x"9b", x"9c", x"9d", x"9d", x"9c", x"9c", 
        x"9d", x"9d", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9c", x"9b", 
        x"9d", x"9b", x"9b", x"9c", x"9d", x"9c", x"9c", x"9d", x"9d", x"9d", x"9d", x"9d", x"9e", x"9d", x"9d", 
        x"9c", x"9c", x"9d", x"9e", x"9f", x"9f", x"9f", x"9e", x"9e", x"9d", x"9d", x"9e", x"9f", x"9f", x"9f", 
        x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9e", x"9d", x"9d", x"a0", x"a0", x"9e", 
        x"9e", x"9f", x"a0", x"a0", x"9f", x"a0", x"a1", x"a0", x"9f", x"a0", x"a0", x"9f", x"9f", x"9f", x"9f", 
        x"9e", x"9f", x"a1", x"a0", x"9e", x"9f", x"a0", x"9f", x"9f", x"9e", x"a0", x"9e", x"a0", x"a2", x"a0", 
        x"a2", x"a4", x"8b", x"73", x"a4", x"a6", x"a9", x"a9", x"a9", x"aa", x"a9", x"a9", x"a8", x"a8", x"ab", 
        x"ab", x"a7", x"a9", x"a7", x"a8", x"b3", x"81", x"42", x"4e", x"4b", x"3d", x"2e", x"28", x"1c", x"10", 
        x"08", x"05", x"04", x"04", x"06", x"0f", x"27", x"45", x"3e", x"3b", x"4b", x"60", x"96", x"83", x"7f", 
        x"79", x"52", x"be", x"e2", x"d5", x"d7", x"d7", x"d8", x"de", x"d2", x"d2", x"d2", x"d1", x"d2", x"d4", 
        x"d4", x"d5", x"d5", x"d5", x"d5", x"d5", x"d5", x"d5", x"d5", x"d4", x"d4", x"d4", x"d4", x"d5", x"d4", 
        x"d5", x"d3", x"d3", x"d5", x"d2", x"d0", x"d5", x"d5", x"d1", x"d3", x"d1", x"d0", x"d3", x"d3", x"d2", 
        x"d4", x"d4", x"d8", x"dd", x"c9", x"ab", x"8b", x"84", x"8a", x"a6", x"c8", x"d8", x"de", x"da", x"d7", 
        x"d7", x"d6", x"e8", x"ee", x"ef", x"ef", x"ef", x"ed", x"ed", x"ef", x"f0", x"f0", x"ef", x"f1", x"f1", 
        x"ec", x"e7", x"e1", x"d9", x"d2", x"cd", x"c3", x"b9", x"b2", x"ae", x"ad", x"ad", x"bd", x"cb", x"d8", 
        x"e3", x"e8", x"ec", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"ee", x"e8", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"ed", x"f2", x"f1", 
        x"f3", x"f3", x"f1", x"f3", x"f3", x"f2", x"f2", x"f3", x"f5", x"f5", x"f0", x"e6", x"dc", x"d5", x"ce", 
        x"c4", x"b8", x"b3", x"bb", x"c7", x"d8", x"e6", x"ee", x"f2", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f4", x"f4", x"f3", x"f2", x"f3", x"f1", x"f0", x"f7", x"f9", x"f9", x"f8", x"f7", x"f6", x"f6", x"f5", 
        x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"f0", x"f2", x"f1", x"f0", x"f3", x"f6", x"f6", x"db", 
        x"63", x"6b", x"62", x"a7", x"ad", x"9f", x"9f", x"9f", x"9e", x"9b", x"98", x"92", x"87", x"7c", x"70", 
        x"67", x"63", x"6e", x"7b", x"85", x"8e", x"93", x"93", x"92", x"99", x"9d", x"94", x"8e", x"91", x"95", 
        x"92", x"90", x"8e", x"94", x"71", x"4e", x"41", x"7d", x"89", x"91", x"90", x"90", x"8e", x"8e", x"8f", 
        x"8f", x"8f", x"8e", x"90", x"8f", x"8e", x"8e", x"8f", x"91", x"91", x"8f", x"8f", x"8f", x"8f", x"8f", 
        x"8e", x"8e", x"8b", x"85", x"9d", x"96", x"5a", x"a0", x"e6", x"de", x"de", x"de", x"dd", x"dc", x"da", 
        x"d8", x"d7", x"d6", x"d5", x"d6", x"d9", x"db", x"db", x"dc", x"dd", x"db", x"d9", x"d8", x"d9", x"d9", 
        x"db", x"dc", x"d8", x"d4", x"d4", x"d7", x"db", x"de", x"df", x"de", x"db", x"d8", x"d6", x"d6", x"d8", 
        x"d9", x"d8", x"da", x"da", x"db", x"dd", x"df", x"df", x"e1", x"de", x"d7", x"d4", x"d4", x"d7", x"da", 
        x"d9", x"d7", x"d7", x"d7", x"d8", x"d8", x"d9", x"de", x"e2", x"e1", x"e3", x"e7", x"e1", x"b5", x"8d", 
        x"99", x"aa", x"b7", x"c3", x"ce", x"d2", x"d3", x"d7", x"d9", x"d7", x"d7", x"d8", x"d8", x"d8", x"d9", 
        x"a1", x"a0", x"9e", x"9c", x"9c", x"9c", x"9d", x"9f", x"9e", x"9d", x"9d", x"9e", x"9e", x"9e", x"9d", 
        x"9c", x"9b", x"9b", x"9d", x"9e", x"9d", x"9c", x"9d", x"9d", x"9d", x"9d", x"9e", x"9d", x"9c", x"9e", 
        x"9f", x"9e", x"9d", x"9e", x"9f", x"9e", x"9c", x"9c", x"9b", x"9d", x"9d", x"9b", x"9e", x"a0", x"a0", 
        x"9e", x"9d", x"9c", x"9c", x"9c", x"9e", x"a0", x"9f", x"9e", x"9f", x"9f", x"a0", x"a0", x"a0", x"9f", 
        x"9e", x"9f", x"a0", x"a0", x"a0", x"9e", x"9f", x"9f", x"9f", x"9f", x"9e", x"9f", x"a0", x"a1", x"a0", 
        x"9f", x"a0", x"a0", x"a0", x"9f", x"a0", x"a1", x"a1", x"a0", x"a0", x"a0", x"9f", x"a0", x"a0", x"9f", 
        x"9d", x"9d", x"9f", x"a0", x"9f", x"a0", x"a0", x"a0", x"9f", x"9f", x"a2", x"a2", x"a1", x"a1", x"9f", 
        x"a1", x"a3", x"8d", x"76", x"a3", x"a4", x"a6", x"a6", x"a8", x"a8", x"a7", x"a9", x"ac", x"a8", x"a4", 
        x"a7", x"a9", x"ae", x"b6", x"a9", x"84", x"59", x"38", x"39", x"33", x"28", x"14", x"0c", x"07", x"06", 
        x"04", x"04", x"08", x"12", x"34", x"62", x"87", x"8f", x"61", x"45", x"4d", x"5b", x"96", x"85", x"7f", 
        x"77", x"53", x"bc", x"e3", x"d8", x"da", x"da", x"d9", x"dd", x"d1", x"d1", x"d0", x"d1", x"d2", x"d3", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d4", x"d4", x"d5", x"d5", x"d5", 
        x"d5", x"d2", x"d3", x"d4", x"d2", x"d0", x"d2", x"d1", x"d0", x"d1", x"cf", x"cf", x"d2", x"d1", x"d6", 
        x"d9", x"d0", x"b7", x"8e", x"72", x"7e", x"9e", x"be", x"cf", x"d7", x"da", x"d9", x"d7", x"d6", x"d7", 
        x"db", x"d6", x"e6", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"ef", x"f0", x"f0", x"ee", x"ed", x"ee", 
        x"ee", x"ef", x"f2", x"f1", x"f0", x"f0", x"ea", x"e7", x"e5", x"dd", x"d2", x"c5", x"bb", x"b5", x"ab", 
        x"a3", x"a4", x"ae", x"ba", x"d1", x"de", x"e7", x"ef", x"f2", x"f2", x"f0", x"ed", x"ed", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"ee", x"ec", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"ed", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ee", x"e8", x"f2", 
        x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"eb", x"f3", x"f0", 
        x"f1", x"f1", x"f1", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f5", x"f4", 
        x"ee", x"e7", x"de", x"d5", x"cb", x"bc", x"b1", x"b4", x"c1", x"d3", x"e1", x"ea", x"f2", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f1", x"f0", x"f2", x"f4", x"f3", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f5", 
        x"f4", x"f3", x"f3", x"f0", x"f2", x"f0", x"f1", x"f8", x"f9", x"f9", x"f8", x"f6", x"f6", x"f5", x"f4", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f2", x"f5", x"f7", x"f6", x"e2", 
        x"6c", x"6c", x"66", x"b0", x"c4", x"a0", x"9f", x"a1", x"9b", x"9a", x"98", x"96", x"9a", x"93", x"90", 
        x"8f", x"87", x"77", x"69", x"59", x"61", x"6f", x"81", x"92", x"9d", x"9f", x"97", x"8e", x"8d", x"90", 
        x"92", x"92", x"8f", x"93", x"71", x"4f", x"3e", x"79", x"87", x"91", x"8f", x"8f", x"8e", x"8d", x"8e", 
        x"8d", x"8c", x"8c", x"8e", x"8e", x"8d", x"8c", x"8d", x"8f", x"90", x"8d", x"8d", x"8c", x"8d", x"8d", 
        x"8c", x"8a", x"89", x"86", x"9f", x"a2", x"5e", x"93", x"e2", x"d9", x"d9", x"de", x"e2", x"e0", x"dc", 
        x"db", x"da", x"d9", x"dd", x"df", x"de", x"db", x"d9", x"d9", x"dd", x"df", x"e0", x"de", x"db", x"d9", 
        x"d9", x"da", x"dd", x"df", x"dd", x"d9", x"d7", x"d7", x"d6", x"d8", x"dc", x"dd", x"de", x"dd", x"de", 
        x"de", x"df", x"e3", x"e3", x"e1", x"dc", x"d7", x"d4", x"d9", x"dc", x"da", x"da", x"d8", x"d7", x"d7", 
        x"d7", x"da", x"dd", x"e1", x"e4", x"e7", x"e9", x"e8", x"e4", x"de", x"d3", x"c9", x"c8", x"c0", x"c6", 
        x"cd", x"d6", x"d5", x"d7", x"d8", x"d7", x"d9", x"db", x"d9", x"d8", x"d8", x"d9", x"d9", x"d6", x"d5", 
        x"a0", x"a0", x"9f", x"9e", x"9d", x"9d", x"9d", x"9e", x"9d", x"9d", x"9d", x"9e", x"9e", x"9d", x"9e", 
        x"9e", x"9d", x"9e", x"9f", x"a0", x"9f", x"9e", x"9d", x"9c", x"9c", x"9e", x"9e", x"9d", x"9d", x"9d", 
        x"9d", x"9d", x"9c", x"9c", x"9d", x"9f", x"9b", x"9b", x"9a", x"9d", x"9d", x"99", x"9d", x"a0", x"a0", 
        x"9f", x"9d", x"9c", x"9c", x"9c", x"9e", x"a0", x"a0", x"a0", x"9f", x"9e", x"9e", x"9e", x"9e", x"9f", 
        x"9f", x"9f", x"a0", x"a0", x"9f", x"9d", x"9e", x"9f", x"a0", x"9f", x"9f", x"9f", x"9f", x"a0", x"a0", 
        x"a0", x"a0", x"9f", x"9f", x"9f", x"a1", x"a2", x"a2", x"a1", x"a0", x"a0", x"9f", x"a1", x"a2", x"a2", 
        x"9f", x"9f", x"a0", x"a0", x"a0", x"a0", x"a0", x"a0", x"a0", x"a0", x"a2", x"a4", x"a2", x"9f", x"a0", 
        x"a1", x"a2", x"8d", x"75", x"9f", x"9f", x"a3", x"a5", x"a5", x"a4", x"a5", x"a7", x"a9", x"a8", x"ad", 
        x"b1", x"ab", x"98", x"74", x"54", x"3a", x"37", x"2e", x"19", x"0c", x"07", x"04", x"05", x"04", x"09", 
        x"15", x"2b", x"5c", x"82", x"92", x"9b", x"9b", x"91", x"5b", x"42", x"50", x"5a", x"92", x"84", x"83", 
        x"7e", x"54", x"bb", x"e1", x"d6", x"d8", x"d8", x"d6", x"dd", x"d1", x"d1", x"d0", x"d0", x"d2", x"d2", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d5", x"d5", x"d5", x"d4", x"d5", 
        x"d3", x"d1", x"d2", x"d2", x"d0", x"cf", x"d0", x"d2", x"d3", x"d5", x"d5", x"d9", x"d8", x"ce", x"b9", 
        x"95", x"79", x"83", x"9f", x"bd", x"ce", x"d0", x"d4", x"d6", x"d5", x"d7", x"d6", x"d7", x"d8", x"d7", 
        x"dc", x"d6", x"e5", x"ef", x"ef", x"ed", x"ed", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ed", x"ef", 
        x"ee", x"ed", x"ee", x"ef", x"ef", x"f0", x"ee", x"ed", x"ef", x"f0", x"ee", x"eb", x"ec", x"eb", x"e8", 
        x"e1", x"d4", x"c6", x"ba", x"b0", x"aa", x"a7", x"aa", x"b3", x"c1", x"cf", x"db", x"e3", x"e7", x"eb", 
        x"ee", x"f1", x"f3", x"f2", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", x"ee", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ee", x"ee", x"ef", x"f0", x"ef", x"ed", x"e7", x"f1", 
        x"f1", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f3", x"f3", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f2", x"ef", x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"ed", x"f6", x"f3", 
        x"f5", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f1", x"ed", x"e9", x"e4", x"da", x"ce", x"c1", x"b5", x"b4", x"bc", x"cd", x"de", 
        x"e9", x"eb", x"ee", x"f0", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f5", 
        x"f4", x"f5", x"f5", x"f2", x"f3", x"f0", x"f1", x"f8", x"f8", x"f8", x"f8", x"f6", x"f5", x"f4", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ee", x"f0", x"f4", x"f5", x"f6", x"f7", x"e9", 
        x"6f", x"64", x"62", x"a7", x"d5", x"a9", x"9e", x"a2", x"9c", x"9c", x"99", x"97", x"93", x"92", x"92", 
        x"91", x"8e", x"8c", x"8d", x"8b", x"84", x"70", x"60", x"60", x"74", x"88", x"95", x"92", x"8f", x"90", 
        x"8f", x"8d", x"8b", x"8f", x"6f", x"51", x"3e", x"77", x"86", x"90", x"8a", x"8b", x"8c", x"8b", x"8b", 
        x"8a", x"8b", x"8b", x"8a", x"8b", x"8c", x"8b", x"8b", x"8c", x"8c", x"8c", x"8a", x"8a", x"8b", x"8b", 
        x"8a", x"88", x"8b", x"83", x"8c", x"92", x"52", x"81", x"e2", x"df", x"dc", x"de", x"df", x"de", x"dd", 
        x"e2", x"e3", x"e0", x"dc", x"da", x"db", x"dd", x"de", x"de", x"de", x"de", x"de", x"de", x"dd", x"dd", 
        x"dc", x"db", x"d9", x"d6", x"d8", x"db", x"dc", x"dc", x"dd", x"df", x"e2", x"e2", x"e3", x"e3", x"e4", 
        x"de", x"da", x"dc", x"da", x"da", x"db", x"db", x"db", x"e0", x"df", x"dc", x"dc", x"dd", x"de", x"e2", 
        x"e6", x"e9", x"e9", x"e5", x"de", x"d9", x"d6", x"ce", x"c9", x"c8", x"c9", x"cc", x"d4", x"d9", x"db", 
        x"d5", x"d7", x"d8", x"da", x"db", x"da", x"d8", x"d8", x"d6", x"da", x"da", x"d8", x"d7", x"d8", x"d6", 
        x"9f", x"a0", x"a0", x"9f", x"9e", x"9d", x"9d", x"9d", x"9c", x"9c", x"9d", x"9e", x"9e", x"9c", x"9b", 
        x"9b", x"9d", x"9d", x"9e", x"9e", x"9f", x"9f", x"9d", x"9c", x"9d", x"9e", x"9e", x"9d", x"9d", x"9e", 
        x"9e", x"9e", x"9e", x"9c", x"9e", x"a0", x"9b", x"9b", x"9a", x"9c", x"9c", x"99", x"9c", x"9e", x"9e", 
        x"9e", x"9d", x"9e", x"9e", x"9f", x"9e", x"9f", x"a1", x"a0", x"9f", x"9d", x"9a", x"9c", x"9e", x"9f", 
        x"a0", x"a0", x"a0", x"a0", x"9f", x"9d", x"9e", x"9f", x"a0", x"a0", x"a0", x"a0", x"9f", x"9f", x"9f", 
        x"a0", x"a0", x"9f", x"9f", x"9f", x"a1", x"a2", x"a1", x"a0", x"a0", x"a0", x"9f", x"a1", x"a3", x"a2", 
        x"a1", x"a0", x"a1", x"a1", x"a0", x"a0", x"a0", x"a0", x"a0", x"a0", x"a0", x"a2", x"a1", x"a0", x"a1", 
        x"a1", x"a2", x"8e", x"77", x"a3", x"a5", x"a9", x"ab", x"ab", x"a6", x"a6", x"a6", x"a9", x"ab", x"a5", 
        x"8e", x"6c", x"47", x"38", x"3b", x"2a", x"17", x"0b", x"0c", x"07", x"04", x"04", x"0b", x"1f", x"43", 
        x"77", x"94", x"a8", x"9d", x"92", x"96", x"94", x"8d", x"5c", x"41", x"4e", x"57", x"91", x"87", x"85", 
        x"7c", x"54", x"b9", x"e2", x"d6", x"d7", x"d8", x"d9", x"df", x"d2", x"d2", x"d1", x"d0", x"d1", x"d1", 
        x"d1", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d3", x"d4", 
        x"d2", x"cf", x"d1", x"d0", x"cf", x"ce", x"cf", x"d2", x"d1", x"d3", x"d0", x"c3", x"a5", x"85", x"7c", 
        x"90", x"ba", x"d2", x"d5", x"d2", x"d1", x"d1", x"d3", x"d2", x"d0", x"d6", x"d7", x"d6", x"d9", x"d8", 
        x"db", x"d7", x"e7", x"f0", x"ee", x"ed", x"ef", x"ef", x"ee", x"ee", x"ef", x"f1", x"f0", x"ee", x"f0", 
        x"ee", x"ed", x"ee", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f1", 
        x"ef", x"ee", x"ee", x"ee", x"ea", x"e6", x"de", x"d1", x"c3", x"b5", x"aa", x"a6", x"a8", x"af", x"ba", 
        x"c8", x"d6", x"e0", x"e6", x"ea", x"ed", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"ee", x"ec", x"ee", x"f0", x"ef", x"ed", x"e8", x"f1", 
        x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"f1", x"f0", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"ec", x"f3", x"f1", 
        x"f3", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f4", x"f4", x"f3", x"f2", x"f3", x"f4", 
        x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", x"ef", x"e9", x"de", x"cd", x"c2", x"bc", 
        x"bb", x"bf", x"cd", x"da", x"e5", x"eb", x"ec", x"ef", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f5", x"f5", x"f4", x"f4", x"ef", x"ef", x"f8", x"f7", x"f7", x"f7", x"f7", x"f5", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"ee", x"ed", x"f1", x"f4", x"f4", x"f4", x"f7", x"ed", 
        x"76", x"65", x"65", x"a1", x"e0", x"ba", x"a1", x"a3", x"9f", x"9f", x"9a", x"97", x"96", x"95", x"93", 
        x"91", x"8e", x"8f", x"8f", x"89", x"8d", x"8f", x"90", x"8c", x"7f", x"6e", x"66", x"6a", x"75", x"85", 
        x"8f", x"90", x"8a", x"8f", x"70", x"54", x"40", x"76", x"86", x"8e", x"87", x"88", x"89", x"8a", x"89", 
        x"89", x"8a", x"89", x"88", x"8a", x"8a", x"8b", x"88", x"89", x"89", x"8a", x"8a", x"8a", x"8a", x"8b", 
        x"89", x"87", x"88", x"83", x"8d", x"a0", x"5c", x"7e", x"de", x"dd", x"dd", x"e1", x"e3", x"e0", x"dc", 
        x"dd", x"df", x"e1", x"e3", x"e1", x"dc", x"d9", x"d9", x"db", x"df", x"e3", x"e3", x"de", x"d7", x"d8", 
        x"da", x"db", x"dd", x"df", x"e0", x"de", x"dc", x"db", x"e0", x"e2", x"e4", x"e2", x"de", x"da", x"d9", 
        x"dd", x"dd", x"df", x"de", x"de", x"dc", x"da", x"dd", x"e4", x"e7", x"e7", x"e8", x"e8", x"e7", x"e4", 
        x"df", x"da", x"d3", x"cc", x"ca", x"cc", x"d0", x"d6", x"d8", x"da", x"d9", x"db", x"dc", x"db", x"da", 
        x"d7", x"da", x"db", x"d8", x"d8", x"da", x"db", x"d9", x"d6", x"da", x"da", x"da", x"da", x"d9", x"d6", 
        x"a1", x"a0", x"a0", x"9f", x"9e", x"9e", x"9e", x"9e", x"9d", x"9d", x"9d", x"9d", x"9d", x"9e", x"9f", 
        x"9d", x"9f", x"9f", x"9c", x"9d", x"9d", x"9c", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9d", 
        x"9d", x"9d", x"9d", x"9d", x"9d", x"9d", x"9b", x"9d", x"9e", x"9d", x"9c", x"9c", x"9c", x"9e", x"a0", 
        x"a1", x"9e", x"9d", x"9f", x"9e", x"9b", x"9d", x"a1", x"9f", x"9e", x"9e", x"9d", x"9f", x"9e", x"9f", 
        x"9e", x"9e", x"a1", x"a0", x"a1", x"9e", x"a0", x"a2", x"a1", x"a0", x"a0", x"9f", x"a0", x"9f", x"9f", 
        x"a0", x"a2", x"a1", x"a0", x"9f", x"a0", x"a1", x"a1", x"9f", x"9f", x"a0", x"a1", x"a1", x"a0", x"a0", 
        x"a1", x"a1", x"a0", x"a0", x"a1", x"a1", x"a1", x"a2", x"a2", x"a2", x"9f", x"9f", x"a2", x"a1", x"9f", 
        x"9e", x"a0", x"8b", x"73", x"a1", x"a3", x"a6", x"a6", x"ab", x"ab", x"af", x"ad", x"9d", x"81", x"5b", 
        x"40", x"36", x"30", x"24", x"13", x"08", x"07", x"0c", x"2c", x"1c", x"08", x"0b", x"3c", x"86", x"a9", 
        x"b1", x"ad", x"a6", x"99", x"90", x"93", x"93", x"8f", x"5e", x"42", x"4f", x"5a", x"90", x"82", x"84", 
        x"7c", x"56", x"b9", x"e3", x"d7", x"d8", x"d7", x"da", x"e0", x"d1", x"d3", x"d1", x"d2", x"d2", x"d1", 
        x"d2", x"d4", x"d3", x"d2", x"d3", x"d4", x"d2", x"d0", x"d1", x"d3", x"d3", x"d4", x"d3", x"d2", x"d3", 
        x"d1", x"d1", x"d4", x"d0", x"d0", x"d4", x"d4", x"d0", x"c2", x"ab", x"8f", x"7d", x"8e", x"af", x"cb", 
        x"d3", x"d6", x"d5", x"d4", x"d3", x"d1", x"d0", x"d1", x"d0", x"d3", x"db", x"da", x"d7", x"d8", x"da", 
        x"dc", x"d7", x"e6", x"f2", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ee", x"ed", x"ed", x"ee", x"ee", x"ec", x"e8", x"e1", x"d8", x"cc", x"be", 
        x"b5", x"ae", x"ac", x"af", x"b8", x"c5", x"d1", x"da", x"e0", x"e5", x"e9", x"ed", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"ee", x"ec", x"ef", x"ef", x"ed", x"ee", x"ef", x"ee", x"ef", x"ed", x"ec", x"ed", x"ef", 
        x"f0", x"f2", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ee", x"ef", x"f2", x"f0", x"ec", x"e9", x"f0", 
        x"f0", x"f1", x"f1", x"f2", x"f3", x"f1", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"ec", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"eb", 
        x"e1", x"d7", x"ca", x"be", x"ba", x"c2", x"ce", x"d9", x"e2", x"e9", x"ee", x"f2", x"f3", x"f2", x"f1", 
        x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f0", x"f0", x"f0", x"f1", 
        x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f5", x"f5", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f4", 
        x"f3", x"f3", x"f2", x"f5", x"f6", x"f0", x"ec", x"f5", x"f7", x"f7", x"f6", x"f5", x"f5", x"f3", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"ef", 
        x"ee", x"f0", x"f1", x"ef", x"ef", x"ef", x"f0", x"ef", x"f1", x"f5", x"f4", x"f4", x"f4", x"f6", x"ef", 
        x"81", x"66", x"67", x"9b", x"e5", x"cd", x"a9", x"9f", x"a0", x"9c", x"9c", x"96", x"96", x"95", x"97", 
        x"96", x"92", x"90", x"90", x"8d", x"8b", x"8c", x"8d", x"90", x"98", x"97", x"94", x"87", x"6a", x"5e", 
        x"6c", x"7b", x"80", x"8d", x"70", x"58", x"46", x"74", x"86", x"8a", x"86", x"87", x"89", x"88", x"89", 
        x"8a", x"88", x"86", x"88", x"87", x"85", x"87", x"85", x"88", x"86", x"88", x"87", x"89", x"88", x"89", 
        x"87", x"87", x"86", x"81", x"91", x"ae", x"5b", x"77", x"e0", x"dc", x"d8", x"db", x"de", x"e0", x"e0", 
        x"e0", x"df", x"df", x"e0", x"df", x"df", x"e2", x"e2", x"dc", x"d6", x"d9", x"dc", x"e0", x"e0", x"e2", 
        x"e0", x"dd", x"dd", x"de", x"e1", x"e3", x"e2", x"df", x"db", x"db", x"df", x"de", x"df", x"de", x"df", 
        x"e0", x"d8", x"d8", x"de", x"e2", x"e6", x"e8", x"e7", x"e7", x"e5", x"e2", x"dd", x"d9", x"d4", x"cf", 
        x"cc", x"cf", x"d3", x"d6", x"d8", x"d8", x"d8", x"d8", x"d9", x"da", x"da", x"db", x"dc", x"dc", x"da", 
        x"da", x"da", x"db", x"db", x"da", x"d9", x"da", x"da", x"d9", x"d9", x"d8", x"d9", x"d9", x"d9", x"d9", 
        x"9f", x"9f", x"a0", x"a0", x"9f", x"9f", x"9f", x"9f", x"9e", x"9e", x"9d", x"9d", x"9d", x"9e", x"9e", 
        x"9d", x"9e", x"9f", x"9d", x"9e", x"9e", x"9d", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9d", 
        x"9d", x"9d", x"9d", x"9d", x"9d", x"9d", x"9d", x"9e", x"9f", x"9e", x"9d", x"9e", x"9f", x"9e", x"a0", 
        x"9f", x"9e", x"9e", x"a0", x"9e", x"9c", x"9e", x"a1", x"9f", x"9e", x"9f", x"9d", x"9e", x"9e", x"a0", 
        x"a0", x"a0", x"a2", x"a0", x"a0", x"9f", x"a0", x"a1", x"a1", x"a0", x"a0", x"a0", x"a0", x"9f", x"9f", 
        x"a0", x"a1", x"a0", x"9f", x"a0", x"a1", x"a0", x"a0", x"a0", x"a0", x"a0", x"a1", x"a1", x"a0", x"a0", 
        x"a1", x"a1", x"a0", x"a0", x"a1", x"a1", x"a2", x"a2", x"a1", x"a1", x"9f", x"9e", x"a1", x"a1", x"a0", 
        x"a0", x"a3", x"90", x"77", x"9e", x"a3", x"aa", x"ab", x"ac", x"a9", x"94", x"73", x"4e", x"34", x"33", 
        x"2f", x"18", x"07", x"08", x"06", x"10", x"26", x"42", x"5b", x"35", x"0e", x"1a", x"79", x"b6", x"af", 
        x"a7", x"a7", x"a9", x"9f", x"8c", x"90", x"97", x"8e", x"5c", x"41", x"4b", x"56", x"94", x"8d", x"88", 
        x"7b", x"4e", x"ba", x"df", x"d6", x"d9", x"d8", x"d8", x"e0", x"d2", x"d4", x"d2", x"d3", x"d2", x"d1", 
        x"d5", x"d6", x"d5", x"d3", x"d2", x"d3", x"d3", x"cf", x"d0", x"d4", x"d4", x"d3", x"d5", x"d4", x"d0", 
        x"ce", x"d2", x"d7", x"d7", x"d3", x"c4", x"ac", x"91", x"79", x"7d", x"a7", x"d0", x"e0", x"dd", x"d4", 
        x"d4", x"d3", x"d2", x"d3", x"d4", x"d3", x"d2", x"d1", x"ce", x"d1", x"d8", x"d9", x"d9", x"d8", x"d9", 
        x"db", x"d5", x"e4", x"f1", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ec", x"ed", x"f0", x"f5", x"f7", 
        x"f5", x"ef", x"e8", x"dc", x"ca", x"bd", x"b1", x"ac", x"ae", x"b2", x"b9", x"c6", x"ce", x"d7", x"e0", 
        x"e6", x"ea", x"eb", x"f0", x"f0", x"ee", x"ed", x"ef", x"f0", x"ee", x"ef", x"ef", x"f0", x"f2", x"f1", 
        x"ee", x"ee", x"f1", x"f3", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"ee", x"e9", x"e5", x"f0", 
        x"f0", x"f1", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f3", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"ed", x"f3", x"f4", 
        x"f2", x"f2", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f4", x"f4", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"ef", x"f0", x"f2", x"f3", 
        x"f4", x"f5", x"f7", x"f3", x"ea", x"dc", x"c9", x"bd", x"bb", x"bf", x"c7", x"d2", x"dc", x"e5", x"ea", 
        x"ed", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f3", x"f4", x"f0", x"f0", x"f4", x"f6", x"f3", x"f0", x"f2", x"f5", x"f4", x"f2", x"f2", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f4", 
        x"f3", x"f3", x"f3", x"f5", x"f6", x"f0", x"ed", x"f7", x"f8", x"f8", x"f6", x"f4", x"f3", x"f3", x"f1", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"ef", 
        x"ef", x"f0", x"f1", x"ef", x"ef", x"ef", x"f1", x"f1", x"f3", x"f6", x"f5", x"f4", x"f3", x"f5", x"ef", 
        x"88", x"65", x"6a", x"96", x"e2", x"d8", x"bd", x"a1", x"9d", x"9f", x"9c", x"96", x"99", x"97", x"97", 
        x"96", x"93", x"93", x"94", x"93", x"8e", x"8e", x"8d", x"8e", x"95", x"99", x"9a", x"a3", x"9c", x"8c", 
        x"79", x"6a", x"5f", x"6c", x"61", x"59", x"4e", x"73", x"84", x"8a", x"89", x"88", x"87", x"84", x"85", 
        x"87", x"87", x"85", x"87", x"86", x"85", x"86", x"85", x"89", x"88", x"83", x"81", x"83", x"83", x"86", 
        x"86", x"85", x"84", x"81", x"89", x"a3", x"50", x"66", x"dd", x"e6", x"e4", x"e2", x"e1", x"e0", x"e0", 
        x"e1", x"e3", x"e5", x"e1", x"db", x"d9", x"dd", x"df", x"e1", x"e5", x"e3", x"e1", x"e0", x"df", x"e0", 
        x"e2", x"e5", x"e3", x"df", x"db", x"db", x"de", x"e1", x"e2", x"e1", x"e2", x"de", x"dd", x"dd", x"df", 
        x"e8", x"e7", x"e7", x"e9", x"e6", x"e1", x"dd", x"d9", x"d6", x"d1", x"ce", x"cd", x"d1", x"d5", x"d8", 
        x"db", x"dc", x"dc", x"dc", x"db", x"da", x"d9", x"d9", x"d9", x"d9", x"da", x"da", x"da", x"da", x"d8", 
        x"d9", x"da", x"db", x"db", x"db", x"da", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"d9", x"d9", 
        x"9e", x"9f", x"a0", x"a1", x"a1", x"a0", x"9f", x"9f", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", 
        x"9d", x"9d", x"9e", x"9d", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", 
        x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9d", x"9d", x"9d", x"9c", x"9b", x"9c", x"9e", x"a0", x"a1", 
        x"9f", x"9e", x"9f", x"a0", x"9d", x"9b", x"9d", x"a0", x"9e", x"9f", x"a1", x"9f", x"9f", x"9e", x"a0", 
        x"a0", x"a1", x"a1", x"a0", x"a0", x"a0", x"9f", x"9f", x"a0", x"a0", x"a0", x"9f", x"a1", x"a0", x"9f", 
        x"a0", x"a1", x"a0", x"9f", x"a0", x"a0", x"9f", x"a0", x"a1", x"a1", x"a0", x"a1", x"a1", x"a0", x"a1", 
        x"a1", x"a1", x"a0", x"a1", x"a2", x"a2", x"a2", x"a1", x"a1", x"a0", x"a1", x"a1", x"a2", x"a2", x"a1", 
        x"a1", x"a4", x"8e", x"72", x"a2", x"a9", x"aa", x"9b", x"7f", x"64", x"4c", x"39", x"31", x"26", x"15", 
        x"0a", x"06", x"09", x"1a", x"2c", x"53", x"7b", x"93", x"70", x"44", x"25", x"26", x"82", x"ac", x"a8", 
        x"a9", x"aa", x"aa", x"9f", x"8e", x"93", x"96", x"8c", x"5f", x"42", x"50", x"5f", x"94", x"7f", x"5e", 
        x"47", x"4a", x"ba", x"e1", x"d8", x"d9", x"d9", x"dc", x"e2", x"d3", x"d5", x"d1", x"d3", x"d2", x"d1", 
        x"d1", x"d1", x"d2", x"d3", x"d2", x"d1", x"d1", x"d3", x"d2", x"d1", x"d0", x"d0", x"d2", x"d3", x"d4", 
        x"d7", x"d5", x"c7", x"aa", x"92", x"87", x"87", x"9e", x"ba", x"d4", x"d9", x"d6", x"d5", x"d6", x"d1", 
        x"d3", x"d3", x"d2", x"d3", x"d4", x"d1", x"d1", x"d1", x"cf", x"d2", x"d8", x"d8", x"d7", x"d7", x"d9", 
        x"d9", x"d4", x"e2", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ec", x"f0", x"f1", x"f0", x"ee", 
        x"ee", x"ee", x"ef", x"f0", x"f0", x"ec", x"ea", x"e7", x"df", x"d4", x"cc", x"c7", x"c1", x"bd", x"bc", 
        x"be", x"c3", x"c9", x"ce", x"d7", x"e0", x"e5", x"eb", x"ef", x"f1", x"f3", x"f2", x"f1", x"f1", x"ef", 
        x"ee", x"ef", x"f1", x"f2", x"f0", x"f1", x"ef", x"f1", x"f0", x"f0", x"f0", x"ee", x"eb", x"e8", x"f2", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ed", x"f2", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f4", x"f1", x"f0", x"f0", x"ee", x"eb", x"e8", x"da", x"d2", x"cc", x"c7", x"c6", x"c8", 
        x"ca", x"d2", x"d8", x"e1", x"ec", x"f3", x"f4", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f4", 
        x"f3", x"f4", x"f4", x"f5", x"f4", x"f0", x"ee", x"f7", x"f8", x"f7", x"f5", x"f3", x"f3", x"f2", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", 
        x"f0", x"f1", x"f1", x"ee", x"ee", x"ee", x"f1", x"f2", x"f4", x"f7", x"f5", x"f5", x"f3", x"f4", x"ef", 
        x"8f", x"61", x"6c", x"8f", x"df", x"d9", x"d1", x"a8", x"9d", x"a0", x"a1", x"99", x"9b", x"98", x"97", 
        x"96", x"94", x"94", x"95", x"92", x"90", x"90", x"8f", x"8e", x"93", x"98", x"99", x"9b", x"94", x"8d", 
        x"8b", x"8b", x"8b", x"85", x"6d", x"5b", x"47", x"69", x"77", x"73", x"78", x"80", x"87", x"89", x"87", 
        x"87", x"85", x"83", x"83", x"84", x"82", x"82", x"80", x"83", x"84", x"84", x"82", x"82", x"82", x"84", 
        x"84", x"83", x"85", x"81", x"82", x"a3", x"61", x"6c", x"dd", x"e2", x"df", x"e3", x"e5", x"e3", x"e0", 
        x"dd", x"da", x"dc", x"e1", x"e3", x"e4", x"e3", x"e1", x"df", x"de", x"e1", x"e3", x"e3", x"e4", x"e0", 
        x"df", x"dc", x"dc", x"de", x"e0", x"e1", x"e0", x"de", x"de", x"e1", x"e7", x"e9", x"e8", x"e5", x"e4", 
        x"e1", x"de", x"de", x"de", x"da", x"d5", x"d2", x"d3", x"d6", x"d6", x"d7", x"d8", x"d9", x"d9", x"da", 
        x"db", x"da", x"d9", x"d9", x"d9", x"d9", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", 
        x"db", x"dc", x"db", x"da", x"d9", x"d9", x"da", x"da", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"d9", 
        x"a0", x"a1", x"a2", x"a2", x"a1", x"a0", x"9e", x"9e", x"9e", x"9e", x"9e", x"9f", x"9f", x"9e", x"9e", 
        x"9f", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", 
        x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9d", x"9c", x"9d", x"9f", x"a0", x"a1", 
        x"9f", x"9e", x"9f", x"a0", x"9d", x"9c", x"9e", x"a0", x"9e", x"9f", x"a1", x"9e", x"9e", x"9f", x"a0", 
        x"a0", x"a1", x"a1", x"a0", x"a1", x"a1", x"9f", x"9f", x"a0", x"a1", x"a0", x"a0", x"a1", x"a0", x"a0", 
        x"a0", x"a2", x"a0", x"9f", x"a1", x"a0", x"9f", x"a0", x"a1", x"a1", x"a0", x"a1", x"a1", x"a1", x"a1", 
        x"a1", x"a1", x"a1", x"a3", x"a3", x"a2", x"a2", x"a1", x"a1", x"a1", x"a3", x"a3", x"a2", x"a2", x"a2", 
        x"a2", x"a4", x"93", x"7b", x"9b", x"8d", x"74", x"5b", x"45", x"38", x"31", x"1c", x"0f", x"07", x"06", 
        x"0c", x"1d", x"3b", x"5b", x"76", x"99", x"aa", x"ae", x"6e", x"49", x"39", x"37", x"8f", x"ac", x"ac", 
        x"ac", x"a7", x"a8", x"a3", x"93", x"90", x"97", x"8d", x"60", x"44", x"52", x"50", x"59", x"44", x"3e", 
        x"48", x"6b", x"c2", x"e1", x"d8", x"da", x"d8", x"d9", x"e3", x"d4", x"d5", x"d1", x"d2", x"d3", x"d2", 
        x"d0", x"d0", x"d2", x"d3", x"d3", x"d1", x"cf", x"d0", x"d0", x"d2", x"d3", x"d1", x"d4", x"d9", x"d2", 
        x"b9", x"9d", x"86", x"82", x"92", x"b0", x"ce", x"db", x"da", x"d6", x"d4", x"d3", x"d4", x"d4", x"d1", 
        x"d3", x"d3", x"d3", x"d5", x"d5", x"d3", x"d0", x"d1", x"d2", x"d5", x"da", x"d8", x"d6", x"d7", x"d9", 
        x"d9", x"d3", x"e2", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ed", x"ed", 
        x"ed", x"ee", x"ef", x"f0", x"ee", x"ed", x"ee", x"f0", x"f3", x"f2", x"f3", x"f4", x"ee", x"e8", x"de", 
        x"d2", x"c9", x"c4", x"bd", x"bf", x"be", x"ba", x"c0", x"cd", x"d8", x"dd", x"e2", x"ea", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f1", x"f4", x"f1", x"f1", x"ee", x"ee", x"ef", x"ef", x"ed", x"e9", x"f3", 
        x"f2", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"ed", x"f2", x"f3", 
        x"f3", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"f3", x"f4", x"f4", x"f3", 
        x"f4", x"f4", x"f2", x"f2", x"f1", x"ef", x"ee", x"f0", x"f4", x"f7", x"f5", x"f1", x"e9", x"df", x"d3", 
        x"ca", x"c6", x"c4", x"c2", x"c8", x"d3", x"df", x"e8", x"f0", x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f4", x"f3", x"f2", x"f3", x"f3", x"f4", x"f4", x"f5", x"f5", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f4", 
        x"f2", x"f5", x"f6", x"f6", x"f3", x"f0", x"ee", x"f6", x"f6", x"f5", x"f3", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"ef", x"ef", x"ee", x"f0", x"f3", x"f5", x"f6", x"f6", x"f5", x"f4", x"f4", x"f0", 
        x"98", x"5c", x"6c", x"89", x"de", x"d7", x"da", x"ba", x"9f", x"9e", x"a2", x"9b", x"9b", x"99", x"97", 
        x"96", x"95", x"95", x"94", x"93", x"91", x"91", x"91", x"8f", x"91", x"97", x"97", x"9a", x"96", x"90", 
        x"8b", x"89", x"8d", x"99", x"86", x"60", x"46", x"68", x"78", x"67", x"64", x"68", x"71", x"78", x"7f", 
        x"85", x"88", x"85", x"83", x"83", x"82", x"80", x"7f", x"80", x"81", x"82", x"80", x"7f", x"80", x"82", 
        x"83", x"82", x"82", x"82", x"82", x"9c", x"62", x"60", x"d8", x"e4", x"e0", x"e1", x"e0", x"e0", x"e0", 
        x"e2", x"e2", x"e4", x"e4", x"e4", x"e2", x"e2", x"e3", x"e3", x"e0", x"e1", x"e1", x"df", x"e2", x"df", 
        x"e2", x"e2", x"df", x"dd", x"e1", x"e5", x"e6", x"e5", x"e6", x"e7", x"e5", x"e1", x"dd", x"d9", x"d8", 
        x"d5", x"d3", x"d5", x"d7", x"d8", x"db", x"dd", x"dd", x"db", x"da", x"d9", x"d9", x"d9", x"d8", x"da", 
        x"dc", x"db", x"da", x"da", x"d9", x"d9", x"d9", x"da", x"db", x"db", x"da", x"da", x"da", x"d9", x"d9", 
        x"db", x"dc", x"db", x"da", x"d9", x"da", x"da", x"da", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"d9", 
        x"a2", x"a2", x"a3", x"a2", x"a1", x"9f", x"9f", x"9f", x"9e", x"9d", x"9e", x"a0", x"9f", x"9d", x"9e", 
        x"a1", x"9f", x"9e", x"9e", x"9d", x"9d", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", x"9e", 
        x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"a0", x"a1", x"9f", x"9f", x"9f", x"a0", x"9d", x"9d", 
        x"9e", x"9e", x"a0", x"a2", x"a0", x"9f", x"9f", x"a1", x"9e", x"9f", x"a1", x"9f", x"9f", x"a1", x"a0", 
        x"a0", x"a1", x"a0", x"a1", x"a1", x"a1", x"a0", x"9f", x"9f", x"a0", x"a1", x"a1", x"a1", x"a0", x"9f", 
        x"a0", x"a1", x"a0", x"9f", x"a2", x"a0", x"9f", x"9f", x"a0", x"a1", x"a1", x"a1", x"a1", x"a2", x"a2", 
        x"a1", x"a1", x"a2", x"a3", x"a3", x"a2", x"a2", x"a1", x"a1", x"a1", x"a3", x"a3", x"a0", x"a2", x"a2", 
        x"a2", x"a7", x"94", x"64", x"58", x"4b", x"40", x"34", x"22", x"16", x"09", x"04", x"05", x"12", x"34", 
        x"52", x"75", x"93", x"a5", x"a8", x"aa", x"a9", x"ac", x"73", x"58", x"42", x"38", x"92", x"ab", x"ab", 
        x"ab", x"aa", x"aa", x"a8", x"9c", x"95", x"9e", x"95", x"5e", x"2e", x"2e", x"34", x"4c", x"65", x"80", 
        x"87", x"82", x"c3", x"e1", x"d8", x"d9", x"d5", x"d4", x"e2", x"d4", x"d3", x"cf", x"d1", x"d2", x"d3", 
        x"d3", x"d3", x"d3", x"d1", x"d2", x"d3", x"d1", x"d3", x"d2", x"d6", x"db", x"d6", x"be", x"95", x"7a", 
        x"88", x"9b", x"b4", x"ce", x"d9", x"d6", x"d2", x"d3", x"d0", x"d1", x"d3", x"d3", x"d4", x"d5", x"d3", 
        x"d5", x"d4", x"d2", x"d3", x"d4", x"d2", x"d1", x"d3", x"d3", x"d5", x"da", x"d8", x"d6", x"d8", x"da", 
        x"da", x"d4", x"e2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f1", x"f0", x"f0", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", x"ee", x"ee", x"f0", x"f1", x"ef", x"ef", x"f1", x"f2", 
        x"f1", x"f0", x"ef", x"e9", x"e8", x"e1", x"d6", x"ce", x"c9", x"c3", x"b9", x"b4", x"b4", x"b9", x"c2", 
        x"cf", x"dc", x"e7", x"ef", x"ef", x"f4", x"f1", x"f3", x"ee", x"ed", x"ec", x"ed", x"ee", x"e8", x"f2", 
        x"f2", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"ec", x"f1", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f0", x"ef", 
        x"f0", x"f1", x"f0", x"f0", x"ef", x"f1", x"f4", x"f3", x"f0", x"f1", x"f2", x"f1", x"f2", x"f3", x"f4", 
        x"f5", x"ef", x"e7", x"df", x"d5", x"cc", x"c3", x"ba", x"ba", x"c2", x"d3", x"e5", x"f1", x"f6", x"f5", 
        x"f2", x"f0", x"f1", x"f0", x"f0", x"ef", x"f2", x"f3", x"f4", x"f3", x"f3", x"f5", x"f5", x"f4", x"f5", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f4", 
        x"f2", x"f6", x"f8", x"f6", x"f2", x"f0", x"ef", x"f6", x"f5", x"f3", x"f1", x"f0", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"f3", x"f5", x"f4", x"f5", x"f6", x"f6", x"f6", x"f1", 
        x"a4", x"58", x"6a", x"83", x"df", x"d7", x"d8", x"d2", x"a9", x"a0", x"9d", x"9c", x"9a", x"9a", x"98", 
        x"96", x"95", x"95", x"93", x"91", x"92", x"92", x"92", x"91", x"91", x"96", x"99", x"9d", x"9a", x"90", 
        x"8a", x"88", x"88", x"91", x"84", x"5e", x"4b", x"70", x"8f", x"85", x"80", x"7b", x"74", x"65", x"5a", 
        x"5c", x"65", x"70", x"7e", x"83", x"85", x"82", x"80", x"7e", x"81", x"82", x"82", x"80", x"80", x"80", 
        x"81", x"82", x"7f", x"80", x"83", x"9b", x"6e", x"61", x"d5", x"e6", x"e1", x"e6", x"e8", x"e6", x"e5", 
        x"e4", x"e1", x"e0", x"e3", x"e6", x"e5", x"e3", x"e4", x"e4", x"e2", x"e2", x"e3", x"e3", x"e6", x"e5", 
        x"e7", x"e7", x"e7", x"e7", x"e6", x"e4", x"e1", x"dd", x"d5", x"d5", x"d5", x"d6", x"d6", x"d7", x"d8", 
        x"d7", x"d9", x"d9", x"d8", x"da", x"dd", x"de", x"dd", x"db", x"db", x"db", x"db", x"da", x"d9", x"d8", 
        x"d9", x"d9", x"da", x"da", x"da", x"da", x"da", x"db", x"db", x"db", x"da", x"da", x"da", x"da", x"d8", 
        x"d9", x"db", x"db", x"da", x"da", x"db", x"db", x"db", x"da", x"d9", x"d9", x"d9", x"d9", x"d9", x"d9", 
        x"a3", x"a2", x"a2", x"a1", x"a1", x"a1", x"a0", x"9f", x"9e", x"9d", x"9f", x"a1", x"a0", x"9d", x"9e", 
        x"a1", x"9f", x"9d", x"9f", x"9e", x"9d", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"a0", 
        x"a0", x"a0", x"a0", x"a0", x"a0", x"9f", x"9d", x"9e", x"a0", x"9f", x"9e", x"9e", x"9e", x"9c", x"9d", 
        x"9e", x"9e", x"9f", x"a2", x"a1", x"9f", x"9e", x"9f", x"9d", x"9f", x"a3", x"a0", x"9f", x"a0", x"a0", 
        x"a2", x"a2", x"a1", x"a2", x"a0", x"a1", x"a1", x"a1", x"a0", x"a1", x"a1", x"a2", x"a0", x"9f", x"9f", 
        x"a0", x"a1", x"a0", x"a0", x"a1", x"a1", x"a0", x"9f", x"9f", x"a0", x"a1", x"a1", x"a2", x"a2", x"a2", 
        x"a1", x"a1", x"a2", x"a3", x"a3", x"a2", x"a2", x"a2", x"a3", x"a3", x"a4", x"a2", x"a1", x"a2", x"a2", 
        x"a1", x"a8", x"92", x"4f", x"36", x"2b", x"1e", x"12", x"06", x"03", x"04", x"05", x"0c", x"25", x"61", 
        x"88", x"9b", x"a9", x"ad", x"aa", x"aa", x"ad", x"ae", x"7a", x"62", x"43", x"32", x"8d", x"ac", x"ab", 
        x"ac", x"ac", x"ab", x"ac", x"ab", x"9a", x"7c", x"59", x"38", x"3e", x"5d", x"76", x"85", x"8d", x"87", 
        x"72", x"5f", x"b9", x"e6", x"dc", x"da", x"d9", x"d9", x"e1", x"d2", x"d4", x"d1", x"d2", x"d2", x"d2", 
        x"d2", x"d4", x"d1", x"cf", x"d2", x"d8", x"d5", x"d8", x"d3", x"c2", x"a7", x"88", x"86", x"94", x"a7", 
        x"c3", x"d2", x"d8", x"d9", x"d6", x"d1", x"d1", x"d2", x"d1", x"d1", x"d3", x"d3", x"d3", x"d4", x"d0", 
        x"d2", x"d2", x"d1", x"d3", x"d4", x"d3", x"d3", x"d5", x"d4", x"d5", x"d9", x"d8", x"d9", x"d9", x"da", 
        x"da", x"d3", x"e2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ed", x"ef", x"f0", x"f0", x"f0", 
        x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ed", x"ee", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"f1", x"f1", x"f0", x"f0", x"ed", x"e7", x"e1", x"db", x"d5", x"cf", x"c8", 
        x"c1", x"be", x"b9", x"bb", x"bf", x"cc", x"d2", x"e1", x"e5", x"ea", x"ec", x"ee", x"ef", x"e5", x"f0", 
        x"f3", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f4", x"f4", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f0", x"f0", x"f1", x"f1", x"f2", x"f3", x"f4", x"f2", x"ec", x"f1", x"f3", 
        x"f4", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f0", x"f0", x"ef", x"f0", x"f4", x"f3", x"ef", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f3", x"f4", x"f3", x"f1", x"ef", x"ec", x"e6", x"dd", x"d3", x"ca", x"c2", x"bd", x"be", x"c7", x"d3", 
        x"df", x"ed", x"f0", x"f2", x"f2", x"f2", x"f3", x"f5", x"f6", x"f3", x"f4", x"f6", x"f5", x"f4", x"f4", 
        x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", x"f4", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f3", 
        x"f2", x"f7", x"f9", x"f7", x"f1", x"f0", x"f0", x"f6", x"f5", x"f4", x"f2", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"ed", x"f0", 
        x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f2", x"f5", x"f2", x"f4", x"f6", x"f5", x"f6", x"f3", 
        x"af", x"58", x"66", x"7f", x"e0", x"d8", x"d4", x"db", x"bc", x"a4", x"9c", x"9c", x"9b", x"9d", x"9a", 
        x"96", x"94", x"97", x"96", x"94", x"96", x"93", x"92", x"92", x"8f", x"90", x"97", x"9e", x"9d", x"94", 
        x"90", x"8c", x"88", x"90", x"87", x"61", x"4e", x"6a", x"8c", x"85", x"85", x"85", x"83", x"7e", x"78", 
        x"74", x"6c", x"64", x"5e", x"64", x"6e", x"76", x"81", x"81", x"83", x"80", x"82", x"81", x"81", x"7e", 
        x"7f", x"80", x"7e", x"7e", x"85", x"97", x"74", x"62", x"d2", x"eb", x"e6", x"e7", x"e6", x"e4", x"e5", 
        x"e9", x"e7", x"e4", x"e5", x"e6", x"e4", x"e1", x"e3", x"e6", x"e7", x"e7", x"e7", x"e6", x"e5", x"e4", 
        x"e2", x"e0", x"de", x"dc", x"d8", x"d7", x"d8", x"d9", x"d6", x"d8", x"d7", x"d9", x"d9", x"db", x"dd", 
        x"da", x"dd", x"db", x"d9", x"db", x"db", x"db", x"db", x"dc", x"db", x"da", x"db", x"dc", x"dc", x"db", 
        x"da", x"da", x"db", x"db", x"db", x"db", x"da", x"da", x"da", x"da", x"db", x"db", x"db", x"db", x"da", 
        x"db", x"da", x"db", x"da", x"da", x"d9", x"db", x"da", x"d8", x"d7", x"d7", x"d9", x"da", x"d9", x"d9", 
        x"a2", x"a1", x"a1", x"a1", x"a1", x"a2", x"a2", x"a0", x"9e", x"9d", x"9f", x"a1", x"a0", x"9d", x"9d", 
        x"9f", x"9e", x"9d", x"a0", x"9e", x"9e", x"a0", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"a0", 
        x"9f", x"9f", x"9f", x"9f", x"9f", x"9f", x"9e", x"a0", x"a1", x"a0", x"9f", x"9f", x"9f", x"9e", x"a0", 
        x"a1", x"9e", x"9e", x"9f", x"9f", x"a0", x"a0", x"a0", x"9d", x"9f", x"a2", x"9f", x"9d", x"a0", x"a0", 
        x"a3", x"a4", x"a1", x"a1", x"a0", x"a2", x"a3", x"a3", x"a1", x"a1", x"a2", x"a3", x"a1", x"9f", x"9f", 
        x"a1", x"a2", x"a1", x"a1", x"a1", x"a2", x"a1", x"9f", x"9f", x"a0", x"a2", x"a1", x"a2", x"a3", x"a2", 
        x"a1", x"a1", x"a2", x"a3", x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", x"a5", x"a4", x"a3", x"a3", x"a1", 
        x"a0", x"a7", x"98", x"5d", x"3b", x"2c", x"19", x"0c", x"04", x"05", x"09", x"17", x"3e", x"5f", x"73", 
        x"79", x"7c", x"7d", x"82", x"87", x"8f", x"9c", x"a2", x"77", x"62", x"3e", x"33", x"90", x"b0", x"ad", 
        x"ae", x"b3", x"b3", x"99", x"6d", x"43", x"39", x"53", x"6c", x"85", x"90", x"8f", x"84", x"74", x"54", 
        x"36", x"3a", x"b0", x"e4", x"dc", x"da", x"d9", x"d8", x"df", x"d2", x"d5", x"d3", x"d4", x"d3", x"d1", 
        x"d0", x"d3", x"d3", x"d3", x"d9", x"dd", x"d4", x"b7", x"89", x"77", x"8a", x"ac", x"c8", x"d0", x"d0", 
        x"d3", x"d3", x"d2", x"d5", x"d4", x"d1", x"d4", x"d1", x"d1", x"d1", x"d2", x"d3", x"d2", x"d0", x"d2", 
        x"d4", x"d4", x"d2", x"d3", x"d3", x"d1", x"d3", x"d6", x"d5", x"d6", x"d9", x"d9", x"d9", x"d9", x"d9", 
        x"d9", x"d2", x"e1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ee", x"ef", x"f0", x"f2", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ed", x"f0", x"f0", x"ef", 
        x"f1", x"f2", x"f0", x"ef", x"f2", x"f2", x"ef", x"ef", x"ef", x"ee", x"f1", x"ee", x"ec", x"ec", x"ea", 
        x"e7", x"e5", x"e0", x"da", x"cc", x"c4", x"b6", x"b3", x"ad", x"b1", x"bc", x"cf", x"e3", x"e5", x"f1", 
        x"f3", x"f1", x"f2", x"f2", x"f1", x"ef", x"ee", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f4", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f0", x"f1", x"f1", x"f2", x"f2", x"f3", x"f4", x"f2", x"ec", x"f0", x"f3", 
        x"f4", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", 
        x"f4", x"f3", x"ef", x"f3", x"f3", x"f1", x"f1", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f0", x"f1", 
        x"f3", x"f1", x"f0", x"f0", x"f1", x"f4", x"f4", x"f2", x"f0", x"ef", x"ec", x"e4", x"db", x"cf", x"c3", 
        x"bb", x"b8", x"bf", x"cd", x"df", x"f0", x"f5", x"f6", x"f6", x"f3", x"f4", x"f6", x"f5", x"f3", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", 
        x"f2", x"f7", x"fa", x"f7", x"f0", x"f0", x"ef", x"f4", x"f4", x"f2", x"f1", x"f1", x"f2", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"ed", x"ef", 
        x"f2", x"f1", x"f1", x"f3", x"f1", x"f0", x"ee", x"f2", x"f4", x"f2", x"f4", x"f7", x"f4", x"f5", x"f4", 
        x"b7", x"58", x"62", x"7b", x"df", x"d6", x"d2", x"d7", x"d2", x"a6", x"a0", x"9b", x"9d", x"9f", x"9b", 
        x"96", x"94", x"98", x"99", x"94", x"96", x"93", x"92", x"94", x"91", x"90", x"94", x"9c", x"9d", x"92", 
        x"92", x"91", x"8a", x"8e", x"84", x"5d", x"4d", x"67", x"8d", x"83", x"82", x"85", x"85", x"83", x"82", 
        x"82", x"80", x"7d", x"7b", x"75", x"69", x"56", x"58", x"64", x"78", x"82", x"86", x"85", x"84", x"7e", 
        x"7d", x"7d", x"7c", x"7a", x"83", x"8e", x"6f", x"5c", x"ce", x"ec", x"e7", x"eb", x"ec", x"ea", x"e7", 
        x"e6", x"e4", x"e2", x"e7", x"eb", x"ea", x"e6", x"e6", x"e8", x"e6", x"e2", x"dd", x"d9", x"d3", x"d3", 
        x"d2", x"d7", x"d7", x"d8", x"db", x"dd", x"dc", x"da", x"dd", x"de", x"db", x"dc", x"d9", x"da", x"db", 
        x"d8", x"dc", x"db", x"d9", x"dd", x"dd", x"db", x"dc", x"dc", x"db", x"d9", x"da", x"da", x"da", x"db", 
        x"db", x"db", x"db", x"db", x"db", x"dc", x"db", x"d9", x"d9", x"da", x"db", x"db", x"dc", x"dc", x"da", 
        x"d9", x"d9", x"da", x"db", x"db", x"da", x"dc", x"da", x"d8", x"d6", x"d6", x"d8", x"da", x"d9", x"d9", 
        x"a0", x"a0", x"a0", x"9f", x"9f", x"9f", x"9f", x"a0", x"9f", x"9e", x"9f", x"a1", x"a1", x"9f", x"9e", 
        x"9d", x"9e", x"9e", x"9f", x"9f", x"9f", x"a0", x"a0", x"a0", x"9f", x"9e", x"9f", x"a1", x"a1", x"a0", 
        x"9f", x"9f", x"9e", x"9d", x"9e", x"9e", x"9e", x"9f", x"a0", x"9f", x"9e", x"9e", x"9f", x"a0", x"a1", 
        x"a1", x"a0", x"9e", x"9f", x"a1", x"9f", x"a0", x"a1", x"a0", x"a1", x"a2", x"9f", x"a0", x"a2", x"a1", 
        x"a1", x"a1", x"a2", x"a2", x"a2", x"a1", x"a2", x"a1", x"a0", x"a1", x"a0", x"a0", x"a3", x"a1", x"a1", 
        x"a2", x"a1", x"a2", x"a3", x"a2", x"a3", x"a4", x"a4", x"a3", x"a2", x"a2", x"a3", x"a3", x"a2", x"a1", 
        x"a1", x"a3", x"a5", x"a3", x"a2", x"a3", x"a4", x"a5", x"a6", x"a6", x"a5", x"a3", x"a2", x"a2", x"a2", 
        x"a2", x"a4", x"a4", x"a1", x"9f", x"98", x"94", x"6f", x"1f", x"27", x"5c", x"75", x"7c", x"77", x"75", 
        x"72", x"73", x"71", x"70", x"76", x"65", x"6c", x"6e", x"5e", x"5f", x"3b", x"37", x"81", x"9c", x"a4", 
        x"99", x"85", x"65", x"51", x"6d", x"86", x"7f", x"8b", x"8b", x"87", x"76", x"5f", x"3f", x"2e", x"34", 
        x"3e", x"4c", x"ba", x"e4", x"d7", x"d8", x"da", x"d9", x"e3", x"d6", x"d5", x"d1", x"d2", x"d1", x"d0", 
        x"d3", x"d2", x"da", x"d3", x"bd", x"99", x"7d", x"82", x"a7", x"c4", x"d4", x"d3", x"d4", x"d6", x"d3", 
        x"d4", x"d4", x"d5", x"d5", x"d3", x"d2", x"d2", x"d1", x"d1", x"d1", x"d2", x"d3", x"d3", x"d3", x"d2", 
        x"d1", x"d3", x"d5", x"d5", x"d4", x"d3", x"d2", x"d3", x"d3", x"d4", x"da", x"d8", x"d8", x"d9", x"da", 
        x"d9", x"d5", x"df", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ed", x"ed", 
        x"ee", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", 
        x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ea", x"e5", x"e0", x"d8", x"cd", x"c4", x"ca", x"bf", x"b4", 
        x"b8", x"c1", x"d3", x"dc", x"e5", x"ea", x"ed", x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f0", x"f1", x"ef", x"f0", x"f0", x"ed", x"ef", x"f3", x"f2", x"f1", x"f2", x"f3", x"f1", x"f0", 
        x"f3", x"f3", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f3", x"f4", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"ee", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", 
        x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"ee", x"ec", 
        x"e8", x"e0", x"d3", x"c8", x"c2", x"c4", x"c9", x"d0", x"df", x"e6", x"ee", x"f1", x"f2", x"f2", x"f4", 
        x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f1", x"f2", x"f3", x"f3", x"f4", x"f5", x"f4", x"f3", x"f4", 
        x"f7", x"f8", x"f8", x"f6", x"f4", x"f1", x"f1", x"f4", x"f5", x"f2", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"ef", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f0", x"f0", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f1", x"f5", x"f5", x"f4", x"f6", x"f6", x"f5", x"f4", 
        x"be", x"54", x"62", x"77", x"dd", x"d6", x"d4", x"d5", x"d9", x"bc", x"9d", x"a0", x"9e", x"9f", x"99", 
        x"98", x"97", x"96", x"99", x"94", x"96", x"94", x"91", x"91", x"91", x"92", x"93", x"99", x"9d", x"94", 
        x"95", x"95", x"8c", x"8d", x"86", x"5f", x"4f", x"62", x"90", x"83", x"86", x"85", x"84", x"81", x"82", 
        x"7f", x"7d", x"7e", x"7f", x"7f", x"81", x"80", x"79", x"6b", x"5f", x"54", x"56", x"63", x"71", x"79", 
        x"7f", x"82", x"81", x"7c", x"87", x"97", x"81", x"5d", x"c5", x"ef", x"e8", x"e6", x"e9", x"ea", x"e9", 
        x"e8", x"e7", x"e4", x"e5", x"e2", x"e0", x"db", x"dc", x"d9", x"d5", x"d4", x"d3", x"d3", x"d5", x"d8", 
        x"d9", x"db", x"da", x"db", x"dd", x"de", x"de", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", 
        x"d9", x"dc", x"da", x"da", x"dd", x"db", x"da", x"dc", x"db", x"da", x"d9", x"d9", x"d9", x"d9", x"da", 
        x"da", x"da", x"db", x"db", x"db", x"dc", x"db", x"da", x"da", x"db", x"dc", x"db", x"db", x"da", x"d9", 
        x"d9", x"d9", x"da", x"da", x"da", x"da", x"db", x"da", x"d9", x"d8", x"d9", x"d7", x"d6", x"d7", x"d8", 
        x"a2", x"a2", x"a1", x"a0", x"9f", x"9e", x"9e", x"9e", x"9e", x"9f", x"9f", x"9e", x"9e", x"9f", x"a0", 
        x"a0", x"a1", x"a1", x"a1", x"a1", x"a1", x"9f", x"9e", x"9e", x"9e", x"9d", x"9e", x"9f", x"a1", x"9f", 
        x"9f", x"a0", x"9f", x"9e", x"9d", x"9d", x"9f", x"a0", x"a0", x"9f", x"9e", x"9e", x"9f", x"a0", x"a1", 
        x"a1", x"a0", x"a0", x"a0", x"a1", x"a0", x"a1", x"a1", x"9f", x"9f", x"a1", x"a0", x"a1", x"a2", x"a1", 
        x"a1", x"a1", x"a1", x"a2", x"a2", x"a0", x"a2", x"a1", x"a1", x"a2", x"a3", x"a2", x"a3", x"a1", x"a2", 
        x"a2", x"a1", x"a2", x"a3", x"a1", x"a2", x"a3", x"a2", x"a1", x"a2", x"a2", x"a4", x"a4", x"a4", x"a3", 
        x"a3", x"a3", x"a4", x"a3", x"a2", x"a2", x"a2", x"a3", x"a5", x"a5", x"a2", x"9f", x"a0", x"a2", x"a4", 
        x"a5", x"a6", x"a4", x"a2", x"a8", x"a5", x"ae", x"8e", x"33", x"53", x"a6", x"b0", x"a7", x"9d", x"96", 
        x"8b", x"85", x"78", x"75", x"76", x"69", x"6c", x"68", x"62", x"65", x"40", x"3a", x"68", x"5b", x"4e", 
        x"41", x"55", x"87", x"bd", x"d7", x"bf", x"87", x"7f", x"6e", x"4f", x"38", x"2e", x"36", x"48", x"5f", 
        x"68", x"6a", x"c2", x"e2", x"d9", x"db", x"db", x"d6", x"e1", x"d4", x"d4", x"d3", x"d2", x"d2", x"d5", 
        x"d5", x"c5", x"a8", x"83", x"76", x"97", x"c0", x"d5", x"da", x"d6", x"d1", x"d0", x"d3", x"d5", x"d1", 
        x"d3", x"d3", x"d4", x"d3", x"d2", x"d1", x"d1", x"d1", x"d1", x"d1", x"d3", x"d4", x"d4", x"d3", x"d3", 
        x"d2", x"d3", x"d5", x"d4", x"d3", x"d3", x"d2", x"d1", x"d2", x"d3", x"db", x"d9", x"d8", x"d8", x"da", 
        x"db", x"d6", x"de", x"f1", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ed", x"ed", 
        x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", 
        x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ed", x"ef", x"ee", x"ec", x"de", x"d4", 
        x"ca", x"b7", x"ab", x"aa", x"ab", x"b3", x"bf", x"cc", x"d8", x"e5", x"e8", x"ec", x"ef", x"f1", x"f1", 
        x"ef", x"ee", x"ee", x"ec", x"ee", x"f0", x"ee", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f0", x"ef", x"f0", x"f0", x"ef", x"f1", x"f2", x"f0", x"ee", x"ef", 
        x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f1", x"e5", x"d5", x"c9", x"be", x"bf", x"c4", x"cd", x"da", x"e5", x"ed", 
        x"f1", x"f3", x"f3", x"f5", x"f6", x"f4", x"f1", x"f4", x"f5", x"f4", x"f3", x"f4", x"f4", x"f5", x"f5", 
        x"f6", x"f7", x"f9", x"f8", x"f4", x"ef", x"ed", x"f1", x"f3", x"f2", x"f0", x"f0", x"f0", x"ef", x"f1", 
        x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f1", x"f5", x"f5", x"f4", x"f5", x"f6", x"f5", x"f5", 
        x"c3", x"56", x"62", x"75", x"da", x"d5", x"d4", x"d5", x"da", x"c4", x"9e", x"a3", x"9e", x"9e", x"99", 
        x"98", x"98", x"96", x"98", x"95", x"97", x"95", x"92", x"91", x"92", x"93", x"93", x"97", x"9d", x"96", 
        x"96", x"98", x"8f", x"8e", x"89", x"64", x"52", x"60", x"8f", x"82", x"87", x"86", x"85", x"83", x"84", 
        x"81", x"7c", x"7c", x"7b", x"7c", x"7d", x"7e", x"80", x"81", x"81", x"7d", x"6e", x"60", x"56", x"56", 
        x"5d", x"67", x"78", x"81", x"81", x"8f", x"7f", x"6d", x"cf", x"f2", x"eb", x"e8", x"e4", x"e0", x"dc", 
        x"da", x"d8", x"d4", x"d6", x"d4", x"d6", x"d5", x"d6", x"d9", x"df", x"dd", x"db", x"db", x"db", x"dc", 
        x"dd", x"dc", x"db", x"db", x"dd", x"de", x"de", x"dd", x"db", x"db", x"db", x"db", x"dc", x"dc", x"db", 
        x"da", x"dc", x"da", x"da", x"dd", x"da", x"da", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dd", x"dd", 
        x"dc", x"db", x"db", x"db", x"da", x"da", x"db", x"dc", x"dd", x"dd", x"dd", x"dd", x"dc", x"db", x"da", 
        x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"d8", x"d7", x"d6", x"d7", 
        x"a3", x"a2", x"a2", x"a1", x"a0", x"a0", x"9f", x"a0", x"a1", x"a3", x"a2", x"a0", x"9f", x"a1", x"a2", 
        x"a1", x"a1", x"a1", x"a1", x"a0", x"a0", x"9f", x"9f", x"a0", x"a0", x"9f", x"a0", x"a1", x"a2", x"9f", 
        x"a0", x"a1", x"a0", x"9f", x"9e", x"9e", x"9f", x"a0", x"a1", x"a0", x"9f", x"9f", x"a0", x"a0", x"a1", 
        x"a0", x"a1", x"a1", x"a1", x"a0", x"a1", x"a2", x"a0", x"9e", x"9f", x"a1", x"a1", x"a1", x"a1", x"a1", 
        x"a1", x"a1", x"a1", x"a1", x"a3", x"a3", x"a4", x"a2", x"a1", x"a2", x"a3", x"a2", x"a3", x"a1", x"a1", 
        x"a2", x"a1", x"a2", x"a3", x"a3", x"a4", x"a4", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", x"a4", x"a4", 
        x"a2", x"a2", x"a1", x"a2", x"a2", x"a1", x"a1", x"a1", x"a3", x"a4", x"a3", x"a1", x"a2", x"a3", x"a4", 
        x"a4", x"a4", x"a3", x"a2", x"a4", x"a4", x"ab", x"88", x"34", x"57", x"9c", x"ab", x"a9", x"ac", x"ae", 
        x"ab", x"ab", x"a8", x"a3", x"9f", x"99", x"95", x"8c", x"6e", x"60", x"3f", x"33", x"4d", x"4c", x"6f", 
        x"a2", x"c2", x"d0", x"d5", x"c8", x"97", x"5c", x"44", x"33", x"35", x"46", x"59", x"69", x"72", x"7a", 
        x"7a", x"7a", x"c2", x"e1", x"d8", x"d9", x"d9", x"d5", x"e1", x"d8", x"d9", x"d8", x"d2", x"c2", x"ac", 
        x"9a", x"8a", x"92", x"ae", x"ca", x"d7", x"d4", x"d1", x"d3", x"d1", x"d3", x"d4", x"d2", x"d3", x"d1", 
        x"d1", x"d2", x"d3", x"d3", x"d2", x"d0", x"d1", x"d2", x"d1", x"d1", x"d3", x"d5", x"d5", x"d2", x"d3", 
        x"d3", x"d5", x"d5", x"d3", x"d2", x"d3", x"d3", x"d1", x"d0", x"d3", x"dc", x"da", x"d7", x"d7", x"db", 
        x"db", x"d5", x"dd", x"f1", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"ef", x"ed", x"ed", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f1", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ec", x"e7", x"ee", 
        x"f0", x"ed", x"e8", x"e2", x"d9", x"cf", x"c5", x"bc", x"b7", x"ba", x"bc", x"c2", x"cb", x"d4", x"da", 
        x"dd", x"e5", x"ea", x"eb", x"ee", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"ef", x"ef", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f1", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f2", x"f2", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f4", x"f3", x"f2", x"f2", x"f3", x"f4", x"f2", x"f0", x"ee", x"e6", x"da", x"ce", x"c7", x"c7", x"c9", 
        x"cc", x"d4", x"dd", x"e6", x"ec", x"f0", x"f3", x"f4", x"f4", x"f5", x"f3", x"f1", x"f2", x"f3", x"f6", 
        x"f7", x"f6", x"f6", x"f7", x"f6", x"f2", x"ef", x"f0", x"f3", x"f3", x"f2", x"f2", x"f1", x"f0", x"f2", 
        x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f1", x"f5", x"f5", x"f4", x"f5", x"f5", x"f4", x"f5", 
        x"ca", x"59", x"63", x"72", x"d8", x"d6", x"d4", x"d5", x"da", x"c6", x"9e", x"a1", x"9d", x"9d", x"99", 
        x"98", x"97", x"96", x"97", x"96", x"97", x"96", x"93", x"92", x"93", x"93", x"93", x"95", x"9d", x"99", 
        x"97", x"9a", x"94", x"8f", x"8b", x"67", x"53", x"5b", x"8c", x"85", x"89", x"87", x"86", x"83", x"85", 
        x"82", x"7d", x"7b", x"7b", x"7d", x"7c", x"7b", x"79", x"7a", x"7c", x"7e", x"7f", x"7d", x"78", x"70", 
        x"69", x"64", x"60", x"58", x"6e", x"9e", x"9b", x"91", x"d0", x"d9", x"d4", x"d2", x"cc", x"c8", x"cb", 
        x"cf", x"d4", x"d7", x"d9", x"da", x"dc", x"dd", x"de", x"dd", x"dd", x"dc", x"db", x"da", x"da", x"db", 
        x"db", x"dd", x"dc", x"dc", x"dd", x"de", x"de", x"dd", x"db", x"db", x"db", x"db", x"dc", x"dc", x"dc", 
        x"dc", x"dd", x"db", x"db", x"dc", x"db", x"db", x"dc", x"dc", x"dc", x"dc", x"dc", x"dd", x"de", x"de", 
        x"dc", x"dc", x"db", x"db", x"da", x"da", x"da", x"dc", x"dc", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", 
        x"db", x"db", x"db", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"d8", x"d8", x"d9", x"da", x"d6", x"d5", 
        x"a2", x"a2", x"a2", x"a2", x"a2", x"a2", x"a2", x"a2", x"a2", x"a2", x"a2", x"a2", x"a1", x"a2", x"a1", 
        x"a0", x"a0", x"9f", x"9f", x"9e", x"9e", x"9e", x"9f", x"a1", x"a1", x"a0", x"a0", x"a1", x"a2", x"a0", 
        x"a0", x"a0", x"a0", x"a0", x"9f", x"9f", x"a1", x"a1", x"a1", x"a1", x"a1", x"a1", x"a1", x"a2", x"a1", 
        x"a1", x"a2", x"a3", x"a2", x"a0", x"a2", x"a2", x"a1", x"a0", x"a0", x"a1", x"a2", x"a2", x"a1", x"a1", 
        x"a2", x"a2", x"a1", x"a1", x"a3", x"a4", x"a3", x"a2", x"a1", x"a1", x"a3", x"a3", x"a2", x"a2", x"a2", 
        x"a2", x"a2", x"a2", x"a2", x"a3", x"a4", x"a5", x"a4", x"a4", x"a3", x"a4", x"a3", x"a3", x"a3", x"a3", 
        x"a3", x"a2", x"a2", x"a2", x"a3", x"a2", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", x"a4", x"a4", x"a3", 
        x"a3", x"a3", x"a3", x"a1", x"a0", x"a7", x"ae", x"8c", x"4c", x"6c", x"9a", x"aa", x"a9", x"a9", x"ab", 
        x"aa", x"a9", x"ac", x"a7", x"a3", x"ac", x"b3", x"b2", x"73", x"55", x"45", x"4e", x"88", x"ba", x"e0", 
        x"e0", x"d2", x"bb", x"98", x"68", x"36", x"2f", x"3c", x"48", x"61", x"6f", x"7b", x"7f", x"80", x"82", 
        x"7d", x"7c", x"c2", x"e3", x"d7", x"d6", x"d9", x"d6", x"e4", x"d9", x"d1", x"bb", x"9d", x"86", x"84", 
        x"a3", x"c5", x"dc", x"dc", x"d4", x"cf", x"d0", x"cf", x"d0", x"cf", x"d2", x"d3", x"d1", x"d2", x"cf", 
        x"cf", x"d0", x"d2", x"d2", x"d1", x"d0", x"d0", x"d3", x"d1", x"d0", x"d3", x"d6", x"d5", x"d3", x"d3", 
        x"d4", x"d5", x"d6", x"d2", x"d1", x"d2", x"d3", x"d1", x"d0", x"d3", x"dc", x"da", x"d7", x"d6", x"db", 
        x"dc", x"d4", x"db", x"f1", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"f0", x"eb", x"ef", 
        x"ed", x"ee", x"eb", x"ee", x"f2", x"f4", x"f3", x"f1", x"ee", x"e5", x"d9", x"c8", x"bd", x"b7", x"b2", 
        x"b1", x"b6", x"bd", x"c7", x"d1", x"db", x"e3", x"e8", x"eb", x"ef", x"f2", x"f3", x"f2", x"f1", x"f0", 
        x"ef", x"f2", x"f3", x"f0", x"ee", x"f1", x"f1", x"f2", x"f2", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f1", x"f0", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f0", x"f1", x"f4", x"f7", x"f3", x"eb", x"e2", 
        x"cf", x"c8", x"c3", x"c2", x"c9", x"d3", x"dd", x"e5", x"ea", x"f0", x"f3", x"f4", x"f5", x"f8", x"f9", 
        x"f8", x"f7", x"f6", x"f6", x"f4", x"f1", x"ee", x"ed", x"f2", x"f2", x"f0", x"f0", x"f1", x"f0", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f1", x"f5", x"f5", x"f4", x"f5", x"f6", x"f5", x"f6", 
        x"d1", x"5b", x"62", x"6e", x"d5", x"d8", x"d5", x"d6", x"d9", x"c7", x"9c", x"9e", x"9c", x"9c", x"9a", 
        x"98", x"97", x"96", x"96", x"96", x"98", x"96", x"94", x"93", x"94", x"93", x"93", x"92", x"9a", x"9a", 
        x"98", x"9d", x"99", x"91", x"8d", x"66", x"4d", x"4d", x"82", x"81", x"87", x"87", x"86", x"83", x"84", 
        x"83", x"7c", x"7a", x"7c", x"7a", x"79", x"79", x"78", x"77", x"76", x"7a", x"80", x"80", x"80", x"81", 
        x"83", x"7e", x"6b", x"6c", x"9f", x"c7", x"bc", x"b6", x"c1", x"c3", x"c8", x"cf", x"d2", x"d6", x"dd", 
        x"e1", x"e0", x"e0", x"e0", x"e0", x"e0", x"df", x"de", x"dd", x"dd", x"dc", x"dc", x"dd", x"dd", x"de", 
        x"de", x"dd", x"dc", x"dc", x"dd", x"de", x"de", x"dd", x"dc", x"db", x"db", x"db", x"dc", x"dd", x"dc", 
        x"dd", x"dc", x"db", x"db", x"db", x"dc", x"dc", x"dc", x"db", x"db", x"da", x"da", x"db", x"db", x"dc", 
        x"db", x"db", x"db", x"db", x"db", x"db", x"da", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"dc", 
        x"dc", x"dc", x"db", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"d8", x"d7", x"d8", x"da", x"d6", x"d6", 
        x"a3", x"a3", x"a2", x"a2", x"a1", x"a1", x"a1", x"a1", x"9f", x"9e", x"9f", x"a2", x"a2", x"a0", x"a0", 
        x"a2", x"a2", x"a2", x"a1", x"a0", x"a0", x"9f", x"9d", x"9f", x"a0", x"9f", x"9e", x"9f", x"a0", x"a0", 
        x"a0", x"a0", x"9f", x"a0", x"a1", x"a2", x"a2", x"a1", x"a1", x"a1", x"a2", x"a2", x"a1", x"a2", x"a1", 
        x"a1", x"a2", x"a3", x"a2", x"a1", x"a1", x"a1", x"a1", x"a2", x"a2", x"a1", x"a1", x"a2", x"a2", x"a2", 
        x"a2", x"a2", x"a2", x"a2", x"a3", x"a1", x"a0", x"a1", x"a1", x"a1", x"a3", x"a4", x"a2", x"a3", x"a2", 
        x"a2", x"a3", x"a3", x"a2", x"a1", x"a3", x"a5", x"a4", x"a3", x"a2", x"a1", x"a2", x"a2", x"a2", x"a2", 
        x"a3", x"a3", x"a4", x"a3", x"a4", x"a4", x"a5", x"a5", x"a5", x"a4", x"a4", x"a3", x"a3", x"a2", x"a3", 
        x"a4", x"a5", x"a5", x"a6", x"a5", x"a4", x"ab", x"8a", x"54", x"77", x"9f", x"ac", x"a9", x"a9", x"a8", 
        x"a8", x"a9", x"a9", x"a9", x"a5", x"a7", x"9b", x"97", x"7b", x"85", x"ac", x"ce", x"df", x"d9", x"c1", 
        x"9b", x"75", x"50", x"3c", x"38", x"45", x"5e", x"69", x"76", x"7f", x"81", x"82", x"83", x"85", x"86", 
        x"7e", x"7a", x"be", x"e0", x"da", x"de", x"dc", x"c9", x"b6", x"9f", x"92", x"98", x"a8", x"c2", x"d3", 
        x"d9", x"d8", x"d2", x"d2", x"d2", x"d1", x"d2", x"d1", x"d2", x"d0", x"d0", x"d2", x"d2", x"d2", x"ce", 
        x"cf", x"d0", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d1", x"d0", x"d3", x"d5", x"d4", x"d2", x"d3", 
        x"d3", x"d5", x"d5", x"d2", x"d2", x"d3", x"d3", x"d1", x"d1", x"d3", x"dc", x"d9", x"d7", x"d6", x"da", 
        x"dc", x"d3", x"da", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"ef", x"f1", x"ee", x"e7", x"f1", 
        x"ef", x"ed", x"ec", x"ee", x"ee", x"ec", x"eb", x"eb", x"ee", x"f1", x"f1", x"f0", x"f0", x"ee", x"e8", 
        x"e1", x"d4", x"cc", x"c4", x"bc", x"b8", x"b8", x"b9", x"ba", x"be", x"c7", x"d3", x"de", x"e6", x"ee", 
        x"f2", x"f5", x"f6", x"f3", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f2", x"f1", x"f2", x"f3", x"f3", x"f4", x"f4", 
        x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", 
        x"f3", x"f1", x"ec", x"e2", x"d7", x"cf", x"ca", x"c8", x"c8", x"cc", x"d0", x"d9", x"e7", x"f4", x"f7", 
        x"f7", x"f7", x"f7", x"f6", x"f4", x"f2", x"ef", x"ef", x"f3", x"f3", x"f0", x"f1", x"f3", x"f2", x"f1", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f1", x"f5", x"f5", x"f4", x"f5", x"f7", x"f6", x"f6", 
        x"d7", x"5e", x"62", x"6b", x"d2", x"d8", x"d4", x"d6", x"d9", x"cb", x"9e", x"9e", x"9d", x"9c", x"9c", 
        x"9a", x"98", x"98", x"96", x"96", x"97", x"96", x"94", x"94", x"94", x"92", x"92", x"90", x"96", x"99", 
        x"98", x"9d", x"9c", x"91", x"8c", x"67", x"4e", x"4a", x"83", x"88", x"89", x"87", x"86", x"82", x"84", 
        x"83", x"7b", x"78", x"79", x"76", x"76", x"77", x"78", x"77", x"75", x"77", x"7e", x"7e", x"7e", x"80", 
        x"83", x"7a", x"90", x"b6", x"cb", x"c7", x"ce", x"d4", x"da", x"dd", x"df", x"df", x"dd", x"de", x"df", 
        x"de", x"de", x"df", x"df", x"df", x"de", x"de", x"dd", x"dd", x"df", x"df", x"de", x"dd", x"dd", x"dd", 
        x"dd", x"dd", x"dc", x"dc", x"dd", x"de", x"de", x"dd", x"dc", x"db", x"db", x"dc", x"dd", x"dd", x"dd", 
        x"dd", x"dc", x"dc", x"dc", x"db", x"dc", x"dd", x"dd", x"dd", x"dc", x"db", x"da", x"da", x"da", x"db", 
        x"da", x"da", x"da", x"db", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", 
        x"dc", x"db", x"db", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"d8", x"d7", x"d7", x"d8", x"d9", x"d9", 
        x"a4", x"a4", x"a3", x"a2", x"a1", x"a0", x"a0", x"a2", x"a1", x"a0", x"a1", x"a2", x"a3", x"a1", x"a1", 
        x"a1", x"a2", x"a2", x"a2", x"a1", x"a1", x"a0", x"9f", x"a0", x"a1", x"a1", x"a0", x"a0", x"a1", x"a0", 
        x"a0", x"a0", x"a0", x"a1", x"a1", x"a2", x"a2", x"a1", x"a0", x"a1", x"a2", x"a2", x"a1", x"a1", x"a2", 
        x"a2", x"a2", x"a2", x"a2", x"a1", x"a2", x"a1", x"a2", x"a4", x"a3", x"a1", x"a1", x"a3", x"a2", x"a2", 
        x"a2", x"a2", x"a2", x"a2", x"a4", x"a2", x"a1", x"a2", x"a2", x"a0", x"a1", x"a3", x"a3", x"a4", x"a4", 
        x"a3", x"a4", x"a4", x"a2", x"a2", x"a5", x"a6", x"a6", x"a5", x"a4", x"a3", x"a2", x"a2", x"a2", x"a3", 
        x"a3", x"a3", x"a3", x"a4", x"a4", x"a5", x"a5", x"a5", x"a5", x"a4", x"a4", x"a4", x"a3", x"a3", x"a3", 
        x"a4", x"a5", x"a4", x"a3", x"a6", x"a1", x"a9", x"88", x"52", x"76", x"9f", x"ad", x"ab", x"ac", x"a8", 
        x"a8", x"aa", x"a8", x"a2", x"93", x"98", x"9d", x"ad", x"c2", x"d2", x"de", x"d1", x"aa", x"88", x"62", 
        x"46", x"3d", x"41", x"53", x"62", x"71", x"7f", x"7f", x"84", x"84", x"86", x"86", x"86", x"86", x"88", 
        x"81", x"78", x"c2", x"e6", x"d0", x"bf", x"ad", x"a1", x"a1", x"a0", x"b3", x"d0", x"dc", x"dc", x"d2", 
        x"d1", x"d8", x"d4", x"d2", x"d4", x"d4", x"d4", x"d3", x"d6", x"d1", x"d0", x"d1", x"d2", x"d2", x"ce", 
        x"d0", x"d0", x"d1", x"d1", x"d2", x"d2", x"d2", x"d1", x"d0", x"d0", x"d2", x"d4", x"d3", x"d3", x"d3", 
        x"d2", x"d3", x"d5", x"d4", x"d2", x"d3", x"d4", x"d2", x"d2", x"d3", x"db", x"d8", x"d6", x"d5", x"da", 
        x"db", x"d4", x"da", x"ef", x"f0", x"f0", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"ed", x"e6", x"f0", 
        x"f1", x"ef", x"ed", x"ee", x"ef", x"ed", x"ec", x"ec", x"ed", x"f1", x"f0", x"ee", x"ef", x"f0", x"f2", 
        x"f2", x"f4", x"f3", x"f0", x"e8", x"de", x"d7", x"ce", x"c3", x"bc", x"b8", x"b8", x"b8", x"ba", x"be", 
        x"c5", x"cf", x"d8", x"e2", x"e9", x"ee", x"f1", x"f1", x"f0", x"f2", x"f0", x"ef", x"f0", x"f3", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f3", x"f3", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f7", x"f5", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f0", x"e6", x"dd", x"d3", x"ca", x"c8", x"cc", x"d3", x"d8", 
        x"de", x"e8", x"f1", x"f4", x"f4", x"f2", x"ef", x"ef", x"f4", x"f4", x"f1", x"f1", x"f3", x"f2", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f1", x"f5", x"f5", x"f4", x"f5", x"f7", x"f7", x"f6", 
        x"dd", x"60", x"62", x"68", x"cf", x"d8", x"d4", x"d6", x"d9", x"cf", x"a0", x"9e", x"9e", x"9c", x"9d", 
        x"9b", x"98", x"98", x"96", x"96", x"97", x"96", x"95", x"95", x"94", x"91", x"91", x"90", x"93", x"96", 
        x"97", x"9b", x"9e", x"94", x"90", x"6a", x"4f", x"46", x"81", x"88", x"88", x"87", x"87", x"83", x"84", 
        x"84", x"7b", x"78", x"7c", x"7b", x"7a", x"79", x"78", x"79", x"78", x"79", x"7f", x"80", x"80", x"80", 
        x"81", x"71", x"bb", x"e4", x"e1", x"e1", x"e1", x"de", x"dd", x"dd", x"dd", x"dd", x"de", x"e0", x"e0", 
        x"de", x"dd", x"df", x"de", x"e0", x"df", x"e1", x"e0", x"e0", x"de", x"de", x"de", x"dd", x"dd", x"dd", 
        x"dd", x"dd", x"dc", x"dc", x"de", x"df", x"df", x"de", x"dc", x"dc", x"dc", x"dc", x"dd", x"dd", x"dd", 
        x"dd", x"db", x"dd", x"dd", x"db", x"dc", x"dd", x"dd", x"dd", x"dd", x"dc", x"db", x"db", x"dc", x"dc", 
        x"da", x"da", x"da", x"db", x"dc", x"dc", x"dc", x"dd", x"dd", x"dc", x"dc", x"dc", x"dd", x"dd", x"db", 
        x"db", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"d9", x"d8", x"d9", 
        x"a2", x"a2", x"a2", x"a2", x"a1", x"a1", x"a1", x"a1", x"a1", x"a2", x"a2", x"a0", x"a0", x"a2", x"a0", 
        x"9e", x"9f", x"9f", x"9f", x"a0", x"a0", x"9f", x"9e", x"a0", x"a1", x"a0", x"9f", x"9f", x"9f", x"9f", 
        x"a0", x"a1", x"a2", x"a2", x"a2", x"a1", x"a2", x"a1", x"a0", x"a1", x"a2", x"a2", x"a1", x"a1", x"a2", 
        x"a2", x"a1", x"a0", x"a1", x"a2", x"a3", x"a1", x"a1", x"a3", x"a3", x"a1", x"a1", x"a4", x"a4", x"a3", 
        x"a2", x"a2", x"a3", x"a4", x"a4", x"a1", x"a1", x"a4", x"a5", x"a2", x"a1", x"a3", x"a3", x"a5", x"a4", 
        x"a4", x"a5", x"a5", x"a2", x"a3", x"a4", x"a5", x"a4", x"a3", x"a3", x"a4", x"a2", x"a2", x"a4", x"a4", 
        x"a4", x"a2", x"a1", x"a3", x"a4", x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", x"a5", x"a5", x"a4", 
        x"a4", x"a3", x"a4", x"a3", x"a4", x"a4", x"a8", x"88", x"55", x"79", x"a0", x"ad", x"a8", x"ac", x"ae", 
        x"a9", x"9c", x"8f", x"94", x"a0", x"bc", x"cd", x"da", x"db", x"bf", x"9a", x"6b", x"44", x"3d", x"40", 
        x"4f", x"5a", x"5f", x"77", x"90", x"8a", x"89", x"88", x"87", x"86", x"87", x"88", x"85", x"85", x"87", 
        x"83", x"7c", x"b1", x"b4", x"8f", x"99", x"b0", x"c4", x"dd", x"d7", x"d6", x"d7", x"d3", x"d5", x"d4", 
        x"cf", x"d6", x"d1", x"d1", x"d3", x"d2", x"d2", x"d1", x"d2", x"cf", x"d2", x"d3", x"d2", x"d1", x"ce", 
        x"d1", x"d1", x"d1", x"d1", x"d2", x"d4", x"d4", x"d0", x"d0", x"d0", x"d1", x"d2", x"d3", x"d3", x"d3", 
        x"d1", x"d2", x"d5", x"d5", x"d4", x"d3", x"d4", x"d3", x"d4", x"d4", x"da", x"d7", x"d5", x"d6", x"d9", 
        x"da", x"d4", x"da", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f1", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f2", x"f2", x"ef", x"e8", x"ef", 
        x"f0", x"ed", x"ed", x"ec", x"ed", x"ef", x"ef", x"ee", x"ee", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f0", x"ef", x"f0", x"ef", x"ef", x"f3", x"f2", x"f1", x"ee", x"e8", x"e0", x"d8", x"d1", x"c9", 
        x"bf", x"b7", x"b1", x"ac", x"ac", x"b2", x"be", x"cc", x"db", x"e9", x"f3", x"f5", x"f7", x"f6", x"f3", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", 
        x"f2", x"f3", x"f3", x"f2", x"f0", x"f1", x"f2", x"f3", x"f5", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f5", x"f5", x"f3", x"f0", x"ea", x"e2", x"da", x"d5", 
        x"d3", x"d0", x"ce", x"ce", x"d6", x"e1", x"e8", x"ee", x"f5", x"f5", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"f1", x"f5", x"f5", x"f4", x"f5", x"f6", x"f6", x"f7", 
        x"e2", x"63", x"62", x"65", x"cd", x"da", x"d5", x"d7", x"d8", x"cf", x"9f", x"9c", x"9d", x"9c", x"9f", 
        x"9c", x"98", x"99", x"96", x"96", x"96", x"95", x"95", x"95", x"94", x"91", x"91", x"91", x"90", x"93", 
        x"96", x"98", x"9d", x"9b", x"99", x"6f", x"50", x"41", x"7d", x"85", x"87", x"89", x"89", x"84", x"86", 
        x"86", x"7d", x"78", x"7b", x"7a", x"79", x"78", x"78", x"78", x"78", x"79", x"7f", x"82", x"82", x"81", 
        x"81", x"6a", x"bf", x"e4", x"dd", x"dd", x"de", x"de", x"dd", x"e0", x"df", x"dd", x"de", x"de", x"de", 
        x"df", x"e1", x"e1", x"df", x"e0", x"dd", x"e0", x"de", x"df", x"de", x"de", x"dd", x"dd", x"dd", x"dc", 
        x"dd", x"dd", x"dd", x"dd", x"de", x"df", x"df", x"de", x"dc", x"dc", x"dc", x"dc", x"dd", x"dd", x"dd", 
        x"dc", x"da", x"dd", x"dd", x"db", x"dd", x"dc", x"db", x"dc", x"dc", x"dc", x"dc", x"dd", x"dd", x"dd", 
        x"db", x"db", x"db", x"db", x"db", x"da", x"db", x"dc", x"db", x"da", x"da", x"da", x"db", x"db", x"d9", 
        x"d9", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"dc", x"de", x"de", x"dd", x"d8", x"d1", 
        x"a4", x"a2", x"a3", x"a2", x"a2", x"a4", x"a2", x"a0", x"a3", x"a2", x"a1", x"a2", x"a0", x"a3", x"a2", 
        x"a0", x"a0", x"9f", x"9f", x"a0", x"a0", x"a0", x"9f", x"a0", x"a0", x"a0", x"a1", x"a1", x"a1", x"a0", 
        x"a1", x"a2", x"a3", x"a3", x"a2", x"a1", x"a1", x"a2", x"9f", x"9f", x"a0", x"9f", x"a0", x"a3", x"a2", 
        x"a0", x"a0", x"a1", x"a2", x"a3", x"a3", x"a2", x"a2", x"a3", x"a3", x"a2", x"a2", x"a2", x"a0", x"a2", 
        x"a4", x"a4", x"a2", x"a2", x"a2", x"a2", x"a4", x"a3", x"a2", x"a3", x"a4", x"a5", x"a5", x"a3", x"a3", 
        x"a5", x"a4", x"a4", x"a5", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a5", x"a5", x"a4", x"a3", x"a3", 
        x"a3", x"a3", x"a4", x"a5", x"a6", x"a5", x"a4", x"a4", x"a5", x"a6", x"a6", x"a6", x"a4", x"a5", x"a6", 
        x"a4", x"a3", x"a5", x"a5", x"a4", x"a5", x"a8", x"89", x"56", x"79", x"a1", x"ac", x"a8", x"a1", x"94", 
        x"92", x"9b", x"b6", x"c7", x"d4", x"da", x"c8", x"a3", x"73", x"52", x"46", x"46", x"4c", x"57", x"64", 
        x"72", x"88", x"a6", x"c5", x"c5", x"96", x"86", x"8b", x"89", x"87", x"88", x"88", x"88", x"87", x"88", 
        x"86", x"7d", x"96", x"b1", x"bf", x"ca", x"d5", x"d7", x"e4", x"d4", x"d0", x"d4", x"d4", x"d5", x"d3", 
        x"d1", x"d2", x"d0", x"d1", x"d3", x"d3", x"d1", x"d1", x"d1", x"d0", x"d2", x"d3", x"d1", x"d0", x"d0", 
        x"d1", x"d2", x"d1", x"d1", x"d3", x"d4", x"d4", x"d2", x"d1", x"d1", x"d3", x"d3", x"d5", x"d4", x"d2", 
        x"d1", x"d3", x"d3", x"d2", x"d4", x"d4", x"d4", x"d6", x"d3", x"d2", x"db", x"d8", x"d6", x"d8", x"da", 
        x"d9", x"d6", x"da", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", x"ef", x"ef", x"f0", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ee", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ed", x"ef", x"ef", x"ee", x"ef", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", x"f0", x"e7", x"ef", 
        x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"f0", x"ee", x"ef", x"f2", x"f2", x"f1", x"f0", x"f1", x"f0", 
        x"ed", x"e8", x"e2", x"da", x"d2", x"ca", x"c0", x"b5", x"af", x"ac", x"aa", x"b3", x"c2", x"d6", x"e3", 
        x"ea", x"ed", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f2", x"f3", x"f4", x"f2", 
        x"f4", x"f4", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f4", x"f3", x"f3", x"f4", x"f5", x"f4", x"f5", x"f3", 
        x"f1", x"eb", x"e4", x"dc", x"d1", x"ca", x"c4", x"c5", x"d1", x"dc", x"e9", x"f0", x"f1", x"f0", x"ef", 
        x"f1", x"f2", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f4", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f1", x"f4", x"f6", x"f6", x"f6", x"f6", x"f6", x"f7", 
        x"e9", x"6c", x"5f", x"66", x"c6", x"da", x"d4", x"d5", x"d9", x"d3", x"a1", x"9e", x"a0", x"9e", x"9d", 
        x"9d", x"9b", x"9a", x"98", x"9a", x"98", x"95", x"93", x"93", x"93", x"92", x"91", x"92", x"91", x"92", 
        x"96", x"97", x"9b", x"9c", x"9c", x"73", x"53", x"44", x"81", x"86", x"89", x"88", x"85", x"86", x"86", 
        x"87", x"7f", x"78", x"76", x"79", x"79", x"78", x"78", x"78", x"78", x"79", x"7e", x"81", x"80", x"7f", 
        x"82", x"68", x"b7", x"e6", x"de", x"dd", x"e0", x"e0", x"dc", x"df", x"e0", x"df", x"de", x"de", x"dd", 
        x"df", x"df", x"df", x"de", x"de", x"dd", x"de", x"dd", x"de", x"df", x"e0", x"df", x"de", x"dc", x"dc", 
        x"dc", x"dc", x"dc", x"dc", x"dd", x"de", x"de", x"dd", x"dc", x"dc", x"db", x"db", x"dc", x"dc", x"dc", 
        x"dd", x"da", x"da", x"db", x"dc", x"dd", x"db", x"d9", x"d9", x"da", x"da", x"da", x"db", x"dc", x"dc", 
        x"db", x"dc", x"dc", x"dc", x"db", x"da", x"da", x"da", x"da", x"d9", x"d9", x"d9", x"da", x"da", x"d9", 
        x"dc", x"dc", x"d9", x"d9", x"db", x"dc", x"dc", x"d8", x"d3", x"cd", x"c5", x"bd", x"b7", x"b7", x"ba", 
        x"a6", x"a4", x"a4", x"a2", x"a1", x"a3", x"a1", x"a1", x"a3", x"a2", x"a1", x"a2", x"a0", x"a2", x"a2", 
        x"a0", x"a0", x"9f", x"9f", x"a0", x"a0", x"a1", x"a0", x"a0", x"a1", x"a1", x"a1", x"a1", x"a1", x"a1", 
        x"a1", x"a2", x"a3", x"a3", x"a2", x"a2", x"a1", x"a3", x"a0", x"a1", x"a2", x"9f", x"a1", x"a2", x"a2", 
        x"a1", x"a1", x"a2", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a1", x"a0", x"a3", 
        x"a4", x"a3", x"a3", x"a2", x"a2", x"a3", x"a5", x"a3", x"a1", x"a3", x"a4", x"a5", x"a5", x"a2", x"a3", 
        x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a5", x"a5", x"a5", x"a5", x"a4", x"a3", x"a2", 
        x"a3", x"a4", x"a6", x"a6", x"a6", x"a5", x"a4", x"a4", x"a5", x"a6", x"a7", x"a7", x"a4", x"a1", x"9f", 
        x"a1", x"a4", x"a5", x"a4", x"a3", x"a5", x"af", x"8c", x"53", x"77", x"9d", x"a0", x"93", x"91", x"a7", 
        x"c1", x"d1", x"d5", x"d2", x"be", x"8f", x"5e", x"43", x"42", x"47", x"52", x"5f", x"69", x"78", x"97", 
        x"bb", x"ca", x"d0", x"d6", x"c6", x"93", x"87", x"8a", x"88", x"89", x"8a", x"89", x"88", x"87", x"87", 
        x"83", x"7f", x"b1", x"d7", x"d9", x"d6", x"d8", x"d3", x"e1", x"d3", x"d0", x"d4", x"d4", x"d6", x"d4", 
        x"d2", x"d2", x"d1", x"d1", x"d2", x"d4", x"d3", x"d2", x"d1", x"d1", x"d1", x"d3", x"d2", x"d0", x"d0", 
        x"d2", x"d4", x"d3", x"d2", x"d3", x"d5", x"d4", x"d3", x"d2", x"d1", x"d3", x"d3", x"d6", x"d4", x"d2", 
        x"d2", x"d5", x"d3", x"d1", x"d3", x"d3", x"d4", x"d7", x"d4", x"d2", x"dc", x"d8", x"d6", x"d8", x"db", 
        x"d9", x"d7", x"d9", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f1", x"f2", x"ef", x"ef", x"f0", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ef", x"ee", x"ec", x"ee", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", x"e7", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", 
        x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", x"ef", x"f1", x"f0", x"f0", x"ef", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f2", x"f0", x"ea", x"e3", x"e1", x"da", x"cb", x"c0", x"b5", x"ab", x"a6", 
        x"a2", x"ac", x"bd", x"cd", x"db", x"e6", x"ec", x"f0", x"f2", x"f3", x"f2", x"f0", x"f1", x"f3", x"f3", 
        x"f1", x"ef", x"f0", x"f3", x"f3", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f0", x"ef", x"f0", 
        x"f4", x"f5", x"f4", x"f1", x"f0", x"f0", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ee", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f2", x"f3", x"f5", x"f2", 
        x"f3", x"f4", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f6", x"f5", x"f4", x"f6", x"f6", 
        x"f7", x"f6", x"f5", x"f3", x"ee", x"e8", x"e0", x"d7", x"d3", x"cc", x"cc", x"ce", x"cf", x"d6", x"e5", 
        x"ea", x"ee", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f3", x"f4", x"f4", x"f1", x"f0", 
        x"f0", x"f1", x"f3", x"f1", x"ef", x"ef", x"f3", x"f3", x"f4", x"f5", x"f5", x"f6", x"f6", x"f7", x"f7", 
        x"ec", x"74", x"5c", x"64", x"c1", x"da", x"d4", x"d5", x"d8", x"d4", x"a2", x"9e", x"a0", x"9f", x"9d", 
        x"9d", x"9c", x"9a", x"99", x"9b", x"99", x"96", x"94", x"93", x"93", x"93", x"92", x"91", x"91", x"92", 
        x"93", x"96", x"9b", x"9d", x"9f", x"76", x"54", x"47", x"82", x"86", x"8a", x"89", x"85", x"87", x"87", 
        x"88", x"7e", x"76", x"76", x"79", x"79", x"77", x"77", x"78", x"79", x"7a", x"7f", x"80", x"7f", x"7d", 
        x"81", x"67", x"b0", x"e5", x"de", x"de", x"df", x"df", x"dd", x"df", x"e0", x"df", x"df", x"de", x"de", 
        x"de", x"de", x"de", x"de", x"de", x"de", x"de", x"de", x"de", x"de", x"df", x"df", x"de", x"dd", x"dc", 
        x"dd", x"dc", x"dc", x"dc", x"dd", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"db", x"db", x"dc", x"dc", 
        x"db", x"da", x"db", x"dc", x"de", x"dd", x"da", x"d9", x"db", x"db", x"db", x"db", x"dc", x"dd", x"db", 
        x"da", x"db", x"dc", x"dd", x"dd", x"dd", x"dd", x"da", x"d9", x"d9", x"d9", x"d9", x"da", x"db", x"d9", 
        x"db", x"de", x"dd", x"d7", x"cd", x"c5", x"ba", x"b5", x"b5", x"b8", x"c0", x"c7", x"cd", x"d2", x"d4", 
        x"a4", x"a2", x"a3", x"a2", x"a1", x"a3", x"a2", x"a2", x"a4", x"a3", x"a1", x"a1", x"a0", x"a1", x"a2", 
        x"a0", x"a0", x"a0", x"a0", x"a0", x"a1", x"a1", x"a0", x"a1", x"a2", x"a2", x"a1", x"9f", x"9f", x"a1", 
        x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", x"a2", x"a3", x"a3", x"a4", x"a4", x"a1", x"a1", x"a1", x"a2", 
        x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a1", x"a2", x"a4", 
        x"a2", x"a1", x"a2", x"a3", x"a2", x"a3", x"a5", x"a4", x"a2", x"a3", x"a5", x"a4", x"a5", x"a3", x"a3", 
        x"a4", x"a4", x"a4", x"a4", x"a2", x"a2", x"a3", x"a4", x"a5", x"a5", x"a5", x"a5", x"a4", x"a3", x"a3", 
        x"a4", x"a5", x"a6", x"a6", x"a5", x"a4", x"a4", x"a4", x"a5", x"a5", x"a4", x"a5", x"a5", x"a3", x"a2", 
        x"a5", x"a7", x"a4", x"a2", x"a2", x"a3", x"ae", x"89", x"4a", x"63", x"82", x"9f", x"b3", x"c7", x"d6", 
        x"d8", x"ce", x"a5", x"78", x"50", x"3f", x"42", x"4d", x"5f", x"63", x"6e", x"8d", x"b2", x"c8", x"d0", 
        x"d1", x"d0", x"cf", x"d4", x"c9", x"98", x"88", x"8c", x"8c", x"8a", x"8a", x"8a", x"88", x"87", x"87", 
        x"80", x"7a", x"c0", x"e1", x"d3", x"d2", x"d7", x"d6", x"e6", x"d7", x"d1", x"d4", x"d3", x"d3", x"d1", 
        x"d2", x"d1", x"d1", x"d1", x"d3", x"d5", x"d5", x"d3", x"d2", x"d2", x"d2", x"d3", x"d2", x"d0", x"d1", 
        x"d3", x"d3", x"d3", x"d2", x"d2", x"d3", x"d4", x"d2", x"d3", x"d3", x"d3", x"d2", x"d4", x"d4", x"d3", 
        x"d2", x"d5", x"d4", x"d2", x"d4", x"d2", x"d4", x"d7", x"d4", x"d3", x"db", x"d8", x"d5", x"d8", x"db", 
        x"d9", x"d7", x"da", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"ef", x"ef", x"f0", 
        x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"ed", x"eb", x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f1", x"e6", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"ef", x"f1", x"f4", x"f4", x"f1", x"f0", x"f2", x"f0", x"ee", x"e9", x"e2", x"de", 
        x"d5", x"c6", x"b5", x"aa", x"a7", x"ac", x"b1", x"b9", x"c5", x"d5", x"e3", x"ea", x"ed", x"ef", x"ef", 
        x"f0", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", x"f1", x"f2", x"f2", x"f0", x"ee", 
        x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ee", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f2", x"f3", x"f4", x"f2", 
        x"f3", x"f4", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f3", x"f4", x"f7", x"f6", x"f4", x"f5", x"f8", 
        x"f9", x"f5", x"f4", x"f3", x"f2", x"f1", x"ed", x"ed", x"f1", x"ee", x"ea", x"e0", x"d5", x"cc", x"c2", 
        x"c3", x"c7", x"d2", x"df", x"ea", x"ef", x"f1", x"f3", x"f3", x"f1", x"f1", x"f1", x"ef", x"ef", x"f1", 
        x"f2", x"f0", x"ef", x"f1", x"f3", x"ef", x"f1", x"f4", x"f7", x"f5", x"f3", x"f3", x"f4", x"f6", x"f7", 
        x"ee", x"79", x"5a", x"62", x"bd", x"da", x"d4", x"d4", x"d8", x"d6", x"a5", x"9e", x"9f", x"9e", x"9d", 
        x"9d", x"9c", x"9a", x"99", x"99", x"99", x"97", x"96", x"95", x"95", x"95", x"94", x"8f", x"91", x"91", 
        x"8f", x"95", x"9a", x"9c", x"a0", x"79", x"54", x"47", x"80", x"87", x"89", x"89", x"85", x"86", x"88", 
        x"8a", x"7f", x"77", x"7a", x"79", x"79", x"78", x"77", x"78", x"7a", x"7a", x"7f", x"80", x"7f", x"7e", 
        x"80", x"68", x"a7", x"e3", x"df", x"de", x"de", x"de", x"df", x"e0", x"e0", x"e0", x"e0", x"e0", x"de", 
        x"dc", x"dd", x"de", x"de", x"de", x"de", x"de", x"de", x"de", x"dd", x"df", x"df", x"de", x"dd", x"dd", 
        x"de", x"de", x"de", x"dd", x"dd", x"dc", x"dc", x"dc", x"dd", x"dd", x"dc", x"db", x"db", x"db", x"dc", 
        x"dd", x"dd", x"dd", x"dd", x"dd", x"db", x"da", x"db", x"dd", x"db", x"db", x"da", x"d9", x"d9", x"da", 
        x"db", x"dc", x"dc", x"dd", x"dd", x"dd", x"dd", x"db", x"da", x"dc", x"dd", x"db", x"db", x"dc", x"d0", 
        x"c5", x"bb", x"b6", x"b4", x"b7", x"be", x"cd", x"d1", x"d4", x"d7", x"da", x"db", x"da", x"d8", x"d8", 
        x"a4", x"a3", x"a3", x"a2", x"a2", x"a2", x"a3", x"a2", x"a3", x"a3", x"a2", x"a1", x"a1", x"a2", x"a2", 
        x"a1", x"a1", x"a1", x"a1", x"a1", x"a1", x"a2", x"a1", x"a1", x"a1", x"a1", x"a0", x"9f", x"9f", x"a1", 
        x"a2", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a2", x"a2", x"a0", x"a2", 
        x"a4", x"a4", x"a3", x"a2", x"a3", x"a1", x"a1", x"a1", x"a1", x"a1", x"a1", x"a1", x"a0", x"a2", x"a4", 
        x"a3", x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", x"a3", x"a4", x"a4", x"a5", x"a4", x"a4", 
        x"a4", x"a4", x"a4", x"a4", x"a2", x"a3", x"a3", x"a4", x"a5", x"a4", x"a3", x"a4", x"a4", x"a4", x"a4", 
        x"a4", x"a5", x"a6", x"a5", x"a5", x"a4", x"a4", x"a4", x"a4", x"a5", x"a4", x"a5", x"a7", x"a7", x"a5", 
        x"a4", x"a6", x"a6", x"a4", x"a1", x"a3", x"a2", x"8a", x"78", x"a8", x"c9", x"d7", x"d8", x"cf", x"b3", 
        x"85", x"52", x"3b", x"3c", x"4c", x"60", x"66", x"6f", x"82", x"a9", x"c6", x"d6", x"d8", x"d2", x"d0", 
        x"d3", x"d2", x"d0", x"d3", x"ca", x"9a", x"88", x"8c", x"8e", x"8c", x"8b", x"8a", x"89", x"89", x"89", 
        x"82", x"7c", x"be", x"dd", x"d4", x"d7", x"d5", x"d7", x"e4", x"d6", x"cf", x"d3", x"d4", x"d4", x"d3", 
        x"d1", x"d0", x"d1", x"d3", x"d4", x"d5", x"d3", x"d2", x"d2", x"d3", x"d3", x"d3", x"d1", x"d0", x"d1", 
        x"d2", x"d2", x"d4", x"d3", x"d0", x"d1", x"d3", x"d2", x"d3", x"d5", x"d4", x"d3", x"d3", x"d4", x"d3", 
        x"d2", x"d5", x"d5", x"d3", x"d4", x"d2", x"d3", x"d6", x"d4", x"d4", x"db", x"d6", x"d5", x"d8", x"da", 
        x"d8", x"d7", x"d9", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"f1", x"e6", x"ee", 
        x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"ee", x"f0", x"ef", x"f0", x"f2", x"f1", x"ee", x"ed", x"ee", x"ef", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"ea", x"e1", x"d8", x"c5", x"b7", x"aa", x"a6", x"ac", x"b4", x"ba", x"cb", 
        x"d7", x"e1", x"e7", x"e9", x"ec", x"f0", x"f1", x"f1", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ee", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f2", 
        x"f2", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f6", x"f9", x"f7", x"f4", x"f5", x"f7", 
        x"f6", x"f4", x"f4", x"f2", x"f1", x"f1", x"ee", x"ef", x"f3", x"f2", x"f2", x"f3", x"f2", x"f3", x"ef", 
        x"e3", x"d0", x"bd", x"b7", x"b9", x"c1", x"cf", x"da", x"e5", x"ec", x"f0", x"f1", x"f0", x"f3", x"f3", 
        x"f1", x"f2", x"f3", x"f2", x"f1", x"f2", x"f4", x"f2", x"f4", x"f5", x"f5", x"f7", x"f5", x"f5", x"f6", 
        x"f0", x"81", x"57", x"5f", x"b7", x"da", x"d3", x"d3", x"d7", x"d9", x"a7", x"9d", x"9f", x"9e", x"9d", 
        x"9d", x"9d", x"9b", x"99", x"97", x"98", x"99", x"98", x"96", x"96", x"96", x"94", x"92", x"91", x"90", 
        x"90", x"94", x"98", x"9b", x"a1", x"7f", x"54", x"4a", x"7e", x"8a", x"8a", x"89", x"87", x"87", x"87", 
        x"8a", x"82", x"7a", x"7c", x"79", x"79", x"7a", x"77", x"78", x"79", x"78", x"7d", x"7f", x"7f", x"7f", 
        x"81", x"6c", x"a1", x"e3", x"e1", x"df", x"e0", x"df", x"df", x"e0", x"e0", x"e2", x"e2", x"e1", x"df", 
        x"dc", x"dc", x"de", x"de", x"de", x"de", x"de", x"de", x"dd", x"dc", x"de", x"df", x"de", x"de", x"de", 
        x"de", x"dd", x"dd", x"dd", x"dd", x"dd", x"dd", x"dd", x"de", x"de", x"dd", x"db", x"db", x"db", x"db", 
        x"da", x"da", x"da", x"db", x"db", x"db", x"db", x"db", x"d9", x"d8", x"d9", x"da", x"da", x"db", x"da", 
        x"db", x"dc", x"dd", x"dd", x"dc", x"da", x"d9", x"d8", x"cf", x"c9", x"c1", x"b6", x"b1", x"b3", x"b9", 
        x"c3", x"d0", x"d9", x"db", x"de", x"e1", x"dd", x"da", x"da", x"da", x"db", x"da", x"d9", x"d8", x"d8", 
        x"a6", x"a6", x"a4", x"a2", x"a2", x"a0", x"a1", x"a1", x"a1", x"a2", x"a2", x"a1", x"a2", x"a4", x"a3", 
        x"a2", x"a1", x"a1", x"a1", x"a2", x"a2", x"a2", x"a2", x"a1", x"a0", x"a0", x"a0", x"a0", x"a1", x"a2", 
        x"a2", x"a3", x"a4", x"a4", x"a3", x"a3", x"a2", x"a1", x"a2", x"a1", x"a1", x"a2", x"a2", x"a1", x"a2", 
        x"a4", x"a4", x"a4", x"a3", x"a3", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a3", x"a3", x"a2", x"a3", 
        x"a5", x"a4", x"a2", x"a1", x"a4", x"a4", x"a3", x"a3", x"a4", x"a4", x"a4", x"a4", x"a4", x"a5", x"a4", 
        x"a3", x"a3", x"a4", x"a4", x"a4", x"a4", x"a5", x"a5", x"a4", x"a3", x"a2", x"a4", x"a5", x"a5", x"a5", 
        x"a5", x"a5", x"a6", x"a5", x"a5", x"a4", x"a4", x"a4", x"a4", x"a5", x"a6", x"a5", x"a3", x"a5", x"a6", 
        x"a4", x"a1", x"a1", x"9f", x"9a", x"a4", x"b2", x"c9", x"cf", x"d8", x"ce", x"bb", x"9b", x"6d", x"49", 
        x"40", x"48", x"56", x"62", x"6c", x"79", x"96", x"b5", x"ca", x"d3", x"d3", x"d1", x"d1", x"d0", x"ce", 
        x"cf", x"d1", x"d2", x"d4", x"c9", x"99", x"88", x"8a", x"8b", x"8c", x"8b", x"8a", x"8a", x"8b", x"8b", 
        x"83", x"7c", x"bf", x"df", x"d4", x"d8", x"d4", x"d7", x"e4", x"d6", x"ce", x"d3", x"d5", x"d3", x"d4", 
        x"d1", x"cf", x"d0", x"d1", x"d2", x"d3", x"d2", x"d1", x"d2", x"d3", x"d3", x"d3", x"d1", x"d0", x"d0", 
        x"d1", x"d1", x"d3", x"d2", x"d0", x"d0", x"d2", x"d2", x"d4", x"d5", x"d4", x"d3", x"d2", x"d4", x"d4", 
        x"d2", x"d5", x"d5", x"d3", x"d4", x"d1", x"d3", x"d6", x"d5", x"d5", x"db", x"d5", x"d5", x"d8", x"da", 
        x"d8", x"d6", x"d8", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f1", x"e6", x"ee", 
        x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ed", x"ed", x"ee", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", 
        x"ef", x"f0", x"f1", x"ef", x"ef", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"ef", x"ee", x"ef", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"ec", x"e7", x"db", x"cc", x"be", x"b4", 
        x"b2", x"b2", x"b4", x"b9", x"c0", x"c7", x"d1", x"da", x"e2", x"e9", x"ec", x"f0", x"f4", x"f5", x"f3", 
        x"f2", x"f2", x"f1", x"f0", x"ee", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"ef", x"f3", 
        x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f3", x"f3", x"f4", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f7", x"f9", x"f7", x"f4", x"f5", x"f8", 
        x"f6", x"f3", x"f3", x"f1", x"f0", x"f1", x"f1", x"f1", x"f5", x"f2", x"f2", x"f2", x"f3", x"f5", x"f1", 
        x"f2", x"f2", x"ef", x"e8", x"de", x"d3", x"c5", x"bf", x"be", x"c2", x"c9", x"d1", x"db", x"e5", x"eb", 
        x"ef", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"ee", x"f2", x"f6", x"f8", x"f7", x"f6", x"f5", x"f6", 
        x"f0", x"87", x"55", x"5d", x"b0", x"da", x"d3", x"d3", x"d6", x"db", x"aa", x"9e", x"9e", x"9d", x"9d", 
        x"9d", x"9d", x"9b", x"9a", x"97", x"98", x"99", x"99", x"97", x"97", x"96", x"93", x"95", x"92", x"8f", 
        x"91", x"92", x"94", x"9a", x"a1", x"85", x"56", x"4c", x"7d", x"8f", x"8c", x"8d", x"8d", x"88", x"85", 
        x"87", x"82", x"7b", x"7a", x"79", x"7a", x"7a", x"78", x"78", x"79", x"7a", x"7f", x"81", x"80", x"80", 
        x"81", x"6d", x"9e", x"e5", x"e1", x"e0", x"e2", x"e2", x"df", x"df", x"e0", x"e1", x"e1", x"e0", x"df", 
        x"dd", x"dd", x"de", x"de", x"de", x"de", x"de", x"de", x"dd", x"dc", x"de", x"df", x"de", x"de", x"de", 
        x"de", x"dd", x"dd", x"dd", x"dd", x"de", x"de", x"de", x"de", x"de", x"dd", x"dc", x"db", x"db", x"db", 
        x"da", x"da", x"da", x"da", x"da", x"d8", x"d7", x"d9", x"da", x"db", x"dc", x"de", x"dd", x"db", x"d9", 
        x"d8", x"d6", x"d2", x"cc", x"c6", x"c1", x"bd", x"ba", x"bb", x"c5", x"cd", x"d0", x"d4", x"da", x"db", 
        x"dd", x"dd", x"db", x"da", x"dc", x"dc", x"db", x"d9", x"d9", x"da", x"db", x"da", x"d9", x"d9", x"d9", 
        x"a5", x"a6", x"a3", x"a2", x"a3", x"a1", x"a3", x"a2", x"a0", x"a3", x"a3", x"a1", x"a3", x"a3", x"a3", 
        x"a2", x"a2", x"a2", x"a2", x"a2", x"a3", x"a3", x"a2", x"a1", x"a0", x"a0", x"a1", x"a2", x"a2", x"a2", 
        x"a3", x"a3", x"a4", x"a4", x"a3", x"a3", x"a2", x"a0", x"a2", x"a1", x"a0", x"a3", x"a2", x"a2", x"a2", 
        x"a3", x"a3", x"a4", x"a4", x"a4", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a3", x"a4", 
        x"a6", x"a4", x"a2", x"a2", x"a4", x"a4", x"a2", x"a4", x"a6", x"a5", x"a4", x"a4", x"a4", x"a6", x"a4", 
        x"a2", x"a3", x"a5", x"a4", x"a4", x"a5", x"a6", x"a5", x"a4", x"a3", x"a1", x"a3", x"a4", x"a4", x"a5", 
        x"a5", x"a5", x"a4", x"a5", x"a5", x"a4", x"a4", x"a4", x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a1", 
        x"9a", x"9b", x"a2", x"ad", x"c2", x"d7", x"d8", x"d5", x"c4", x"a7", x"7f", x"59", x"43", x"3e", x"4c", 
        x"5e", x"6b", x"79", x"8f", x"aa", x"c5", x"d3", x"d6", x"d0", x"cf", x"d1", x"d2", x"d0", x"d1", x"d2", 
        x"d1", x"cf", x"d0", x"d5", x"cb", x"9a", x"89", x"8a", x"8a", x"8d", x"8a", x"89", x"8a", x"8c", x"8c", 
        x"85", x"7c", x"be", x"e1", x"d5", x"d7", x"d1", x"d5", x"e5", x"d8", x"ce", x"d2", x"d4", x"d2", x"d3", 
        x"d3", x"d1", x"cf", x"cf", x"d0", x"d1", x"d1", x"d2", x"d2", x"d4", x"d4", x"d3", x"d2", x"d1", x"d0", 
        x"cf", x"d1", x"d2", x"d1", x"d0", x"d0", x"d2", x"d2", x"d3", x"d4", x"d4", x"d4", x"d1", x"d3", x"d6", 
        x"d4", x"d6", x"d5", x"d4", x"d4", x"d2", x"d3", x"d5", x"d5", x"d7", x"dc", x"d5", x"d5", x"d8", x"da", 
        x"d8", x"d5", x"d9", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"f0", x"ef", x"ee", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", x"e6", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ee", x"ed", x"ee", 
        x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", 
        x"ee", x"ef", x"f1", x"f1", x"f1", x"f1", x"ef", x"ee", x"f0", x"ef", x"f0", x"ef", x"f0", x"f2", x"f0", 
        x"ee", x"ee", x"f0", x"f1", x"f0", x"ef", x"ee", x"f0", x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"ef", 
        x"e8", x"de", x"d4", x"c7", x"b9", x"ac", x"a9", x"ad", x"b5", x"be", x"c6", x"d0", x"d9", x"e2", x"eb", 
        x"ec", x"ee", x"f1", x"f1", x"f1", x"f0", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"ef", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f4", x"f3", x"f2", x"f4", 
        x"f3", x"f2", x"f4", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f3", x"f7", x"fa", x"f7", x"f4", x"f5", x"f7", 
        x"f4", x"f2", x"f4", x"f3", x"f1", x"f2", x"f1", x"ef", x"f3", x"f1", x"f1", x"f1", x"f1", x"f3", x"f2", 
        x"f3", x"f2", x"f1", x"f1", x"f3", x"f4", x"f3", x"ef", x"e6", x"d8", x"c9", x"bd", x"bc", x"c5", x"cc", 
        x"d4", x"db", x"e3", x"eb", x"ef", x"f2", x"f3", x"ef", x"f2", x"f5", x"f6", x"f5", x"f5", x"f5", x"f6", 
        x"f1", x"8f", x"55", x"5b", x"a9", x"d9", x"d3", x"d3", x"d6", x"dc", x"ad", x"9d", x"9e", x"9d", x"9d", 
        x"9d", x"9d", x"9c", x"9a", x"98", x"98", x"98", x"98", x"97", x"96", x"96", x"93", x"96", x"93", x"91", 
        x"92", x"91", x"92", x"98", x"a2", x"8a", x"56", x"4b", x"78", x"91", x"8c", x"8d", x"8e", x"87", x"85", 
        x"87", x"85", x"7b", x"79", x"79", x"79", x"78", x"77", x"78", x"7a", x"7b", x"80", x"82", x"81", x"81", 
        x"80", x"6f", x"9a", x"e5", x"e3", x"e0", x"e2", x"e1", x"df", x"df", x"e0", x"e0", x"e0", x"e0", x"e0", 
        x"df", x"de", x"de", x"de", x"de", x"de", x"de", x"de", x"dd", x"dd", x"df", x"df", x"de", x"dd", x"dd", 
        x"dd", x"dd", x"dd", x"dd", x"de", x"de", x"de", x"de", x"de", x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", 
        x"dc", x"db", x"da", x"db", x"dc", x"dd", x"dd", x"dd", x"dc", x"d9", x"d7", x"d4", x"cf", x"c9", x"c2", 
        x"bd", x"bb", x"ba", x"bd", x"c4", x"ca", x"d1", x"d7", x"d9", x"de", x"e0", x"dd", x"da", x"da", x"dc", 
        x"dc", x"da", x"d9", x"da", x"dc", x"da", x"dc", x"db", x"d8", x"d7", x"d8", x"d9", x"d9", x"d9", x"d9", 
        x"a5", x"a6", x"a3", x"a2", x"a3", x"a1", x"a3", x"a3", x"a0", x"a3", x"a3", x"a0", x"a1", x"a1", x"a2", 
        x"a3", x"a2", x"a2", x"a2", x"a2", x"a3", x"a3", x"a1", x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", x"a2", 
        x"a3", x"a3", x"a4", x"a4", x"a4", x"a4", x"a2", x"a0", x"a3", x"a3", x"a2", x"a5", x"a3", x"a4", x"a3", 
        x"a2", x"a3", x"a4", x"a4", x"a4", x"a4", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a4", x"a5", x"a5", 
        x"a3", x"a2", x"a2", x"a3", x"a4", x"a3", x"a2", x"a3", x"a6", x"a5", x"a4", x"a4", x"a4", x"a6", x"a4", 
        x"a2", x"a3", x"a5", x"a4", x"a3", x"a4", x"a6", x"a6", x"a5", x"a4", x"a2", x"a2", x"a3", x"a4", x"a4", 
        x"a5", x"a4", x"a4", x"a5", x"a6", x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a7", x"a5", x"a0", x"9f", 
        x"a9", x"bc", x"cc", x"da", x"df", x"d0", x"a9", x"7f", x"5c", x"45", x"3d", x"47", x"59", x"62", x"72", 
        x"8e", x"aa", x"c4", x"d3", x"d9", x"d3", x"cf", x"d0", x"ce", x"cf", x"cf", x"d1", x"d3", x"d2", x"d0", 
        x"d0", x"d3", x"d2", x"d2", x"c9", x"9a", x"8a", x"8c", x"8e", x"8e", x"8b", x"89", x"8a", x"8b", x"8b", 
        x"84", x"7f", x"bd", x"e3", x"d7", x"da", x"d3", x"d3", x"e4", x"d9", x"ce", x"d2", x"d4", x"d1", x"d3", 
        x"d4", x"d4", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d2", x"d4", x"d4", x"d3", x"d2", x"d2", x"d0", 
        x"cf", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d2", x"d2", x"d4", x"d4", x"d6", x"d1", x"d2", x"d6", 
        x"d4", x"d4", x"d4", x"d3", x"d4", x"d1", x"d3", x"d4", x"d5", x"d7", x"dc", x"d4", x"d5", x"d8", x"da", 
        x"d7", x"d5", x"d8", x"ed", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"f0", x"f0", x"ef", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f2", x"e7", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"f1", x"f2", x"f1", x"ef", x"ef", 
        x"ee", x"ef", x"f0", x"ef", x"f0", x"f1", x"f0", x"ee", x"ef", x"ef", x"f1", x"ef", x"f0", x"f2", x"f0", 
        x"f1", x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"ef", 
        x"ef", x"f1", x"f3", x"f3", x"f2", x"f2", x"e8", x"dc", x"ce", x"bf", x"b8", x"b3", x"b0", x"b2", x"b5", 
        x"b6", x"bc", x"c7", x"d6", x"e3", x"eb", x"f3", x"f6", x"f7", x"f7", x"f4", x"f2", x"f1", x"f1", x"f0", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"ef", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f4", x"f3", x"f2", x"f4", 
        x"f2", x"f2", x"f4", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f3", x"f7", x"fa", x"f6", x"f4", x"f6", x"f9", 
        x"f6", x"f2", x"f5", x"f4", x"ef", x"f0", x"f0", x"ef", x"f3", x"f2", x"f2", x"f3", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f4", x"f2", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"ee", x"e8", x"dc", x"d2", 
        x"c5", x"bf", x"c1", x"c9", x"cf", x"d6", x"e0", x"ea", x"f4", x"f7", x"f7", x"f8", x"f6", x"f5", x"f7", 
        x"f2", x"95", x"57", x"5a", x"a2", x"d9", x"d3", x"d2", x"d5", x"de", x"af", x"9c", x"9e", x"9d", x"9d", 
        x"9d", x"9d", x"9c", x"9b", x"99", x"98", x"97", x"96", x"97", x"96", x"94", x"94", x"94", x"95", x"94", 
        x"90", x"91", x"91", x"95", x"a2", x"8f", x"55", x"4a", x"73", x"90", x"8c", x"8d", x"8e", x"88", x"87", 
        x"89", x"85", x"79", x"78", x"7a", x"78", x"75", x"76", x"7a", x"7a", x"78", x"7d", x"81", x"82", x"84", 
        x"84", x"74", x"94", x"e5", x"e4", x"df", x"de", x"de", x"e1", x"df", x"df", x"df", x"df", x"e0", x"e1", 
        x"e1", x"df", x"de", x"de", x"de", x"de", x"de", x"de", x"de", x"df", x"e0", x"e0", x"de", x"dd", x"dc", 
        x"dd", x"de", x"de", x"de", x"de", x"dd", x"dd", x"dd", x"de", x"dd", x"dd", x"dd", x"dc", x"dc", x"de", 
        x"de", x"dd", x"df", x"e0", x"de", x"d8", x"d0", x"c8", x"c1", x"bc", x"ba", x"bc", x"bf", x"c1", x"c3", 
        x"c9", x"d1", x"da", x"df", x"e0", x"df", x"dc", x"da", x"d9", x"da", x"da", x"da", x"d9", x"db", x"db", 
        x"db", x"da", x"da", x"d9", x"da", x"dc", x"db", x"da", x"d9", x"d9", x"db", x"db", x"db", x"d8", x"d7", 
        x"a6", x"a6", x"a4", x"a3", x"a3", x"a1", x"a1", x"a2", x"a2", x"a3", x"a4", x"a1", x"a2", x"a1", x"a2", 
        x"a3", x"a4", x"a3", x"a2", x"a2", x"a1", x"a2", x"a1", x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", x"a3", 
        x"a3", x"a2", x"a2", x"a3", x"a3", x"a3", x"a2", x"a2", x"a5", x"a5", x"a3", x"a3", x"a2", x"a4", x"a3", 
        x"a2", x"a3", x"a3", x"a4", x"a4", x"a2", x"a2", x"a4", x"a4", x"a4", x"a3", x"a3", x"a3", x"a5", x"a5", 
        x"a3", x"a3", x"a4", x"a5", x"a5", x"a4", x"a3", x"a4", x"a5", x"a5", x"a5", x"a4", x"a4", x"a6", x"a4", 
        x"a3", x"a4", x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a5", x"a5", x"a4", x"a4", x"a5", x"a6", 
        x"a6", x"a5", x"a4", x"a5", x"a6", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a4", x"9f", x"b4", x"c0", 
        x"cd", x"db", x"d3", x"b8", x"85", x"5e", x"45", x"38", x"41", x"53", x"60", x"70", x"88", x"a2", x"bd", 
        x"cf", x"d6", x"d3", x"d2", x"d0", x"d0", x"d1", x"d1", x"d1", x"d1", x"d3", x"d3", x"d2", x"d1", x"d1", 
        x"d2", x"d2", x"d1", x"d5", x"ca", x"9a", x"89", x"8c", x"90", x"8e", x"8b", x"89", x"8a", x"8b", x"8b", 
        x"85", x"7a", x"bb", x"e1", x"d4", x"d9", x"d7", x"d5", x"e4", x"d6", x"ce", x"d2", x"d2", x"d2", x"d2", 
        x"d2", x"d2", x"d1", x"d3", x"d4", x"d3", x"d3", x"d2", x"d2", x"d3", x"d4", x"d3", x"d1", x"d0", x"cf", 
        x"d0", x"d1", x"d1", x"d2", x"d4", x"d5", x"d5", x"d2", x"d3", x"d3", x"d2", x"d3", x"d2", x"d3", x"d3", 
        x"d1", x"d4", x"d4", x"d3", x"d5", x"d3", x"d2", x"d4", x"d6", x"d7", x"dd", x"d5", x"d5", x"d7", x"db", 
        x"d8", x"d5", x"d7", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ee", x"ec", x"ee", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"f2", x"e8", x"ee", 
        x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ee", x"ef", x"f0", x"ef", 
        x"ef", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f0", x"ef", x"f0", 
        x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"eb", x"e2", x"da", x"d1", 
        x"c8", x"bf", x"ba", x"b7", x"b5", x"b6", x"ba", x"c3", x"ce", x"da", x"e6", x"ed", x"f1", x"f2", x"f3", 
        x"f3", x"f2", x"f1", x"f2", x"f3", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f2", x"f1", x"ee", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f4", 
        x"f3", x"f2", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f3", x"f3", x"f1", x"f2", x"f4", x"f3", x"f4", x"f5", x"f8", x"fa", x"f6", x"f3", x"f6", x"f6", 
        x"f3", x"f2", x"f2", x"f2", x"f0", x"f1", x"f0", x"f0", x"f3", x"f0", x"f2", x"f3", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"ef", x"ef", x"f1", x"f1", x"f3", x"f3", 
        x"ef", x"e8", x"e1", x"d8", x"ce", x"ca", x"c9", x"c8", x"cd", x"da", x"e7", x"ef", x"f4", x"f5", x"f6", 
        x"f2", x"9b", x"54", x"5b", x"9d", x"d8", x"d3", x"d3", x"d7", x"dd", x"b2", x"9e", x"9e", x"9d", x"9b", 
        x"9b", x"9b", x"9a", x"99", x"98", x"99", x"99", x"99", x"96", x"95", x"95", x"95", x"93", x"93", x"92", 
        x"91", x"91", x"90", x"92", x"9f", x"91", x"53", x"4e", x"73", x"91", x"8d", x"8e", x"8b", x"8b", x"8a", 
        x"89", x"84", x"79", x"79", x"78", x"77", x"77", x"77", x"79", x"7a", x"78", x"7f", x"81", x"84", x"85", 
        x"82", x"76", x"8f", x"e3", x"e3", x"de", x"e0", x"e0", x"e1", x"e0", x"e0", x"e0", x"e0", x"e0", x"e1", 
        x"e1", x"e1", x"df", x"de", x"de", x"df", x"e0", x"df", x"de", x"de", x"e1", x"e1", x"df", x"dc", x"dc", 
        x"dd", x"df", x"df", x"de", x"de", x"dd", x"db", x"db", x"dd", x"de", x"df", x"df", x"de", x"de", x"de", 
        x"d6", x"ce", x"c6", x"c0", x"bd", x"bf", x"c3", x"c6", x"c7", x"c8", x"cc", x"d2", x"da", x"e0", x"e2", 
        x"df", x"de", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"dc", x"dd", x"dc", x"dc", x"da", 
        x"d9", x"da", x"d9", x"d8", x"d9", x"db", x"db", x"d9", x"d8", x"d9", x"d9", x"d9", x"db", x"da", x"d9", 
        x"a6", x"a6", x"a5", x"a4", x"a3", x"a2", x"a1", x"a2", x"a3", x"a3", x"a3", x"a2", x"a2", x"a2", x"a1", 
        x"a3", x"a4", x"a3", x"a2", x"a2", x"a2", x"a2", x"a3", x"a2", x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", 
        x"a3", x"a2", x"a2", x"a2", x"a3", x"a4", x"a4", x"a4", x"a3", x"a2", x"a2", x"a2", x"a2", x"a3", x"a4", 
        x"a3", x"a3", x"a3", x"a3", x"a3", x"a2", x"a3", x"a5", x"a5", x"a5", x"a4", x"a3", x"a3", x"a3", x"a3", 
        x"a3", x"a4", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a4", x"a4", x"a4", x"a4", x"a4", x"a5", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a4", x"a5", x"a6", x"a6", 
        x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a8", x"a5", x"a2", x"cc", x"dc", 
        x"ce", x"a6", x"74", x"4b", x"33", x"36", x"48", x"51", x"5f", x"72", x"96", x"ae", x"c4", x"d5", x"d7", 
        x"d5", x"cf", x"d0", x"d1", x"d1", x"d0", x"d1", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", 
        x"d2", x"d2", x"d2", x"d7", x"ca", x"99", x"89", x"8b", x"8e", x"8e", x"8d", x"8b", x"88", x"89", x"87", 
        x"84", x"7a", x"bb", x"e3", x"d5", x"d6", x"d3", x"d5", x"e3", x"d3", x"cd", x"d2", x"d1", x"d4", x"d3", 
        x"d1", x"d2", x"d1", x"d5", x"d5", x"d3", x"d3", x"d0", x"d0", x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", 
        x"d3", x"d2", x"d2", x"d2", x"d3", x"d4", x"d4", x"d2", x"d3", x"d3", x"d2", x"d2", x"d3", x"d3", x"d2", 
        x"d0", x"d3", x"d3", x"d2", x"d5", x"d4", x"d3", x"d4", x"d6", x"d7", x"dd", x"d5", x"d5", x"d7", x"dc", 
        x"d9", x"d5", x"d8", x"ef", x"ef", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"ef", x"ee", x"ec", x"ee", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", 
        x"f0", x"f1", x"ef", x"ee", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ee", x"f2", x"e9", x"ec", 
        x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ed", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"f0", x"f2", x"f4", x"f4", x"f4", x"f4", x"f3", 
        x"f2", x"ef", x"e9", x"df", x"d4", x"cc", x"c2", x"bb", x"b4", x"af", x"b2", x"b6", x"bb", x"c7", x"d6", 
        x"e5", x"ee", x"f2", x"f4", x"f5", x"f2", x"f2", x"f3", x"f1", x"f0", x"f2", x"f3", x"f2", x"f3", x"f4", 
        x"f4", x"f4", x"f3", x"f1", x"f0", x"f1", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f4", x"f4", x"f5", x"f4", x"f4", x"f2", x"f1", x"f3", x"f1", x"ed", x"f3", 
        x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", 
        x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", 
        x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f2", x"f3", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f3", x"f4", x"f2", x"f3", x"f5", x"f3", x"f5", x"f7", x"f9", x"fa", x"f6", x"f3", x"f5", x"f4", 
        x"f3", x"f4", x"f3", x"f1", x"f1", x"f2", x"f0", x"f0", x"f2", x"ef", x"f1", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", 
        x"f1", x"f1", x"f4", x"f3", x"ed", x"ea", x"e4", x"d6", x"ce", x"ce", x"cc", x"cc", x"d0", x"d8", x"e0", 
        x"e9", x"a1", x"57", x"5d", x"96", x"d9", x"d4", x"d2", x"d5", x"da", x"b5", x"a0", x"9f", x"9d", x"9b", 
        x"9a", x"9b", x"9b", x"9b", x"99", x"98", x"97", x"96", x"95", x"94", x"94", x"96", x"94", x"93", x"92", 
        x"93", x"93", x"90", x"91", x"9d", x"95", x"55", x"54", x"73", x"92", x"8e", x"90", x"8a", x"8d", x"8c", 
        x"89", x"86", x"7c", x"7a", x"77", x"78", x"7a", x"78", x"78", x"79", x"79", x"80", x"82", x"84", x"84", 
        x"82", x"79", x"8a", x"e0", x"e2", x"df", x"e1", x"e2", x"e1", x"e0", x"df", x"e1", x"e2", x"e2", x"e1", 
        x"df", x"e0", x"e1", x"e0", x"e0", x"e1", x"e1", x"e0", x"de", x"dc", x"de", x"df", x"dd", x"dc", x"de", 
        x"e0", x"df", x"df", x"dd", x"dd", x"de", x"df", x"e0", x"e0", x"dd", x"d5", x"cb", x"c2", x"bd", x"bc", 
        x"bd", x"c0", x"c3", x"c6", x"c9", x"cf", x"d6", x"dc", x"de", x"df", x"de", x"dc", x"dc", x"dc", x"dc", 
        x"dc", x"dc", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"db", x"dc", x"dd", x"dc", x"da", x"da", 
        x"d9", x"d9", x"d9", x"d9", x"d9", x"da", x"db", x"d9", x"d9", x"db", x"db", x"d9", x"da", x"d9", x"d9", 
        x"a6", x"a5", x"a4", x"a3", x"a3", x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", x"a2", x"a2", x"a1", x"a3", 
        x"a4", x"a3", x"a2", x"a2", x"a3", x"a4", x"a4", x"a4", x"a3", x"a3", x"a2", x"a2", x"a3", x"a3", x"a4", 
        x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", x"a5", x"a4", x"a2", x"a1", x"a1", x"a3", x"a4", x"a4", x"a4", 
        x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a5", x"a5", x"a6", x"a5", x"a5", x"a5", x"a5", x"a4", 
        x"a4", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a4", x"a4", x"a4", x"a3", x"a4", x"a5", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a4", x"a4", x"a5", x"a5", 
        x"a6", x"a7", x"a8", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"ab", x"af", x"8b", 
        x"59", x"36", x"32", x"3f", x"52", x"5f", x"6d", x"89", x"ac", x"c2", x"d0", x"d7", x"d6", x"d3", x"cf", 
        x"d2", x"d2", x"d3", x"d2", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", 
        x"d2", x"d2", x"d1", x"d6", x"ca", x"9a", x"8a", x"8b", x"8c", x"8c", x"8e", x"8b", x"87", x"8a", x"8c", 
        x"86", x"7e", x"b9", x"e3", x"d8", x"d8", x"d6", x"d7", x"e5", x"d5", x"ce", x"d2", x"d2", x"d3", x"d3", 
        x"d3", x"d3", x"d2", x"d6", x"d5", x"d2", x"d0", x"ce", x"ce", x"d0", x"d2", x"d4", x"d4", x"d5", x"d3", 
        x"d0", x"d1", x"d1", x"d1", x"d2", x"d3", x"d3", x"d2", x"d3", x"d4", x"d4", x"d4", x"d3", x"d3", x"d4", 
        x"d2", x"d3", x"d2", x"d1", x"d3", x"d3", x"d4", x"d5", x"d6", x"d6", x"dc", x"d5", x"d6", x"d8", x"db", 
        x"d9", x"d5", x"d8", x"ef", x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ee", x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"f0", x"f1", x"f0", x"ef", 
        x"f0", x"f0", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f2", x"e9", x"ec", 
        x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ed", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"ef", x"f0", x"f1", x"f2", x"f2", x"f0", x"ee", x"ed", x"e8", x"e1", x"d7", x"ce", x"c6", x"b7", x"b1", 
        x"a9", x"a2", x"a8", x"b6", x"c7", x"d9", x"e4", x"ed", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", x"f2", x"f3", x"f1", x"ed", x"f3", 
        x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f2", x"f0", x"f0", x"f1", 
        x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f2", x"f3", x"f3", x"f2", x"f3", x"f4", x"f4", x"f6", x"f7", x"f9", x"f9", x"f5", x"f3", x"f5", x"f3", 
        x"f3", x"f3", x"f3", x"f1", x"f1", x"f2", x"f0", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", 
        x"f0", x"ee", x"f0", x"f1", x"ef", x"ef", x"f4", x"f5", x"f3", x"f0", x"e8", x"e2", x"d9", x"cd", x"c5", 
        x"c1", x"82", x"48", x"5b", x"92", x"d8", x"d8", x"d5", x"d6", x"db", x"b7", x"9e", x"a1", x"9f", x"9c", 
        x"9d", x"9e", x"9c", x"9a", x"98", x"98", x"99", x"98", x"96", x"94", x"94", x"94", x"94", x"93", x"93", 
        x"93", x"92", x"90", x"90", x"98", x"95", x"56", x"55", x"6e", x"92", x"8e", x"93", x"8d", x"8d", x"8c", 
        x"8a", x"88", x"7c", x"78", x"78", x"7a", x"7a", x"79", x"78", x"78", x"78", x"7f", x"80", x"82", x"83", 
        x"83", x"7e", x"84", x"d9", x"e2", x"e0", x"e2", x"e1", x"e1", x"e0", x"e0", x"e1", x"e1", x"e2", x"e2", 
        x"e2", x"e0", x"de", x"df", x"e0", x"df", x"de", x"de", x"de", x"df", x"df", x"df", x"de", x"dd", x"dd", 
        x"de", x"e2", x"e2", x"e2", x"dc", x"d3", x"c8", x"c0", x"bc", x"bd", x"bf", x"c3", x"c8", x"d0", x"d6", 
        x"da", x"db", x"dc", x"dc", x"dd", x"df", x"e1", x"dd", x"da", x"db", x"dc", x"db", x"dc", x"dd", x"de", 
        x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", x"dc", x"dc", x"db", x"db", x"db", x"dc", x"dc", x"dc", x"dc", 
        x"db", x"da", x"d9", x"d9", x"d9", x"da", x"da", x"d8", x"d8", x"da", x"db", x"da", x"d9", x"db", x"da", 
        x"a5", x"a4", x"a3", x"a3", x"a2", x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", x"a2", x"a2", x"a2", x"a3", 
        x"a4", x"a2", x"a2", x"a3", x"a5", x"a5", x"a4", x"a3", x"a4", x"a4", x"a4", x"a3", x"a3", x"a3", x"a4", 
        x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", 
        x"a4", x"a5", x"a5", x"a4", x"a4", x"a5", x"a4", x"a3", x"a3", x"a4", x"a5", x"a6", x"a6", x"a6", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a5", x"a6", x"a5", x"a5", x"a5", x"a4", x"a4", x"a4", x"a4", x"a5", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a5", x"a5", x"a5", x"a5", 
        x"a5", x"a6", x"a8", x"a7", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", x"a7", x"a2", x"90", 
        x"7a", x"5e", x"59", x"66", x"86", x"a6", x"c0", x"d5", x"d8", x"d3", x"d2", x"d0", x"d0", x"d2", x"d0", 
        x"d2", x"d5", x"d6", x"d4", x"d2", x"d2", x"d1", x"d0", x"d2", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", 
        x"d2", x"d2", x"d1", x"d5", x"ca", x"9b", x"8a", x"8a", x"8b", x"8a", x"8b", x"8b", x"88", x"8a", x"88", 
        x"80", x"7d", x"ba", x"e4", x"d5", x"d7", x"d9", x"d5", x"e5", x"d6", x"d0", x"d2", x"d2", x"d1", x"d1", 
        x"d3", x"d1", x"d0", x"d3", x"d4", x"d3", x"d3", x"d1", x"d0", x"d1", x"d2", x"d3", x"d3", x"d3", x"d2", 
        x"d1", x"d3", x"d4", x"d4", x"d3", x"d2", x"d3", x"d3", x"d2", x"d4", x"d6", x"d7", x"d4", x"d2", x"d5", 
        x"d4", x"d2", x"d1", x"d0", x"d2", x"d2", x"d2", x"d2", x"d4", x"d6", x"de", x"d7", x"d8", x"d8", x"db", 
        x"d8", x"d6", x"d9", x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"ef", x"ee", x"ed", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"f0", x"f2", x"f0", x"ef", 
        x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"f2", x"e9", x"ec", 
        x"f0", x"ef", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f4", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"f2", x"f3", x"f3", x"f1", x"f1", x"f4", x"f4", x"f4", x"f4", x"f3", x"f1", x"f0", x"ea", x"e6", 
        x"e0", x"d5", x"c8", x"ba", x"b0", x"a7", x"a8", x"ac", x"b2", x"be", x"cf", x"df", x"e7", x"eb", x"f0", 
        x"f2", x"f2", x"f2", x"f1", x"f0", x"f2", x"f4", x"f4", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f0", x"ed", x"f3", 
        x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f5", x"f5", x"f7", x"f8", x"f8", x"f7", x"f5", x"f3", x"f4", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f0", x"ef", x"f2", x"f2", x"f1", x"f0", x"f1", x"f3", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", 
        x"f3", x"f2", x"f1", x"f1", x"f0", x"f1", x"f4", x"f2", x"f1", x"f3", x"f3", x"f5", x"f5", x"f1", x"ed", 
        x"e7", x"9e", x"4e", x"54", x"73", x"a9", x"b3", x"bf", x"cb", x"d7", x"bb", x"a0", x"a0", x"a0", x"9f", 
        x"9b", x"98", x"98", x"9a", x"9a", x"9a", x"99", x"97", x"95", x"96", x"96", x"94", x"94", x"94", x"94", 
        x"92", x"91", x"90", x"90", x"93", x"95", x"59", x"57", x"6c", x"99", x"90", x"93", x"8e", x"8e", x"8b", 
        x"8b", x"89", x"7d", x"78", x"78", x"79", x"79", x"78", x"78", x"78", x"79", x"7f", x"81", x"81", x"81", 
        x"82", x"80", x"7e", x"d3", x"e3", x"e1", x"e2", x"e2", x"e2", x"e0", x"df", x"e0", x"e0", x"e0", x"e0", 
        x"e0", x"df", x"dd", x"dd", x"dd", x"de", x"df", x"df", x"df", x"e0", x"e1", x"e2", x"e1", x"dc", x"d6", 
        x"cf", x"ca", x"c4", x"bd", x"bb", x"c0", x"c9", x"d1", x"d5", x"d8", x"db", x"dc", x"dc", x"dd", x"de", 
        x"dc", x"db", x"dc", x"dd", x"de", x"de", x"dd", x"dc", x"dd", x"de", x"de", x"dd", x"de", x"de", x"de", 
        x"de", x"de", x"dd", x"dd", x"dd", x"dd", x"dc", x"dc", x"db", x"db", x"db", x"db", x"dc", x"dc", x"dc", 
        x"dc", x"dc", x"dc", x"db", x"da", x"d9", x"d9", x"d8", x"d9", x"da", x"db", x"da", x"db", x"dc", x"dc", 
        x"a5", x"a4", x"a3", x"a2", x"a2", x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", 
        x"a3", x"a3", x"a3", x"a5", x"a6", x"a4", x"a3", x"a1", x"a3", x"a5", x"a5", x"a5", x"a3", x"a3", x"a4", 
        x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", x"a2", x"a3", x"a5", x"a5", x"a5", x"a3", x"a3", x"a3", x"a4", 
        x"a4", x"a5", x"a5", x"a4", x"a4", x"a5", x"a4", x"a2", x"a2", x"a3", x"a5", x"a5", x"a6", x"a6", x"a6", 
        x"a6", x"a6", x"a5", x"a5", x"a5", x"a6", x"a6", x"a5", x"a5", x"a5", x"a5", x"a4", x"a5", x"a5", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a5", 
        x"a5", x"a5", x"a6", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a9", x"a6", x"a4", x"a5", x"aa", 
        x"a5", x"8b", x"90", x"b7", x"d0", x"d6", x"d3", x"d8", x"d5", x"d0", x"d2", x"d2", x"d3", x"d6", x"d2", 
        x"d2", x"d2", x"d5", x"d4", x"d2", x"d2", x"d1", x"d0", x"d2", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", 
        x"d3", x"d2", x"d1", x"d5", x"ca", x"9b", x"8a", x"8a", x"8d", x"8d", x"8a", x"8b", x"88", x"8a", x"8b", 
        x"85", x"7d", x"bc", x"e6", x"d4", x"d5", x"d7", x"d3", x"e4", x"d7", x"d0", x"d1", x"d1", x"cf", x"d1", 
        x"d2", x"cf", x"cf", x"d2", x"d4", x"d4", x"d4", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"cf", 
        x"ce", x"d2", x"d5", x"d5", x"d3", x"d1", x"d1", x"d2", x"d2", x"d3", x"d6", x"d7", x"d4", x"d2", x"d5", 
        x"d5", x"d2", x"d1", x"d1", x"d2", x"d3", x"d0", x"d1", x"d5", x"d7", x"df", x"d7", x"d7", x"d8", x"da", 
        x"d7", x"d7", x"da", x"f0", x"f2", x"f0", x"f1", x"f0", x"ef", x"ee", x"ee", x"ec", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"f2", x"e9", x"ec", 
        x"f0", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f4", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f1", x"f0", 
        x"ef", x"f0", x"f1", x"f2", x"f0", x"f0", x"ef", x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f5", x"f3", x"ef", x"eb", x"e5", x"df", x"d3", x"c1", x"b2", x"a7", x"a3", x"a8", x"b0", x"be", 
        x"cd", x"d9", x"e4", x"e9", x"eb", x"ee", x"f0", x"f1", x"f1", x"f0", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f0", x"ec", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f4", x"f3", x"f3", x"f4", x"f4", x"f4", x"f5", x"f7", x"f9", x"f8", x"f6", x"f4", x"f4", x"f3", x"f2", 
        x"f2", x"f3", x"f2", x"f0", x"f0", x"f1", x"f0", x"ef", x"f1", x"f3", x"f1", x"ef", x"f1", x"f3", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f4", x"f4", x"f2", x"f0", x"f0", x"f6", x"f8", x"f4", x"f2", x"f6", x"f5", x"f4", x"f5", x"f5", x"f6", 
        x"f6", x"b3", x"56", x"5b", x"83", x"c3", x"b4", x"a3", x"9e", x"a7", x"9b", x"8d", x"99", x"9d", x"a0", 
        x"a2", x"a1", x"9e", x"9b", x"9c", x"9a", x"99", x"98", x"96", x"93", x"91", x"93", x"94", x"94", x"93", 
        x"92", x"91", x"91", x"91", x"93", x"95", x"5a", x"57", x"67", x"9b", x"90", x"91", x"8e", x"8e", x"8b", 
        x"8b", x"8a", x"7d", x"78", x"79", x"79", x"77", x"77", x"78", x"79", x"79", x"7f", x"83", x"83", x"82", 
        x"81", x"80", x"7c", x"d0", x"e5", x"e2", x"e1", x"e0", x"e0", x"e1", x"e1", x"e0", x"df", x"df", x"df", 
        x"e0", x"e0", x"de", x"dc", x"dc", x"df", x"e0", x"df", x"dc", x"d8", x"cf", x"c6", x"c1", x"be", x"bd", 
        x"bd", x"c4", x"cb", x"d4", x"dc", x"df", x"df", x"de", x"de", x"e0", x"e0", x"df", x"de", x"de", x"de", 
        x"db", x"da", x"dc", x"dd", x"de", x"de", x"dd", x"dd", x"de", x"de", x"de", x"dc", x"dc", x"dc", x"dd", 
        x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", x"db", x"dc", x"dc", x"db", x"db", x"db", x"dc", x"dc", x"dc", 
        x"dd", x"de", x"dd", x"dc", x"da", x"d8", x"d5", x"d9", x"dd", x"de", x"de", x"dc", x"db", x"dc", x"dc", 
        x"a5", x"a3", x"a2", x"a2", x"a2", x"a2", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", 
        x"a3", x"a4", x"a5", x"a5", x"a4", x"a3", x"a2", x"a2", x"a3", x"a5", x"a5", x"a5", x"a4", x"a4", x"a4", 
        x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a3", x"a4", x"a4", x"a4", x"a4", x"a5", x"a4", x"a4", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a5", x"a4", x"a3", x"a2", x"a2", x"a3", x"a4", x"a5", x"a5", x"a6", x"a6", 
        x"a6", x"a6", x"a6", x"a5", x"a5", x"a6", x"a6", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", 
        x"a5", x"a5", x"a5", x"a6", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a9", x"a8", x"aa", x"a8", x"a5", 
        x"a3", x"bf", x"d6", x"d7", x"d0", x"cf", x"d1", x"d9", x"d3", x"d0", x"d2", x"d4", x"d1", x"d3", x"d6", 
        x"d7", x"d4", x"d4", x"d4", x"d3", x"d2", x"d2", x"d2", x"d2", x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", 
        x"d4", x"d2", x"d0", x"d5", x"c9", x"99", x"89", x"8a", x"8b", x"86", x"84", x"88", x"87", x"8a", x"8e", 
        x"89", x"81", x"ba", x"e0", x"d5", x"d8", x"d6", x"d2", x"e3", x"d7", x"d0", x"d0", x"d1", x"ce", x"d0", 
        x"d1", x"cf", x"d3", x"d4", x"d4", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"cd", 
        x"c8", x"ce", x"d2", x"d2", x"d1", x"d0", x"d1", x"d2", x"d1", x"d1", x"d4", x"d6", x"d4", x"d2", x"d4", 
        x"d5", x"d2", x"d2", x"d2", x"d1", x"d3", x"d3", x"d3", x"d7", x"d8", x"de", x"d5", x"d5", x"d8", x"da", 
        x"d7", x"d7", x"d9", x"ee", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", 
        x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"f2", x"e9", x"ec", 
        x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ef", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f0", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f3", x"f4", x"f2", x"ec", x"e5", x"de", x"d7", x"cb", x"b8", 
        x"aa", x"a6", x"aa", x"b1", x"ba", x"c4", x"cf", x"da", x"e3", x"e9", x"ec", x"ee", x"f0", x"f1", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f3", x"f3", x"f3", x"f0", x"ec", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f3", x"f1", 
        x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f4", x"f3", x"f3", x"f5", x"f4", x"f4", x"f5", x"f8", x"f9", x"f8", x"f4", x"f4", x"f4", x"f2", x"f1", 
        x"f2", x"f3", x"f2", x"f0", x"f0", x"f1", x"f1", x"ee", x"f0", x"f4", x"f1", x"ef", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"ef", x"ee", x"f1", x"f5", x"f4", x"ef", x"f0", x"f6", x"f7", x"f5", x"f7", x"f7", x"f5", 
        x"f7", x"bd", x"55", x"57", x"83", x"d2", x"d6", x"d7", x"d2", x"c8", x"a5", x"7a", x"70", x"74", x"7e", 
        x"88", x"91", x"95", x"97", x"9a", x"9c", x"99", x"94", x"8f", x"91", x"95", x"97", x"95", x"93", x"92", 
        x"92", x"92", x"92", x"90", x"90", x"92", x"5b", x"56", x"62", x"9b", x"92", x"91", x"90", x"8f", x"8b", 
        x"8b", x"89", x"7c", x"78", x"7b", x"79", x"76", x"77", x"79", x"79", x"79", x"7e", x"84", x"83", x"83", 
        x"81", x"80", x"7c", x"cf", x"e7", x"e2", x"e1", x"e0", x"de", x"de", x"df", x"e0", x"e1", x"e1", x"df", 
        x"dd", x"dd", x"dd", x"d9", x"d6", x"d1", x"ca", x"c4", x"bf", x"bf", x"c2", x"c7", x"d1", x"d9", x"dd", 
        x"e0", x"e1", x"e0", x"df", x"de", x"de", x"de", x"df", x"dd", x"de", x"df", x"de", x"dc", x"dc", x"dc", 
        x"dc", x"dc", x"dd", x"dc", x"dc", x"dd", x"dd", x"dd", x"dd", x"de", x"dd", x"dc", x"dc", x"dc", x"dd", 
        x"dd", x"dd", x"dc", x"dc", x"dc", x"dc", x"db", x"dc", x"dc", x"dc", x"db", x"db", x"dc", x"dc", x"dc", 
        x"dd", x"dd", x"dd", x"dc", x"db", x"da", x"db", x"dd", x"dc", x"db", x"dc", x"dd", x"dd", x"dc", x"dd", 
        x"a6", x"a4", x"a3", x"a2", x"a2", x"a4", x"a5", x"a3", x"a3", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", 
        x"a4", x"a4", x"a4", x"a3", x"a2", x"a3", x"a5", x"a4", x"a4", x"a3", x"a3", x"a3", x"a4", x"a5", x"a5", 
        x"a4", x"a4", x"a4", x"a4", x"a5", x"a4", x"a3", x"a3", x"a3", x"a3", x"a4", x"a5", x"a5", x"a5", x"a5", 
        x"a5", x"a4", x"a4", x"a5", x"a5", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a5", x"a5", x"a4", x"a4", 
        x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a4", x"a5", x"a6", x"a6", 
        x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a6", x"a7", x"a8", x"a6", x"a7", 
        x"a7", x"c9", x"d2", x"cf", x"d0", x"d2", x"cf", x"d6", x"d1", x"d1", x"d4", x"d6", x"d4", x"d3", x"d1", 
        x"d4", x"d4", x"d2", x"d3", x"d3", x"d1", x"d2", x"d3", x"d2", x"d2", x"d3", x"d3", x"d3", x"d3", x"d3", 
        x"d3", x"d2", x"d1", x"d6", x"c9", x"98", x"88", x"8a", x"8c", x"87", x"85", x"8d", x"8f", x"91", x"89", 
        x"71", x"5c", x"ae", x"e2", x"d6", x"d7", x"d3", x"d2", x"e1", x"d5", x"d0", x"cf", x"d1", x"cc", x"d0", 
        x"d2", x"d0", x"d5", x"d4", x"d2", x"d0", x"d1", x"d3", x"d2", x"d2", x"d1", x"d1", x"d1", x"d2", x"d0", 
        x"d0", x"d4", x"d6", x"d4", x"d1", x"d0", x"d2", x"d2", x"d1", x"d1", x"d2", x"d4", x"d4", x"d2", x"d3", 
        x"d4", x"d2", x"d2", x"d3", x"d0", x"d2", x"d4", x"d4", x"d6", x"d6", x"dd", x"d5", x"d5", x"d9", x"da", 
        x"d6", x"d7", x"d8", x"ec", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"ee", x"ef", x"f0", x"f0", 
        x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f2", x"e9", x"ec", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"f0", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f3", x"f4", x"f4", 
        x"f3", x"f1", x"f0", x"f1", x"f2", x"f5", x"f4", x"f1", x"f0", x"f0", x"f0", x"ef", x"f3", x"f4", x"f4", 
        x"f2", x"ed", x"e1", x"d3", x"c1", x"b1", x"a8", x"a5", x"aa", x"b5", x"be", x"c6", x"d1", x"d9", x"e3", 
        x"ec", x"f1", x"f4", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f0", x"ec", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f3", x"f1", 
        x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f4", x"f3", x"f3", x"f6", x"f4", x"f4", x"f5", x"f8", x"fa", x"f8", x"f3", x"f3", x"f4", x"f2", x"f0", 
        x"f1", x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"ee", x"ef", x"f3", x"f2", x"f0", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f1", 
        x"f0", x"f0", x"f0", x"ef", x"f3", x"f7", x"f7", x"f2", x"f1", x"f6", x"f6", x"f5", x"f6", x"f9", x"f7", 
        x"f5", x"c2", x"53", x"52", x"7f", x"d2", x"d6", x"d5", x"d7", x"dc", x"c8", x"a3", x"a4", x"9e", x"8d", 
        x"7b", x"71", x"74", x"7c", x"84", x"89", x"90", x"96", x"99", x"99", x"99", x"99", x"95", x"91", x"90", 
        x"92", x"92", x"92", x"90", x"93", x"92", x"5e", x"57", x"60", x"9a", x"96", x"97", x"93", x"90", x"8a", 
        x"8b", x"8a", x"7c", x"77", x"7b", x"7a", x"77", x"77", x"79", x"79", x"78", x"7c", x"83", x"83", x"85", 
        x"83", x"82", x"7a", x"ca", x"e5", x"e1", x"e3", x"e4", x"e4", x"e4", x"e2", x"df", x"da", x"d5", x"d1", 
        x"ce", x"c7", x"c0", x"bf", x"be", x"c1", x"c9", x"d4", x"dd", x"e3", x"e2", x"e0", x"df", x"de", x"dd", 
        x"dc", x"df", x"df", x"df", x"de", x"de", x"dd", x"dd", x"dc", x"dd", x"e0", x"e0", x"df", x"de", x"de", 
        x"dd", x"de", x"df", x"de", x"dd", x"dc", x"de", x"dd", x"de", x"de", x"de", x"dc", x"dd", x"dd", x"de", 
        x"de", x"de", x"dd", x"dd", x"dd", x"dd", x"db", x"db", x"dc", x"dd", x"dc", x"db", x"db", x"dc", x"dd", 
        x"dc", x"db", x"db", x"db", x"dc", x"dc", x"dd", x"df", x"de", x"de", x"df", x"db", x"d2", x"cc", x"bf", 
        x"a6", x"a5", x"a4", x"a3", x"a3", x"a3", x"a5", x"a4", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", x"a3", 
        x"a4", x"a4", x"a4", x"a3", x"a3", x"a4", x"a5", x"a5", x"a4", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", 
        x"a4", x"a4", x"a5", x"a5", x"a5", x"a4", x"a3", x"a2", x"a3", x"a4", x"a4", x"a5", x"a5", x"a5", x"a5", 
        x"a5", x"a4", x"a4", x"a5", x"a6", x"a5", x"a4", x"a4", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a4", 
        x"a5", x"a5", x"a5", x"a6", x"a7", x"a7", x"a7", x"a6", x"a5", x"a5", x"a4", x"a4", x"a5", x"a5", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a5", x"a5", x"a5", x"a6", x"a7", 
        x"a6", x"a6", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a6", x"a6", x"a8", x"a9", x"a8", 
        x"a4", x"ca", x"d2", x"d1", x"cf", x"d2", x"d2", x"d7", x"d0", x"d1", x"d5", x"d3", x"d1", x"d3", x"d1", 
        x"d1", x"d2", x"d2", x"d2", x"d3", x"d1", x"d2", x"d4", x"d2", x"d3", x"d3", x"d2", x"d2", x"d3", x"d3", 
        x"d3", x"d3", x"d1", x"d5", x"cb", x"99", x"87", x"8b", x"8f", x"8f", x"8e", x"8d", x"78", x"5b", x"41", 
        x"28", x"2e", x"a1", x"e5", x"d7", x"d7", x"d5", x"d4", x"e1", x"d6", x"cf", x"cf", x"d1", x"ce", x"d0", 
        x"d1", x"d1", x"d5", x"d4", x"d2", x"d1", x"d2", x"d3", x"d3", x"d2", x"d0", x"d0", x"d1", x"d1", x"d1", 
        x"d1", x"d3", x"d4", x"d2", x"d1", x"d2", x"d4", x"d4", x"d3", x"d1", x"d1", x"d3", x"d3", x"d2", x"d4", 
        x"d4", x"d2", x"d3", x"d4", x"d2", x"d3", x"d4", x"d5", x"d5", x"d5", x"dc", x"d5", x"d7", x"d9", x"da", 
        x"d8", x"d7", x"d9", x"ec", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", 
        x"ed", x"ec", x"ed", x"ee", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f2", x"e8", x"eb", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f3", x"f0", x"f1", x"f2", x"f2", x"f1", x"f2", x"f1", x"f0", 
        x"f1", x"f3", x"f3", x"f1", x"ef", x"ed", x"e8", x"e2", x"d8", x"cb", x"be", x"b5", x"b1", x"b3", x"b6", 
        x"bc", x"c3", x"ca", x"d0", x"dd", x"e6", x"ee", x"f2", x"f3", x"f2", x"f3", x"f3", x"f2", x"ee", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f1", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f4", x"f3", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f4", x"f8", x"f8", x"f6", x"f3", x"f2", x"f3", x"f2", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f0", x"f2", x"f2", x"ee", x"ef", x"f4", x"f2", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f4", x"f4", x"f5", x"f1", x"f0", x"f5", x"f5", x"f5", x"f6", x"f6", x"f7", 
        x"f8", x"c9", x"58", x"52", x"7b", x"d1", x"d8", x"d5", x"d4", x"d8", x"c7", x"9d", x"a5", x"a4", x"a1", 
        x"a0", x"9b", x"94", x"8e", x"7f", x"74", x"74", x"79", x"80", x"85", x"8a", x"91", x"96", x"98", x"95", 
        x"93", x"93", x"92", x"90", x"91", x"93", x"60", x"57", x"5e", x"96", x"96", x"99", x"95", x"91", x"8c", 
        x"8c", x"8b", x"7d", x"77", x"7a", x"7a", x"79", x"79", x"78", x"78", x"77", x"7c", x"82", x"82", x"84", 
        x"83", x"83", x"78", x"c4", x"e7", x"de", x"db", x"d5", x"d2", x"d0", x"cd", x"c8", x"c4", x"c3", x"c7", 
        x"cb", x"cf", x"d5", x"dc", x"e0", x"e0", x"e0", x"e1", x"e1", x"e0", x"de", x"dd", x"de", x"df", x"e0", 
        x"e0", x"de", x"de", x"df", x"df", x"df", x"de", x"de", x"df", x"df", x"df", x"de", x"dd", x"de", x"de", 
        x"dd", x"dd", x"de", x"de", x"dd", x"dd", x"df", x"df", x"de", x"de", x"de", x"dd", x"dc", x"dc", x"dd", 
        x"de", x"de", x"dd", x"dd", x"dd", x"dd", x"dd", x"dc", x"dc", x"dd", x"dc", x"da", x"da", x"dc", x"dd", 
        x"dd", x"df", x"df", x"e1", x"e1", x"dd", x"d7", x"cc", x"c0", x"b1", x"9d", x"8a", x"7c", x"6e", x"62", 
        x"a5", x"a5", x"a5", x"a3", x"a2", x"a2", x"a3", x"a5", x"a4", x"a3", x"a3", x"a4", x"a3", x"a2", x"a2", 
        x"a2", x"a3", x"a3", x"a4", x"a4", x"a4", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", x"a3", x"a3", x"a3", 
        x"a4", x"a5", x"a6", x"a6", x"a5", x"a4", x"a2", x"a2", x"a3", x"a3", x"a4", x"a5", x"a5", x"a4", x"a5", 
        x"a6", x"a5", x"a4", x"a5", x"a6", x"a5", x"a4", x"a4", x"a5", x"a6", x"a5", x"a3", x"a5", x"a7", x"a6", 
        x"a5", x"a5", x"a5", x"a6", x"a7", x"a7", x"a7", x"a6", x"a6", x"a5", x"a4", x"a4", x"a6", x"a5", x"a5", 
        x"a5", x"a7", x"a6", x"a5", x"a6", x"a6", x"a7", x"a7", x"a6", x"a5", x"a5", x"a6", x"a6", x"a7", x"a7", 
        x"a5", x"a6", x"a7", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a8", x"a5", x"a7", x"a9", x"a6", 
        x"a4", x"cc", x"d3", x"d0", x"d1", x"d2", x"d0", x"d6", x"d1", x"d1", x"d4", x"d3", x"d1", x"d0", x"d0", 
        x"d1", x"d2", x"d2", x"d2", x"d4", x"d2", x"d0", x"d3", x"d2", x"d1", x"d2", x"d0", x"d2", x"d2", x"d1", 
        x"d3", x"d3", x"d3", x"d2", x"c9", x"9b", x"8f", x"93", x"8f", x"80", x"63", x"48", x"2c", x"13", x"0e", 
        x"16", x"35", x"a6", x"e3", x"d5", x"d8", x"d9", x"d2", x"e0", x"d7", x"ce", x"d0", x"d2", x"d1", x"d1", 
        x"cf", x"d2", x"d6", x"d7", x"d6", x"d4", x"d2", x"cf", x"d2", x"d3", x"d0", x"d1", x"d1", x"d1", x"d2", 
        x"d2", x"d3", x"d2", x"d1", x"cf", x"d0", x"d2", x"d4", x"d5", x"d3", x"d2", x"d5", x"d5", x"d4", x"d4", 
        x"d3", x"d3", x"d4", x"d4", x"d4", x"d3", x"d4", x"d6", x"d4", x"d5", x"db", x"d5", x"d7", x"da", x"da", 
        x"da", x"d6", x"d7", x"ed", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ee", 
        x"ec", x"eb", x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"ee", x"ee", x"ed", x"ef", x"f1", x"f0", x"e8", x"ea", 
        x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"ef", x"ef", x"f1", x"f2", x"f4", x"f5", x"f7", x"f4", x"e9", x"de", x"d0", 
        x"c2", x"b6", x"b0", x"ae", x"b2", x"b8", x"ba", x"c2", x"cc", x"d8", x"e6", x"ee", x"f2", x"f1", x"f4", 
        x"f5", x"f4", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f0", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", 
        x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f6", x"f7", x"f5", x"f3", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f1", x"f0", x"ef", x"f1", x"f3", x"f2", x"ee", x"f1", x"f3", x"f2", x"f3", x"f2", x"f3", x"f4", 
        x"f2", x"f2", x"f1", x"f2", x"f1", x"ef", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f3", x"f4", x"f2", x"f6", x"f2", x"ef", x"f6", x"f6", x"f6", x"f8", x"f5", x"f6", 
        x"f7", x"d0", x"5f", x"54", x"75", x"cc", x"da", x"d8", x"d5", x"d8", x"ca", x"9c", x"a4", x"a3", x"9a", 
        x"9c", x"9a", x"9f", x"a3", x"a5", x"9b", x"94", x"8e", x"80", x"74", x"72", x"76", x"7d", x"83", x"88", 
        x"8e", x"95", x"99", x"97", x"94", x"95", x"61", x"57", x"5f", x"95", x"96", x"99", x"93", x"8f", x"8c", 
        x"8c", x"8b", x"80", x"77", x"79", x"78", x"79", x"7a", x"77", x"77", x"77", x"7d", x"82", x"81", x"83", 
        x"83", x"81", x"76", x"ab", x"ce", x"c3", x"c3", x"c2", x"c0", x"c7", x"cc", x"d4", x"db", x"e0", x"e3", 
        x"e5", x"e5", x"e2", x"e0", x"df", x"de", x"de", x"df", x"e0", x"e0", x"df", x"df", x"df", x"df", x"df", 
        x"e0", x"de", x"df", x"e0", x"e0", x"df", x"de", x"de", x"e0", x"e0", x"e0", x"df", x"de", x"dd", x"dd", 
        x"db", x"dc", x"dc", x"dc", x"dc", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", x"dd", x"dd", x"dc", x"dc", 
        x"dd", x"de", x"de", x"de", x"dc", x"db", x"db", x"dc", x"dc", x"dc", x"de", x"e0", x"e3", x"e4", x"e0", 
        x"da", x"d4", x"c6", x"b8", x"a7", x"94", x"83", x"72", x"63", x"58", x"49", x"42", x"44", x"43", x"47", 
        x"a6", x"a5", x"a4", x"a4", x"a4", x"a3", x"a3", x"a5", x"a4", x"a3", x"a3", x"a4", x"a4", x"a3", x"a3", 
        x"a2", x"a3", x"a3", x"a4", x"a3", x"a3", x"a2", x"a2", x"a4", x"a5", x"a5", x"a4", x"a3", x"a3", x"a3", 
        x"a4", x"a5", x"a5", x"a5", x"a4", x"a4", x"a5", x"a5", x"a5", x"a4", x"a4", x"a5", x"a5", x"a4", x"a5", 
        x"a5", x"a5", x"a4", x"a5", x"a6", x"a4", x"a4", x"a5", x"a5", x"a5", x"a4", x"a4", x"a6", x"a7", x"a6", 
        x"a5", x"a5", x"a5", x"a6", x"a5", x"a4", x"a5", x"a7", x"a7", x"a7", x"a6", x"a5", x"a6", x"a5", x"a5", 
        x"a6", x"a7", x"a6", x"a5", x"a4", x"a5", x"a6", x"a7", x"a7", x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", 
        x"a6", x"a6", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a5", x"a6", x"a7", x"a6", 
        x"a3", x"ca", x"d2", x"d0", x"d3", x"d3", x"cf", x"d3", x"d1", x"d3", x"d4", x"d4", x"d3", x"d2", x"d2", 
        x"d2", x"d2", x"d2", x"d1", x"d4", x"d3", x"d1", x"d3", x"d2", x"d1", x"d4", x"cf", x"d0", x"d0", x"d0", 
        x"d2", x"d0", x"d3", x"dc", x"d4", x"a2", x"7a", x"5a", x"3f", x"27", x"13", x"0e", x"18", x"28", x"37", 
        x"3e", x"4b", x"ad", x"e5", x"d4", x"d4", x"d6", x"d3", x"e0", x"d7", x"cf", x"d2", x"d4", x"d4", x"d4", 
        x"d2", x"d1", x"d3", x"d4", x"d4", x"d2", x"d0", x"cf", x"d2", x"d2", x"d1", x"d3", x"d0", x"cf", x"d1", 
        x"d3", x"d3", x"d3", x"d3", x"d2", x"d1", x"d0", x"d1", x"d3", x"d5", x"d5", x"d7", x"d7", x"d5", x"d2", 
        x"d3", x"d5", x"d6", x"d5", x"d3", x"d2", x"d4", x"d6", x"d4", x"d5", x"db", x"d5", x"d8", x"db", x"da", 
        x"da", x"d6", x"d5", x"ed", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ee", x"f0", x"f0", x"e9", x"ea", 
        x"f2", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"f2", x"f5", 
        x"f6", x"f2", x"ed", x"e6", x"da", x"d4", x"c7", x"bf", x"b9", x"b5", x"b4", x"b1", x"b6", x"bd", x"cc", 
        x"db", x"e7", x"ee", x"f4", x"f5", x"f5", x"f5", x"f4", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", x"f4", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f5", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f5", x"f6", x"f5", x"f3", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"ed", x"f0", x"f3", x"f2", x"f3", x"f3", x"f2", x"f3", 
        x"f2", x"f2", x"f1", x"f2", x"f1", x"f0", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f5", x"f6", x"f4", x"f7", x"f3", x"f0", x"f5", x"f5", x"f4", x"f7", x"f6", x"f5", 
        x"f8", x"d3", x"61", x"52", x"70", x"c9", x"d9", x"d6", x"d6", x"da", x"cd", x"9e", x"a2", x"ac", x"a7", 
        x"9c", x"99", x"9c", x"9c", x"9a", x"9a", x"9a", x"9c", x"9c", x"99", x"93", x"8e", x"84", x"7a", x"75", 
        x"70", x"70", x"78", x"83", x"8f", x"9b", x"67", x"53", x"58", x"91", x"97", x"99", x"96", x"93", x"8f", 
        x"8c", x"8d", x"81", x"77", x"7b", x"79", x"79", x"7a", x"79", x"79", x"76", x"7b", x"81", x"81", x"84", 
        x"84", x"83", x"72", x"99", x"c8", x"d0", x"d8", x"dc", x"dc", x"e0", x"e3", x"e4", x"e3", x"e2", x"e1", 
        x"e2", x"e1", x"df", x"df", x"df", x"df", x"df", x"e0", x"e0", x"df", x"e0", x"df", x"df", x"df", x"df", 
        x"df", x"de", x"de", x"df", x"e0", x"df", x"de", x"df", x"e0", x"de", x"dd", x"de", x"df", x"de", x"dd", 
        x"dd", x"dd", x"dc", x"db", x"db", x"dc", x"dc", x"db", x"db", x"dc", x"dd", x"de", x"de", x"dc", x"db", 
        x"dc", x"db", x"db", x"dc", x"de", x"e0", x"e2", x"e4", x"e5", x"e1", x"d7", x"c9", x"b2", x"9d", x"8b", 
        x"75", x"68", x"60", x"5c", x"59", x"54", x"4e", x"4b", x"45", x"45", x"44", x"44", x"46", x"48", x"3e", 
        x"a8", x"a6", x"a5", x"a5", x"a5", x"a5", x"a4", x"a5", x"a4", x"a3", x"a4", x"a5", x"a4", x"a3", x"a3", 
        x"a2", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a3", x"a4", x"a5", x"a6", x"a5", x"a4", x"a3", x"a3", 
        x"a3", x"a4", x"a4", x"a4", x"a4", x"a4", x"a6", x"a6", x"a6", x"a6", x"a5", x"a6", x"a5", x"a4", x"a5", 
        x"a5", x"a5", x"a5", x"a6", x"a6", x"a4", x"a5", x"a6", x"a6", x"a5", x"a4", x"a5", x"a7", x"a7", x"a7", 
        x"a6", x"a6", x"a6", x"a6", x"a5", x"a4", x"a6", x"a7", x"a7", x"a6", x"a5", x"a5", x"a6", x"a6", x"a6", 
        x"a6", x"a7", x"a7", x"a5", x"a4", x"a5", x"a6", x"a7", x"a6", x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", 
        x"a6", x"a6", x"a7", x"a7", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a7", x"a5", x"a6", x"a7", x"a6", 
        x"a2", x"c9", x"d2", x"d1", x"d3", x"d3", x"cf", x"d2", x"d2", x"d4", x"d5", x"d4", x"d3", x"d3", x"d2", 
        x"d2", x"d3", x"d2", x"d1", x"d5", x"d4", x"d1", x"d2", x"d2", x"cf", x"d4", x"d1", x"cf", x"cf", x"d3", 
        x"d8", x"d6", x"d0", x"b8", x"91", x"53", x"2e", x"1d", x"15", x"18", x"25", x"34", x"41", x"4a", x"52", 
        x"51", x"4d", x"a8", x"e4", x"d6", x"d5", x"d7", x"d4", x"df", x"d6", x"ce", x"d1", x"d4", x"d3", x"d3", 
        x"d3", x"d2", x"d2", x"d2", x"d3", x"d2", x"d0", x"cf", x"d0", x"cf", x"d0", x"d4", x"d1", x"ce", x"d1", 
        x"d3", x"d3", x"d3", x"d4", x"d3", x"d1", x"cf", x"d1", x"d3", x"d5", x"d6", x"d5", x"d5", x"d3", x"d1", 
        x"d4", x"d6", x"d6", x"d5", x"d3", x"d2", x"d4", x"d6", x"d5", x"d6", x"dc", x"d5", x"d8", x"da", x"da", 
        x"da", x"d5", x"d5", x"ed", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f1", x"f2", x"e9", x"e9", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f3", x"f5", x"f4", x"f1", x"ed", x"e7", x"de", x"d6", x"cd", x"c9", x"c0", x"bf", 
        x"bf", x"be", x"be", x"c1", x"c9", x"d5", x"e2", x"ec", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f3", x"f2", x"f0", x"f1", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f5", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f5", x"f5", x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f0", x"ed", x"f0", x"f3", x"f1", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f3", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f1", x"f2", x"f2", x"f5", x"f3", x"f0", x"f5", x"f5", x"f4", x"f6", x"f7", x"f5", 
        x"f9", x"d8", x"68", x"52", x"6c", x"c7", x"d9", x"d4", x"d6", x"da", x"ce", x"9e", x"a0", x"b3", x"ba", 
        x"9c", x"99", x"9d", x"99", x"9a", x"9c", x"99", x"96", x"97", x"9b", x"9b", x"9d", x"98", x"92", x"90", 
        x"8c", x"83", x"7a", x"71", x"6f", x"7a", x"5a", x"54", x"5c", x"8d", x"96", x"99", x"9a", x"98", x"92", 
        x"8d", x"8c", x"81", x"77", x"7c", x"7a", x"79", x"7a", x"7a", x"7c", x"77", x"7b", x"80", x"81", x"83", 
        x"84", x"84", x"73", x"a3", x"e3", x"e5", x"e4", x"e4", x"e2", x"e1", x"e1", x"e0", x"df", x"df", x"df", 
        x"e0", x"df", x"de", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"e0", x"e0", x"e0", x"df", 
        x"de", x"dd", x"dd", x"de", x"df", x"df", x"df", x"df", x"df", x"de", x"de", x"df", x"df", x"e0", x"df", 
        x"de", x"de", x"dd", x"dc", x"dc", x"dc", x"db", x"dd", x"de", x"dd", x"dd", x"db", x"dc", x"dd", x"de", 
        x"df", x"e0", x"e0", x"dd", x"d5", x"cb", x"c0", x"af", x"9c", x"85", x"74", x"66", x"5c", x"58", x"56", 
        x"4e", x"4f", x"4b", x"46", x"45", x"4a", x"4a", x"49", x"4a", x"4a", x"43", x"42", x"3d", x"37", x"28", 
        x"a8", x"a6", x"a5", x"a5", x"a6", x"a5", x"a4", x"a5", x"a5", x"a4", x"a4", x"a5", x"a4", x"a3", x"a3", 
        x"a2", x"a3", x"a4", x"a3", x"a3", x"a2", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a4", x"a3", 
        x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", x"a5", x"a5", x"a5", x"a6", x"a6", x"a7", x"a7", x"a5", x"a5", 
        x"a4", x"a5", x"a5", x"a6", x"a6", x"a4", x"a5", x"a6", x"a5", x"a4", x"a4", x"a5", x"a7", x"a7", x"a7", 
        x"a7", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a5", x"a5", x"a6", x"a7", x"a6", 
        x"a6", x"a7", x"a7", x"a6", x"a5", x"a6", x"a6", x"a7", x"a6", x"a5", x"a5", x"a6", x"a6", x"a6", x"a7", 
        x"a7", x"a7", x"a6", x"a7", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a7", x"a7", x"a8", x"a7", x"a8", 
        x"a4", x"c9", x"d4", x"d2", x"d2", x"d1", x"d0", x"d4", x"d4", x"d3", x"d5", x"d4", x"d2", x"d1", x"d1", 
        x"d3", x"d4", x"cf", x"ce", x"d2", x"d5", x"d3", x"d2", x"ce", x"d1", x"d5", x"d1", x"d6", x"df", x"de", 
        x"ca", x"9e", x"68", x"39", x"21", x"11", x"14", x"21", x"32", x"43", x"51", x"59", x"57", x"52", x"52", 
        x"4e", x"4d", x"a4", x"e3", x"d6", x"d5", x"d8", x"d5", x"e0", x"d6", x"ce", x"d1", x"d2", x"d1", x"d2", 
        x"d3", x"d2", x"d1", x"d1", x"d2", x"d2", x"d0", x"d1", x"d2", x"d0", x"d0", x"d3", x"cf", x"cd", x"d0", 
        x"d2", x"d2", x"d2", x"d3", x"d3", x"d0", x"ce", x"d0", x"d2", x"d3", x"d4", x"d2", x"d4", x"d4", x"d2", 
        x"d4", x"d6", x"d5", x"d3", x"d2", x"d3", x"d4", x"d6", x"d5", x"d6", x"dc", x"d5", x"d7", x"d9", x"d9", 
        x"da", x"d7", x"d7", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f2", x"f2", x"ea", x"e9", 
        x"f1", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"f0", x"f1", x"f1", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f0", x"f1", x"f5", x"f4", x"f3", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"ea", x"eb", 
        x"e9", x"e2", x"dd", x"ce", x"c3", x"ba", x"b5", x"b5", x"bb", x"c1", x"cf", x"dc", x"e7", x"f1", x"f6", 
        x"f6", x"f4", x"f0", x"ef", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f4", x"f5", x"f5", x"f5", x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f4", x"f4", x"f4", x"f2", x"f2", x"f1", x"f0", x"ed", x"f0", x"f2", x"f1", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f2", x"f1", x"ef", x"f4", x"f6", x"f6", x"f6", x"f6", x"f5", 
        x"fa", x"df", x"72", x"53", x"6b", x"c4", x"da", x"d4", x"d6", x"d8", x"cf", x"9e", x"9e", x"b4", x"ce", 
        x"a7", x"97", x"9e", x"98", x"9a", x"98", x"95", x"94", x"99", x"9b", x"99", x"93", x"95", x"95", x"93", 
        x"93", x"95", x"92", x"91", x"8a", x"88", x"64", x"54", x"53", x"75", x"84", x"8e", x"95", x"98", x"94", 
        x"90", x"90", x"84", x"76", x"7b", x"78", x"76", x"77", x"77", x"7a", x"79", x"7c", x"80", x"81", x"83", 
        x"83", x"83", x"72", x"a4", x"e3", x"dc", x"e0", x"e3", x"e2", x"e1", x"e0", x"e0", x"e1", x"e2", x"e2", 
        x"e3", x"e1", x"de", x"df", x"e0", x"e0", x"df", x"de", x"de", x"df", x"df", x"e0", x"e1", x"e0", x"df", 
        x"de", x"dd", x"de", x"de", x"de", x"df", x"e0", x"e0", x"dd", x"de", x"e0", x"e1", x"e0", x"df", x"de", 
        x"df", x"de", x"dd", x"dd", x"de", x"dc", x"db", x"dc", x"de", x"df", x"e1", x"e5", x"e5", x"e3", x"dd", 
        x"cf", x"bd", x"a3", x"88", x"71", x"5f", x"56", x"55", x"51", x"51", x"51", x"4e", x"4d", x"4d", x"47", 
        x"42", x"3a", x"2c", x"20", x"23", x"32", x"41", x"3b", x"33", x"27", x"19", x"17", x"15", x"0f", x"0a", 
        x"a8", x"a6", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a4", x"a4", x"a5", x"a5", x"a4", x"a4", 
        x"a4", x"a4", x"a4", x"a4", x"a3", x"a3", x"a4", x"a6", x"a4", x"a3", x"a3", x"a4", x"a5", x"a6", x"a4", 
        x"a4", x"a4", x"a4", x"a4", x"a5", x"a6", x"a4", x"a4", x"a4", x"a5", x"a6", x"a7", x"a7", x"a5", x"a4", 
        x"a4", x"a5", x"a6", x"a6", x"a5", x"a5", x"a6", x"a6", x"a5", x"a5", x"a5", x"a6", x"a7", x"a7", x"a7", 
        x"a8", x"a8", x"a7", x"a6", x"a6", x"a6", x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a7", x"a7", 
        x"a7", x"a6", x"a6", x"a7", x"a7", x"a8", x"a8", x"a7", x"a6", x"a5", x"a5", x"a6", x"a7", x"a6", x"a6", 
        x"a7", x"a7", x"a6", x"a7", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a7", x"a8", x"a9", x"a7", x"a8", 
        x"a4", x"c8", x"d4", x"d3", x"d1", x"d1", x"d2", x"d6", x"d4", x"d1", x"d4", x"d3", x"d2", x"d1", x"d1", 
        x"d2", x"d3", x"d4", x"d4", x"d3", x"ce", x"cd", x"d3", x"d4", x"d5", x"d6", x"d2", x"bc", x"98", x"69", 
        x"38", x"25", x"20", x"1e", x"28", x"37", x"47", x"4f", x"55", x"56", x"54", x"51", x"50", x"51", x"52", 
        x"4c", x"4a", x"a5", x"e5", x"d5", x"d6", x"d8", x"d5", x"e3", x"d9", x"d0", x"d2", x"d4", x"d2", x"d2", 
        x"d2", x"d1", x"d2", x"d2", x"d2", x"d1", x"d0", x"d1", x"d3", x"d2", x"d0", x"d2", x"d0", x"d0", x"d2", 
        x"d2", x"d2", x"d2", x"d2", x"d1", x"d0", x"cf", x"d3", x"d3", x"d3", x"d3", x"ce", x"d2", x"d3", x"d3", 
        x"d5", x"d5", x"d5", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d6", x"dc", x"d4", x"d6", x"d7", x"d8", 
        x"db", x"d8", x"d7", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"f1", x"ea", x"e9", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f3", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"ef", x"f0", x"f3", x"f2", x"f1", x"f2", x"f2", x"f4", x"f3", x"ed", x"ef", 
        x"f2", x"f2", x"f0", x"f0", x"ef", x"ed", x"e9", x"e1", x"d7", x"cf", x"c3", x"bb", x"b8", x"b7", x"bd", 
        x"c8", x"d3", x"e1", x"ea", x"ee", x"f0", x"f0", x"f1", x"f2", x"f4", x"f3", x"f2", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f4", x"f5", x"f6", x"f4", x"f4", x"f5", x"f5", x"f4", x"f3", x"f3", x"f5", 
        x"f6", x"f5", x"f4", x"f2", x"f2", x"f1", x"f0", x"ed", x"ef", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f2", x"f3", x"f1", x"f1", x"f2", x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f1", x"f2", x"f3", x"f0", x"f1", x"ef", x"ef", x"f3", x"f7", x"f7", x"f6", x"f5", x"f5", 
        x"f9", x"e3", x"7b", x"53", x"69", x"c1", x"db", x"d4", x"d5", x"d6", x"d0", x"a1", x"9f", x"af", x"d7", 
        x"c2", x"9a", x"9c", x"99", x"97", x"9b", x"9f", x"9d", x"99", x"97", x"98", x"97", x"97", x"97", x"95", 
        x"93", x"93", x"94", x"94", x"92", x"9a", x"73", x"54", x"59", x"7b", x"80", x"7c", x"7c", x"7a", x"77", 
        x"7c", x"87", x"83", x"79", x"7a", x"79", x"7a", x"79", x"7a", x"7e", x"7b", x"7b", x"80", x"82", x"83", 
        x"82", x"81", x"71", x"9d", x"e3", x"de", x"e1", x"e0", x"e0", x"e0", x"df", x"df", x"e1", x"e2", x"e3", 
        x"e2", x"e0", x"df", x"e0", x"e0", x"e0", x"df", x"de", x"de", x"df", x"e0", x"e0", x"e0", x"e0", x"df", 
        x"df", x"df", x"de", x"de", x"de", x"de", x"df", x"e0", x"df", x"df", x"df", x"dd", x"dd", x"df", x"e0", 
        x"e1", x"e0", x"de", x"df", x"e0", x"df", x"dd", x"db", x"d3", x"c5", x"b7", x"a4", x"8c", x"73", x"60", 
        x"57", x"53", x"50", x"52", x"53", x"54", x"52", x"51", x"53", x"4f", x"49", x"44", x"3f", x"37", x"23", 
        x"16", x"0c", x"07", x"08", x"08", x"0c", x"0e", x"0f", x"12", x"0e", x"11", x"12", x"15", x"23", x"3b", 
        x"a6", x"a6", x"a6", x"a5", x"a4", x"a4", x"a5", x"a6", x"a5", x"a4", x"a5", x"a5", x"a5", x"a4", x"a5", 
        x"a5", x"a5", x"a5", x"a4", x"a3", x"a3", x"a4", x"a5", x"a5", x"a4", x"a4", x"a5", x"a5", x"a5", x"a5", 
        x"a4", x"a4", x"a4", x"a4", x"a5", x"a6", x"a4", x"a4", x"a4", x"a5", x"a5", x"a6", x"a6", x"a5", x"a4", 
        x"a3", x"a4", x"a6", x"a6", x"a5", x"a6", x"a6", x"a5", x"a4", x"a5", x"a6", x"a6", x"a6", x"a7", x"a7", 
        x"a8", x"a8", x"a7", x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a5", x"a5", x"a6", x"a8", x"a8", 
        x"a7", x"a6", x"a6", x"a7", x"a7", x"a7", x"a8", x"a8", x"a7", x"a7", x"a7", x"a7", x"a6", x"a6", x"a6", 
        x"a7", x"a7", x"a6", x"a7", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a7", x"a8", x"a9", x"a6", x"a8", 
        x"a3", x"c7", x"d3", x"d1", x"d2", x"d3", x"d3", x"d4", x"d4", x"d1", x"d2", x"d3", x"d3", x"d3", x"d3", 
        x"d2", x"d2", x"d1", x"d3", x"d6", x"d3", x"d5", x"d9", x"d3", x"c6", x"a2", x"6f", x"3a", x"20", x"1a", 
        x"23", x"33", x"3b", x"43", x"50", x"59", x"55", x"52", x"54", x"51", x"50", x"4e", x"4d", x"4c", x"4c", 
        x"44", x"43", x"a4", x"e6", x"d4", x"d7", x"d9", x"d4", x"e1", x"d7", x"cf", x"d2", x"d3", x"d3", x"d3", 
        x"d0", x"d1", x"d2", x"d2", x"d2", x"d1", x"d1", x"d0", x"d1", x"d3", x"d0", x"d3", x"d3", x"d3", x"d4", 
        x"d3", x"d3", x"d3", x"d1", x"d1", x"d1", x"d2", x"d6", x"d6", x"d5", x"d4", x"cd", x"d1", x"d3", x"d4", 
        x"d4", x"d4", x"d5", x"d5", x"d4", x"d3", x"d2", x"d4", x"d4", x"d6", x"db", x"d4", x"d5", x"d7", x"d8", 
        x"da", x"d7", x"d7", x"ed", x"ed", x"ed", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ee", x"ed", x"ec", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f1", x"f0", x"f0", x"f0", x"ed", x"ed", x"f1", x"ea", x"e8", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f0", x"ef", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f5", x"f3", x"f2", x"f3", x"f1", x"f3", x"f2", x"ec", x"f0", 
        x"f3", x"f3", x"f2", x"f3", x"f4", x"f3", x"f3", x"f2", x"f0", x"ef", x"ef", x"ed", x"e8", x"e0", x"d1", 
        x"c4", x"b9", x"b8", x"bd", x"bf", x"c4", x"cb", x"d7", x"e4", x"ec", x"ee", x"ef", x"f1", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", 
        x"f5", x"f5", x"f3", x"f3", x"f3", x"f5", x"f6", x"f4", x"f4", x"f5", x"f5", x"f4", x"f4", x"f3", x"f6", 
        x"f8", x"f6", x"f3", x"f1", x"f1", x"f1", x"f0", x"ed", x"ef", x"f2", x"f0", x"f2", x"f1", x"f1", x"f1", 
        x"f3", x"f4", x"f2", x"f2", x"f3", x"f4", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"ef", x"f2", x"f6", x"f6", x"f6", x"f4", x"f5", 
        x"f6", x"e4", x"80", x"50", x"66", x"bd", x"db", x"d4", x"d6", x"d5", x"d2", x"a4", x"9f", x"ac", x"d5", 
        x"d5", x"a7", x"98", x"9a", x"9b", x"9b", x"9a", x"98", x"99", x"9a", x"9a", x"98", x"97", x"96", x"96", 
        x"93", x"92", x"96", x"93", x"90", x"9b", x"75", x"4e", x"59", x"80", x"92", x"97", x"97", x"90", x"82", 
        x"76", x"71", x"6b", x"6b", x"6c", x"6e", x"75", x"76", x"78", x"7e", x"7a", x"7a", x"80", x"83", x"84", 
        x"83", x"82", x"73", x"95", x"e0", x"dd", x"e1", x"e3", x"e2", x"e1", x"e0", x"df", x"e0", x"e1", x"e1", 
        x"e0", x"df", x"de", x"df", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"df", x"df", x"df", x"df", x"e0", 
        x"e0", x"e0", x"df", x"de", x"de", x"de", x"de", x"e0", x"e2", x"e0", x"df", x"e1", x"e3", x"e1", x"de", 
        x"e0", x"de", x"d9", x"d0", x"c2", x"ad", x"9b", x"82", x"6b", x"5b", x"50", x"4d", x"52", x"58", x"5b", 
        x"5a", x"59", x"5b", x"5c", x"5b", x"57", x"55", x"55", x"50", x"40", x"30", x"22", x"17", x"0e", x"08", 
        x"06", x"06", x"0a", x"0f", x"11", x"18", x"0c", x"0d", x"2a", x"39", x"51", x"65", x"67", x"68", x"6f", 
        x"a6", x"a7", x"a7", x"a5", x"a4", x"a4", x"a5", x"a6", x"a6", x"a5", x"a6", x"a6", x"a6", x"a4", x"a5", 
        x"a5", x"a5", x"a5", x"a5", x"a4", x"a4", x"a4", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a6", 
        x"a4", x"a4", x"a4", x"a5", x"a5", x"a7", x"a7", x"a7", x"a6", x"a5", x"a5", x"a5", x"a5", x"a4", x"a4", 
        x"a4", x"a5", x"a6", x"a6", x"a6", x"a7", x"a6", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", 
        x"a8", x"a8", x"a7", x"a6", x"a6", x"a7", x"a7", x"a7", x"a7", x"a6", x"a4", x"a3", x"a6", x"a8", x"a8", 
        x"a7", x"a6", x"a7", x"a8", x"a7", x"a7", x"a8", x"a8", x"a8", x"a9", x"a9", x"a8", x"a7", x"a6", x"a7", 
        x"a8", x"a8", x"a7", x"a8", x"a9", x"a9", x"a9", x"a9", x"a9", x"a9", x"a7", x"a7", x"a8", x"a5", x"a6", 
        x"a2", x"c5", x"d2", x"d0", x"d3", x"d4", x"d4", x"d2", x"d3", x"d2", x"d2", x"d3", x"d4", x"d3", x"d4", 
        x"d3", x"d0", x"d7", x"d8", x"d6", x"d4", x"ca", x"ab", x"7a", x"49", x"23", x"19", x"1c", x"2e", x"44", 
        x"58", x"6d", x"6e", x"5e", x"55", x"56", x"52", x"50", x"52", x"50", x"4d", x"4b", x"4b", x"49", x"47", 
        x"3e", x"3f", x"a3", x"e4", x"d0", x"d4", x"d7", x"d4", x"de", x"d5", x"ce", x"d1", x"d3", x"d3", x"d2", 
        x"d1", x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", x"d0", x"d3", x"d4", x"d3", x"d3", x"d3", x"d2", x"d3", 
        x"d4", x"d4", x"d3", x"d1", x"d1", x"d1", x"d1", x"d2", x"d3", x"d4", x"d5", x"d0", x"d3", x"d5", x"d4", 
        x"d5", x"d5", x"d6", x"d6", x"d5", x"d3", x"d2", x"d4", x"d4", x"d5", x"db", x"d4", x"d4", x"d8", x"d8", 
        x"d9", x"d6", x"d7", x"ed", x"ee", x"ed", x"ef", x"f0", x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", x"ee", 
        x"ef", x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"f1", x"e9", x"e5", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f2", x"f2", x"f0", x"f2", x"f1", x"f2", x"f5", x"f3", x"f3", x"f0", x"eb", x"ee", 
        x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f2", x"f0", 
        x"ee", x"ed", x"eb", x"e5", x"da", x"ca", x"bd", x"b7", x"b7", x"bc", x"c3", x"c8", x"d0", x"d9", x"e1", 
        x"e9", x"ec", x"ee", x"f0", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f5", x"f4", x"f4", x"f4", x"f4", x"f4", x"f5", 
        x"f7", x"f6", x"f5", x"f3", x"f3", x"f4", x"f6", x"f4", x"f4", x"f5", x"f5", x"f5", x"f4", x"f3", x"f6", 
        x"f8", x"f6", x"f3", x"f1", x"f2", x"f2", x"f1", x"ee", x"ef", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f4", x"f2", x"f3", x"f4", x"f3", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"f2", x"f7", x"f6", x"f6", x"f4", x"f5", 
        x"f5", x"e5", x"84", x"4e", x"63", x"b8", x"dc", x"d4", x"d6", x"d6", x"d5", x"a6", x"9e", x"ad", x"d2", 
        x"dd", x"bf", x"9c", x"99", x"99", x"99", x"98", x"99", x"9b", x"9a", x"96", x"95", x"96", x"95", x"93", 
        x"92", x"92", x"92", x"93", x"8f", x"99", x"7c", x"50", x"55", x"74", x"8a", x"94", x"9b", x"9d", x"95", 
        x"8d", x"8b", x"7a", x"61", x"5e", x"60", x"65", x"66", x"67", x"6f", x"73", x"74", x"7e", x"85", x"85", 
        x"84", x"83", x"74", x"90", x"e3", x"de", x"df", x"e3", x"e4", x"e2", x"e2", x"e0", x"e0", x"e1", x"e3", 
        x"e1", x"df", x"de", x"de", x"e0", x"e1", x"e0", x"e0", x"e0", x"df", x"e0", x"df", x"df", x"df", x"df", 
        x"df", x"e0", x"df", x"df", x"e0", x"e2", x"e3", x"e2", x"e2", x"dc", x"d9", x"d7", x"d0", x"c0", x"b2", 
        x"a1", x"91", x"7c", x"6a", x"5d", x"55", x"55", x"57", x"5a", x"5b", x"59", x"56", x"53", x"51", x"51", 
        x"50", x"52", x"56", x"52", x"44", x"31", x"21", x"17", x"12", x"0d", x"0d", x"0d", x"12", x"19", x"20", 
        x"27", x"31", x"3e", x"4d", x"5b", x"65", x"29", x"27", x"69", x"77", x"77", x"88", x"83", x"80", x"79", 
        x"a4", x"a6", x"a7", x"a4", x"a4", x"a5", x"a4", x"a5", x"a6", x"a8", x"a8", x"a7", x"a5", x"a4", x"a3", 
        x"a2", x"a3", x"a3", x"a3", x"a4", x"a4", x"a4", x"a4", x"a5", x"a6", x"a6", x"a5", x"a4", x"a5", x"a5", 
        x"a2", x"a2", x"a4", x"a4", x"a4", x"a7", x"a9", x"a8", x"a7", x"a5", x"a4", x"a5", x"a5", x"a5", x"a5", 
        x"a5", x"a6", x"a6", x"a6", x"a7", x"a6", x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", x"a6", x"a5", x"a6", 
        x"a7", x"a7", x"a6", x"a5", x"a6", x"a7", x"a6", x"a6", x"a7", x"a7", x"a4", x"a3", x"a4", x"a5", x"a6", 
        x"a7", x"a7", x"a6", x"a6", x"a7", x"a7", x"a6", x"a6", x"a7", x"a8", x"a8", x"a9", x"a9", x"a9", x"a9", 
        x"a8", x"a7", x"a7", x"a7", x"a8", x"a8", x"a8", x"a8", x"a9", x"a9", x"a9", x"a8", x"a7", x"a6", x"a5", 
        x"a3", x"c3", x"d6", x"d1", x"d0", x"d3", x"d5", x"cf", x"d1", x"d2", x"d2", x"d3", x"d1", x"ce", x"d3", 
        x"d8", x"d8", x"da", x"d2", x"b0", x"7f", x"52", x"27", x"0a", x"10", x"25", x"3b", x"57", x"6e", x"80", 
        x"7f", x"7a", x"66", x"59", x"50", x"50", x"50", x"4d", x"4d", x"47", x"45", x"45", x"46", x"45", x"43", 
        x"3d", x"40", x"a2", x"e3", x"d3", x"d3", x"d5", x"d4", x"dd", x"d5", x"d0", x"d4", x"d7", x"d5", x"d2", 
        x"d5", x"d5", x"d3", x"d2", x"d2", x"d3", x"d3", x"d3", x"d2", x"d3", x"d4", x"d4", x"d3", x"d2", x"d3", 
        x"d4", x"d3", x"d3", x"d3", x"d2", x"d2", x"d0", x"cd", x"d0", x"d4", x"d4", x"d3", x"d3", x"d3", x"d4", 
        x"d7", x"d7", x"d5", x"d5", x"d5", x"d5", x"d3", x"d6", x"d7", x"d5", x"d9", x"d5", x"d3", x"d8", x"da", 
        x"d8", x"d5", x"d7", x"ec", x"ef", x"eb", x"ed", x"ef", x"ee", x"f0", x"ee", x"ed", x"ef", x"ed", x"ee", 
        x"f1", x"f2", x"ef", x"ee", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ee", 
        x"ee", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"ed", x"ee", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"f0", x"e9", x"e4", 
        x"f3", x"f1", x"f2", x"f3", x"f1", x"ef", x"f1", x"f1", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f3", x"f1", x"ee", x"ef", x"f1", x"f0", x"ed", x"ed", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"f1", x"f1", 
        x"f2", x"f3", x"f1", x"f0", x"ef", x"f0", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"ef", 
        x"f0", x"f1", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f3", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"ed", x"ef", 
        x"f5", x"f4", x"f1", x"f3", x"f3", x"f1", x"f0", x"f1", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f5", x"f7", x"f9", x"f9", x"f4", x"ec", x"e0", x"cd", x"bf", x"af", x"aa", x"ae", 
        x"ba", x"c4", x"cd", x"d4", x"db", x"e3", x"ea", x"ef", x"f0", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", 
        x"f1", x"f1", x"f1", x"ef", x"f0", x"f1", x"f3", x"f4", x"f4", x"f2", x"ef", x"f1", x"f3", x"f3", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f5", x"f5", x"f5", x"f4", x"f4", x"f5", x"f5", x"f6", x"f7", 
        x"f9", x"f8", x"f6", x"f5", x"f5", x"f5", x"f5", x"f4", x"f4", x"f5", x"f6", x"f5", x"f4", x"f2", x"f5", 
        x"f9", x"f7", x"f3", x"f2", x"f4", x"f4", x"f3", x"f1", x"ef", x"f2", x"f0", x"f0", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"f4", x"f8", x"f6", x"f4", x"f5", x"f7", 
        x"f4", x"e7", x"8d", x"4e", x"5e", x"b2", x"df", x"d6", x"d4", x"d6", x"d7", x"aa", x"9f", x"a9", x"c4", 
        x"d6", x"d6", x"ae", x"9a", x"9a", x"99", x"9a", x"9b", x"99", x"98", x"98", x"99", x"97", x"96", x"94", 
        x"92", x"92", x"92", x"95", x"92", x"93", x"7e", x"4c", x"4e", x"69", x"86", x"8e", x"97", x"97", x"90", 
        x"8e", x"93", x"8e", x"81", x"7e", x"75", x"6a", x"61", x"59", x"59", x"5e", x"5f", x"6f", x"7e", x"7f", 
        x"82", x"85", x"7a", x"87", x"de", x"dd", x"e2", x"e3", x"e2", x"e2", x"e3", x"e1", x"de", x"e0", x"e3", 
        x"e2", x"e0", x"e1", x"e0", x"e2", x"e2", x"df", x"e0", x"df", x"db", x"e0", x"e0", x"df", x"e0", x"e0", 
        x"e1", x"e4", x"e2", x"e3", x"e0", x"da", x"d2", x"c6", x"ba", x"a7", x"94", x"7f", x"6a", x"57", x"4f", 
        x"4c", x"54", x"55", x"5e", x"63", x"5a", x"5b", x"5c", x"51", x"4b", x"46", x"46", x"42", x"38", x"31", 
        x"22", x"10", x"08", x"06", x"04", x"07", x"0f", x"17", x"21", x"2d", x"36", x"41", x"4f", x"5d", x"6e", 
        x"80", x"8e", x"93", x"97", x"99", x"95", x"3c", x"27", x"6a", x"6f", x"6e", x"83", x"88", x"83", x"7f", 
        x"a5", x"a7", x"a6", x"a4", x"a5", x"a6", x"a4", x"a5", x"a6", x"a6", x"a6", x"a6", x"a5", x"a4", x"a4", 
        x"a3", x"a3", x"a4", x"a4", x"a4", x"a5", x"a4", x"a4", x"a5", x"a6", x"a6", x"a5", x"a4", x"a5", x"a6", 
        x"a3", x"a3", x"a5", x"a5", x"a5", x"a7", x"a6", x"a5", x"a5", x"a5", x"a5", x"a6", x"a7", x"a5", x"a5", 
        x"a5", x"a6", x"a6", x"a6", x"a7", x"a6", x"a6", x"a5", x"a6", x"a6", x"a6", x"a7", x"a7", x"a7", x"a6", 
        x"a6", x"a6", x"a6", x"a7", x"a8", x"a8", x"a7", x"a7", x"a7", x"a7", x"a5", x"a3", x"a5", x"a6", x"a6", 
        x"a7", x"a7", x"a6", x"a6", x"a9", x"a8", x"a7", x"a6", x"a6", x"a6", x"a7", x"a8", x"a9", x"a9", x"a8", 
        x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a9", x"a9", x"a9", x"a8", x"a7", x"a7", x"a8", 
        x"a3", x"c0", x"d6", x"d4", x"d1", x"d1", x"d5", x"d3", x"d4", x"d4", x"d3", x"d4", x"d9", x"db", x"d6", 
        x"c6", x"ac", x"7a", x"53", x"31", x"17", x"23", x"3b", x"28", x"1a", x"45", x"6f", x"7d", x"79", x"73", 
        x"73", x"78", x"67", x"59", x"4e", x"4b", x"49", x"46", x"44", x"42", x"44", x"43", x"43", x"45", x"46", 
        x"41", x"44", x"a3", x"e4", x"d5", x"d5", x"d6", x"d4", x"de", x"d6", x"ce", x"d1", x"d4", x"d4", x"d2", 
        x"d3", x"d2", x"d2", x"d2", x"d3", x"d4", x"d6", x"d4", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d2", 
        x"d1", x"d2", x"d2", x"d3", x"d4", x"d4", x"d3", x"d1", x"d3", x"d5", x"d5", x"d4", x"d4", x"d3", x"d3", 
        x"d6", x"d6", x"d5", x"d5", x"d5", x"d5", x"d6", x"d7", x"d8", x"d7", x"da", x"d6", x"d4", x"d7", x"d9", 
        x"d9", x"d7", x"d8", x"ec", x"f0", x"ec", x"ed", x"ef", x"ed", x"ef", x"ed", x"ee", x"f1", x"ef", x"ee", 
        x"ef", x"f0", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", 
        x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"f3", x"e7", x"b9", 
        x"bc", x"c7", x"d6", x"df", x"ea", x"f0", x"f3", x"f4", x"f5", x"f6", x"f5", x"f3", x"f1", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ee", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"ee", x"ef", x"f0", x"ef", x"ee", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f2", x"f2", 
        x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"ed", x"ee", 
        x"f4", x"f4", x"f1", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f4", x"f5", x"f5", x"f5", x"f4", x"f2", x"f1", x"f1", x"f0", x"ea", x"e2", 
        x"d7", x"cf", x"c6", x"c1", x"be", x"bc", x"bf", x"c3", x"c7", x"ce", x"d9", x"e6", x"f0", x"f3", x"f3", 
        x"f3", x"f4", x"f3", x"f1", x"f0", x"f1", x"f2", x"f4", x"f5", x"f4", x"f1", x"f2", x"f3", x"f2", x"f1", 
        x"f1", x"f0", x"f3", x"f4", x"f5", x"f5", x"f4", x"f4", x"f6", x"f4", x"f4", x"f4", x"f5", x"f6", x"f7", 
        x"f8", x"f7", x"f6", x"f5", x"f5", x"f4", x"f4", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f5", 
        x"f7", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ef", x"f2", x"f1", x"f0", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f1", x"f0", x"f3", x"f7", x"f6", x"f5", x"f5", x"f8", 
        x"f4", x"e9", x"92", x"4d", x"5b", x"ad", x"de", x"d5", x"d4", x"d6", x"d8", x"ac", x"9a", x"9b", x"9e", 
        x"a3", x"ab", x"a2", x"9d", x"9a", x"98", x"99", x"99", x"97", x"96", x"97", x"98", x"97", x"95", x"94", 
        x"92", x"93", x"93", x"94", x"91", x"93", x"81", x"4e", x"4e", x"66", x"85", x"8c", x"96", x"9a", x"96", 
        x"90", x"91", x"8a", x"7c", x"7d", x"7e", x"7b", x"77", x"71", x"70", x"6c", x"64", x"66", x"69", x"69", 
        x"70", x"75", x"70", x"7e", x"de", x"df", x"df", x"e3", x"e3", x"df", x"e0", x"e1", x"df", x"df", x"e0", 
        x"e1", x"e1", x"e2", x"e2", x"e1", x"e0", x"e0", x"e3", x"e5", x"e3", x"e6", x"e7", x"e7", x"e2", x"d8", 
        x"ca", x"bb", x"ad", x"9d", x"8d", x"80", x"76", x"6e", x"64", x"62", x"60", x"55", x"53", x"55", x"4d", 
        x"45", x"49", x"30", x"35", x"42", x"34", x"2e", x"2d", x"25", x"20", x"1a", x"13", x"0d", x"0c", x"0e", 
        x"0e", x"16", x"24", x"2f", x"38", x"48", x"59", x"64", x"70", x"7e", x"85", x"89", x"8e", x"90", x"8f", 
        x"8f", x"8d", x"8b", x"8b", x"8b", x"8a", x"40", x"22", x"69", x"72", x"70", x"82", x"83", x"82", x"7f", 
        x"a7", x"a7", x"a5", x"a4", x"a6", x"a7", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a5", x"a6", x"a5", 
        x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a5", x"a4", x"a5", x"a5", x"a5", x"a5", x"a4", x"a5", x"a7", 
        x"a4", x"a4", x"a5", x"a6", x"a6", x"a7", x"a6", x"a6", x"a5", x"a5", x"a5", x"a5", x"a4", x"a5", x"a5", 
        x"a5", x"a6", x"a6", x"a6", x"a7", x"a6", x"a6", x"a5", x"a6", x"a6", x"a6", x"a7", x"a8", x"a8", x"a7", 
        x"a6", x"a6", x"a7", x"a8", x"a8", x"a8", x"a7", x"a7", x"a8", x"a7", x"a6", x"a5", x"a7", x"a7", x"a7", 
        x"a7", x"a7", x"a6", x"a5", x"a8", x"a8", x"a7", x"a7", x"a7", x"a7", x"a8", x"a9", x"a9", x"a9", x"a9", 
        x"a9", x"a9", x"a9", x"a8", x"a8", x"a8", x"a8", x"a9", x"aa", x"aa", x"a8", x"aa", x"ac", x"a9", x"a7", 
        x"a4", x"c2", x"d8", x"d3", x"d5", x"d3", x"d1", x"d2", x"d4", x"d5", x"d8", x"d6", x"cf", x"b5", x"86", 
        x"5b", x"35", x"12", x"0e", x"15", x"14", x"26", x"48", x"40", x"24", x"47", x"66", x"72", x"76", x"74", 
        x"74", x"78", x"67", x"55", x"48", x"46", x"45", x"45", x"45", x"45", x"48", x"48", x"47", x"4a", x"4d", 
        x"47", x"45", x"a0", x"e2", x"d5", x"d6", x"d6", x"d4", x"e0", x"d7", x"cf", x"d0", x"d2", x"d4", x"d3", 
        x"d4", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d4", x"d3", x"d2", x"d2", x"d3", x"d3", x"d3", 
        x"d1", x"d2", x"d3", x"d3", x"d4", x"d4", x"d5", x"d3", x"d4", x"d5", x"d4", x"d3", x"d4", x"d3", x"d3", 
        x"d5", x"d6", x"d5", x"d6", x"d5", x"d5", x"d5", x"d4", x"d6", x"d7", x"dc", x"d7", x"d6", x"d6", x"d9", 
        x"dc", x"d6", x"d6", x"ec", x"f0", x"ec", x"ee", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ed", 
        x"ee", x"ef", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"eb", x"eb", x"ee", 
        x"ee", x"f0", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"ef", x"ef", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"f0", x"f3", x"dc", x"7e", 
        x"6a", x"7b", x"86", x"90", x"9e", x"a9", x"b2", x"be", x"cb", x"d5", x"de", x"e7", x"ed", x"f0", x"f1", 
        x"f1", x"f2", x"f1", x"ef", x"ef", x"f0", x"f1", x"ee", x"ee", x"f0", x"f2", x"f2", x"ef", x"ee", x"ed", 
        x"ef", x"ee", x"ec", x"ef", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"f0", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"ed", x"ee", 
        x"f4", x"f4", x"f2", x"f2", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f4", x"f5", x"f5", x"f3", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f5", 
        x"f6", x"f6", x"f3", x"ef", x"e7", x"dc", x"ce", x"c2", x"ba", x"b7", x"ba", x"be", x"c2", x"c6", x"ce", 
        x"d6", x"e0", x"e6", x"ec", x"f1", x"f2", x"f3", x"f3", x"f1", x"f0", x"ef", x"f2", x"f4", x"f2", x"f0", 
        x"f2", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f5", x"f4", x"f5", x"f6", x"f6", x"f6", x"f6", 
        x"f7", x"f7", x"f6", x"f6", x"f5", x"f4", x"f3", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f5", 
        x"f4", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"ef", x"ef", x"f2", x"f1", x"f1", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f1", x"ef", x"f1", x"f4", x"f0", x"f2", x"f6", x"f6", x"f5", x"f5", x"f6", 
        x"f4", x"ec", x"9a", x"4c", x"57", x"a7", x"dc", x"d5", x"d4", x"d6", x"d9", x"af", x"9c", x"a1", x"9b", 
        x"96", x"97", x"9a", x"9b", x"9b", x"98", x"98", x"98", x"97", x"96", x"97", x"97", x"96", x"95", x"94", 
        x"93", x"93", x"94", x"93", x"92", x"96", x"85", x"4f", x"4f", x"62", x"85", x"8d", x"92", x"96", x"96", 
        x"90", x"92", x"8e", x"7c", x"7a", x"7b", x"79", x"79", x"78", x"7a", x"7a", x"77", x"7a", x"7a", x"73", 
        x"71", x"6b", x"60", x"6c", x"d6", x"e1", x"df", x"e4", x"e4", x"e0", x"e0", x"e1", x"df", x"df", x"e0", 
        x"e2", x"e3", x"e3", x"e4", x"e3", x"e3", x"e3", x"e0", x"dc", x"d5", x"c8", x"ba", x"ab", x"9d", x"8c", 
        x"7c", x"6e", x"64", x"59", x"57", x"56", x"55", x"58", x"54", x"4d", x"45", x"35", x"29", x"20", x"15", 
        x"0f", x"19", x"0b", x"14", x"1e", x"15", x"0d", x"09", x"09", x"0d", x"13", x"1a", x"24", x"31", x"3e", 
        x"48", x"57", x"6a", x"78", x"82", x"8a", x"90", x"92", x"93", x"92", x"8e", x"8b", x"89", x"8a", x"89", 
        x"85", x"83", x"84", x"86", x"88", x"8a", x"48", x"1f", x"66", x"72", x"71", x"81", x"83", x"81", x"81", 
        x"a8", x"a7", x"a5", x"a4", x"a6", x"a7", x"a5", x"a6", x"a6", x"a6", x"a5", x"a5", x"a6", x"a7", x"a6", 
        x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a5", x"a5", x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", 
        x"a5", x"a4", x"a5", x"a7", x"a7", x"a6", x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a5", x"a5", x"a5", 
        x"a5", x"a6", x"a6", x"a6", x"a7", x"a6", x"a6", x"a5", x"a6", x"a6", x"a6", x"a7", x"a7", x"a7", x"a7", 
        x"a7", x"a7", x"a7", x"a7", x"a6", x"a6", x"a7", x"a8", x"a9", x"a9", x"a8", x"a9", x"a8", x"a8", x"a9", 
        x"a8", x"a7", x"a7", x"a6", x"a7", x"a7", x"a8", x"a8", x"a9", x"a9", x"aa", x"a9", x"a8", x"a8", x"a8", 
        x"a8", x"a8", x"a9", x"a9", x"a9", x"a9", x"a9", x"aa", x"ab", x"ab", x"a8", x"a8", x"a9", x"a7", x"a7", 
        x"a5", x"c1", x"d3", x"cf", x"d3", x"d2", x"d6", x"e1", x"e2", x"d6", x"b0", x"7f", x"55", x"2f", x"16", 
        x"10", x"0d", x"12", x"16", x"17", x"19", x"2d", x"48", x"4e", x"2d", x"48", x"65", x"75", x"76", x"71", 
        x"6e", x"6f", x"64", x"52", x"49", x"47", x"44", x"45", x"44", x"49", x"4c", x"4e", x"4d", x"4e", x"50", 
        x"4c", x"46", x"9d", x"e0", x"d4", x"d5", x"d5", x"d2", x"df", x"d8", x"d1", x"d2", x"d4", x"d4", x"d4", 
        x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", 
        x"d3", x"d4", x"d4", x"d3", x"d3", x"d4", x"d5", x"d4", x"d4", x"d4", x"d3", x"d2", x"d3", x"d2", x"d3", 
        x"d5", x"d6", x"d6", x"d7", x"d5", x"d4", x"d4", x"d3", x"d5", x"d7", x"dc", x"d5", x"d3", x"d3", x"d6", 
        x"d8", x"d4", x"d5", x"ec", x"ef", x"ed", x"ee", x"ef", x"ed", x"ec", x"ed", x"ef", x"f0", x"f0", x"ef", 
        x"ee", x"ee", x"ee", x"ed", x"ed", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"e8", x"e9", x"ee", 
        x"ef", x"f1", x"ee", x"ec", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f2", x"f1", x"f1", x"e1", x"69", 
        x"45", x"54", x"5c", x"67", x"71", x"75", x"79", x"7f", x"83", x"81", x"84", x"8a", x"92", x"9e", x"b0", 
        x"c0", x"d3", x"e3", x"ef", x"f4", x"f5", x"f7", x"f7", x"f2", x"f2", x"f4", x"f2", x"ee", x"ec", x"ed", 
        x"f0", x"f0", x"ee", x"ef", x"ee", x"ed", x"ee", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"ed", x"ed", 
        x"f3", x"f4", x"f2", x"f1", x"f3", x"f3", x"f3", x"f4", x"f3", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f4", x"f5", x"f6", x"f4", x"f3", x"f3", x"f4", x"f5", x"f5", x"f4", x"f3", x"f2", 
        x"f1", x"f2", x"f2", x"f3", x"f4", x"f4", x"f5", x"f4", x"f3", x"e9", x"e3", x"d9", x"d0", x"c7", x"be", 
        x"b8", x"b2", x"b2", x"b5", x"bb", x"c7", x"d8", x"e9", x"f3", x"f4", x"f4", x"f5", x"f5", x"f2", x"f0", 
        x"f1", x"f2", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f4", x"f5", x"f6", x"f7", x"f6", x"f6", x"f5", 
        x"f6", x"f7", x"f7", x"f6", x"f5", x"f4", x"f3", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f5", 
        x"f3", x"f0", x"f2", x"f3", x"f2", x"f0", x"f2", x"f0", x"ef", x"f2", x"f2", x"f1", x"f2", x"f1", x"f2", 
        x"f3", x"f5", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"f2", x"f6", x"f1", x"f1", x"f6", x"f7", x"f5", x"f5", x"f5", 
        x"f4", x"ee", x"a3", x"4c", x"55", x"a4", x"de", x"d7", x"d5", x"d3", x"d7", x"b2", x"9e", x"a2", x"9e", 
        x"a0", x"a1", x"a0", x"9a", x"9b", x"99", x"99", x"99", x"98", x"96", x"98", x"95", x"95", x"95", x"95", 
        x"94", x"94", x"92", x"93", x"92", x"96", x"88", x"53", x"52", x"61", x"86", x"89", x"8d", x"93", x"98", 
        x"91", x"93", x"91", x"7e", x"78", x"7b", x"79", x"79", x"78", x"77", x"76", x"78", x"81", x"87", x"87", 
        x"88", x"82", x"78", x"73", x"d2", x"e2", x"e0", x"e4", x"e1", x"e0", x"e1", x"e2", x"e4", x"e7", x"e9", 
        x"ea", x"e9", x"e4", x"dd", x"ca", x"b3", x"9b", x"89", x"7d", x"6f", x"6b", x"67", x"64", x"61", x"5e", 
        x"5a", x"55", x"53", x"4f", x"4b", x"42", x"37", x"34", x"2a", x"1d", x"13", x"09", x"04", x"04", x"02", 
        x"02", x"06", x"10", x"29", x"30", x"2d", x"2f", x"36", x"43", x"51", x"5e", x"6d", x"79", x"82", x"86", 
        x"87", x"8a", x"8c", x"8b", x"89", x"87", x"84", x"83", x"83", x"83", x"83", x"84", x"85", x"87", x"87", 
        x"84", x"84", x"85", x"85", x"88", x"8f", x"4e", x"1e", x"61", x"71", x"70", x"7a", x"82", x"81", x"7f", 
        x"a7", x"a7", x"a5", x"a4", x"a5", x"a6", x"a5", x"a6", x"a6", x"a6", x"a5", x"a5", x"a6", x"a7", x"a7", 
        x"a6", x"a6", x"a6", x"a6", x"a6", x"a6", x"a5", x"a5", x"a5", x"a4", x"a4", x"a5", x"a5", x"a6", x"a5", 
        x"a5", x"a4", x"a5", x"a7", x"a7", x"a5", x"a5", x"a6", x"a6", x"a7", x"a7", x"a6", x"a5", x"a5", x"a5", 
        x"a5", x"a6", x"a6", x"a6", x"a7", x"a6", x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", x"a6", x"a6", x"a7", 
        x"a8", x"a8", x"a7", x"a6", x"a6", x"a6", x"a7", x"a9", x"a9", x"a9", x"aa", x"aa", x"a8", x"a9", x"a9", 
        x"a9", x"a8", x"a8", x"a8", x"a9", x"a9", x"a9", x"a9", x"a9", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", 
        x"a8", x"a9", x"a9", x"a9", x"a9", x"a9", x"aa", x"aa", x"ab", x"ab", x"aa", x"a8", x"a9", x"aa", x"a7", 
        x"a2", x"c2", x"d6", x"d2", x"da", x"d9", x"ce", x"b3", x"85", x"5b", x"36", x"1b", x"11", x"0f", x"11", 
        x"17", x"1b", x"1c", x"1b", x"18", x"1b", x"31", x"49", x"4f", x"37", x"4f", x"60", x"6e", x"6f", x"6d", 
        x"6d", x"6d", x"63", x"53", x"4c", x"4d", x"49", x"4a", x"4a", x"4d", x"4e", x"51", x"51", x"4e", x"4f", 
        x"4e", x"4c", x"9f", x"e3", x"d5", x"d6", x"d5", x"d2", x"dd", x"d7", x"d2", x"d3", x"d5", x"d5", x"d4", 
        x"d3", x"d3", x"d4", x"d5", x"d5", x"d3", x"d2", x"d2", x"d3", x"d2", x"d2", x"d2", x"d2", x"d3", x"d2", 
        x"d2", x"d3", x"d5", x"d3", x"d4", x"d5", x"d6", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d3", 
        x"d5", x"d6", x"d6", x"d7", x"d5", x"d1", x"d4", x"d4", x"d5", x"d7", x"dd", x"d7", x"d4", x"d8", x"da", 
        x"dd", x"dd", x"d8", x"e5", x"eb", x"ed", x"ed", x"f0", x"f0", x"ee", x"ed", x"ef", x"ee", x"ef", x"ef", 
        x"ed", x"ec", x"ed", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ec", x"ec", x"ee", 
        x"ee", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f0", x"e1", x"5f", 
        x"1b", x"1b", x"20", x"26", x"2d", x"34", x"3f", x"4c", x"56", x"61", x"69", x"73", x"78", x"7a", x"7e", 
        x"80", x"82", x"89", x"92", x"9b", x"a7", x"b6", x"c0", x"d1", x"dd", x"e5", x"eb", x"ee", x"f0", x"f2", 
        x"f1", x"f1", x"f2", x"f1", x"ee", x"ee", x"ef", x"f0", x"f0", x"ee", x"ee", x"ee", x"ee", x"f0", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"ec", x"ed", 
        x"f3", x"f4", x"f3", x"f1", x"f3", x"f3", x"f4", x"f4", x"f3", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f3", 
        x"f3", x"f3", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f4", x"f3", x"f2", x"f3", x"f2", x"ec", 
        x"e5", x"dd", x"d6", x"ce", x"c3", x"bb", x"b7", x"b6", x"ba", x"be", x"c6", x"d7", x"e5", x"ec", x"ee", 
        x"f1", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f4", x"f5", x"f5", x"f5", x"f6", x"f6", x"f7", x"f7", 
        x"f7", x"f6", x"f6", x"f5", x"f5", x"f4", x"f3", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f1", x"f2", x"f3", x"f2", x"f1", x"f2", x"f0", x"ee", x"f1", x"f2", x"f2", x"f2", x"f1", x"f3", 
        x"f4", x"f5", x"f4", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"f3", x"f7", x"f1", x"f1", x"f7", x"f7", x"f5", x"f5", x"f5", 
        x"f5", x"f0", x"ab", x"4c", x"52", x"9d", x"dc", x"d6", x"d5", x"d3", x"d8", x"b6", x"9d", x"a1", x"9e", 
        x"a0", x"9d", x"9c", x"9a", x"9b", x"99", x"9a", x"9a", x"98", x"97", x"98", x"96", x"95", x"95", x"95", 
        x"95", x"93", x"92", x"92", x"92", x"92", x"87", x"50", x"4e", x"57", x"7f", x"85", x"8a", x"92", x"98", 
        x"91", x"92", x"92", x"81", x"77", x"7a", x"79", x"78", x"78", x"77", x"77", x"77", x"7d", x"83", x"85", 
        x"87", x"83", x"82", x"7b", x"cf", x"e5", x"e2", x"e5", x"e6", x"e5", x"e1", x"dd", x"d8", x"cc", x"b9", 
        x"a8", x"99", x"84", x"79", x"70", x"6e", x"6c", x"64", x"61", x"5a", x"59", x"57", x"51", x"4b", x"49", 
        x"49", x"45", x"3f", x"39", x"32", x"26", x"18", x"15", x"15", x"10", x"15", x"18", x"1e", x"28", x"2e", 
        x"17", x"07", x"1a", x"4a", x"54", x"46", x"49", x"5f", x"76", x"80", x"81", x"7d", x"7d", x"80", x"81", 
        x"84", x"85", x"87", x"8a", x"89", x"86", x"84", x"85", x"85", x"85", x"85", x"85", x"86", x"87", x"87", 
        x"86", x"86", x"86", x"84", x"86", x"8e", x"55", x"1e", x"60", x"76", x"74", x"78", x"81", x"81", x"7d", 
        x"a6", x"a7", x"a5", x"a2", x"a3", x"a5", x"a5", x"a7", x"a7", x"a6", x"a5", x"a5", x"a5", x"a6", x"a7", 
        x"a7", x"a7", x"a6", x"a6", x"a5", x"a5", x"a5", x"a6", x"a5", x"a4", x"a4", x"a5", x"a6", x"a6", x"a4", 
        x"a5", x"a4", x"a4", x"a6", x"a7", x"a5", x"a7", x"a8", x"a8", x"a7", x"a6", x"a5", x"a5", x"a5", x"a5", 
        x"a5", x"a6", x"a6", x"a6", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a8", x"a8", x"a7", x"a7", x"a7", 
        x"a8", x"a8", x"a7", x"a7", x"a6", x"a6", x"a8", x"a9", x"a8", x"a8", x"a8", x"a9", x"a8", x"a8", x"a9", 
        x"a9", x"a8", x"a8", x"a8", x"a8", x"a9", x"a9", x"a9", x"a8", x"a7", x"a6", x"a7", x"a7", x"a8", x"a8", 
        x"a9", x"a9", x"a9", x"a9", x"a9", x"a9", x"a9", x"aa", x"aa", x"aa", x"a9", x"a6", x"ab", x"ad", x"a6", 
        x"a3", x"c5", x"dc", x"da", x"c0", x"94", x"60", x"34", x"1d", x"17", x"11", x"0e", x"13", x"17", x"18", 
        x"19", x"19", x"18", x"19", x"18", x"1c", x"2f", x"45", x"4e", x"39", x"56", x"60", x"6a", x"70", x"6d", 
        x"6e", x"6b", x"5f", x"4d", x"47", x"4a", x"47", x"4d", x"4b", x"4c", x"4d", x"4f", x"4f", x"4f", x"52", 
        x"50", x"4d", x"9e", x"e4", x"d6", x"d6", x"d6", x"d4", x"db", x"d5", x"d0", x"d2", x"d4", x"d5", x"d5", 
        x"d4", x"d4", x"d5", x"d6", x"d5", x"d2", x"d0", x"d0", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", 
        x"d2", x"d4", x"d5", x"d3", x"d3", x"d5", x"d6", x"d3", x"d1", x"d2", x"d3", x"d3", x"d2", x"d1", x"d3", 
        x"d5", x"d6", x"d6", x"d7", x"d3", x"d0", x"d6", x"d7", x"d6", x"d6", x"dd", x"da", x"d7", x"e0", x"df", 
        x"d1", x"b8", x"a1", x"aa", x"ad", x"b2", x"ba", x"c5", x"d4", x"dc", x"e4", x"ec", x"ed", x"ef", x"f3", 
        x"f2", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", 
        x"ed", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"ef", x"f0", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"eb", x"ed", x"f2", x"e2", x"63", 
        x"13", x"0c", x"0c", x"09", x"06", x"05", x"08", x"0e", x"15", x"1c", x"20", x"27", x"32", x"40", x"50", 
        x"5d", x"6c", x"6f", x"73", x"79", x"7e", x"7d", x"7b", x"7b", x"81", x"88", x"94", x"a7", x"bc", x"ce", 
        x"db", x"e7", x"ef", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"ec", x"ed", 
        x"f3", x"f4", x"f3", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f3", x"f1", x"f0", x"f1", x"f4", x"f5", 
        x"f3", x"f3", x"f3", x"f2", x"ef", x"ea", x"e2", x"dc", x"d3", x"c7", x"bb", x"b5", x"b6", x"b8", x"ba", 
        x"c3", x"d3", x"df", x"ea", x"f2", x"f4", x"f4", x"f4", x"f4", x"f5", x"f6", x"f8", x"f7", x"f7", x"f6", 
        x"f7", x"f7", x"f5", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f1", x"ed", x"f0", x"f1", x"f2", x"f2", x"f1", x"f4", 
        x"f5", x"f6", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f4", x"f7", x"f1", x"f1", x"f7", x"f7", x"f5", x"f5", x"f6", 
        x"f6", x"f2", x"b1", x"4d", x"51", x"99", x"dc", x"d7", x"d5", x"d1", x"d7", x"b8", x"9b", x"9f", x"9e", 
        x"9f", x"9e", x"9b", x"99", x"9a", x"99", x"9a", x"9a", x"99", x"97", x"98", x"97", x"96", x"95", x"94", 
        x"93", x"93", x"92", x"91", x"90", x"91", x"89", x"54", x"52", x"56", x"80", x"87", x"8b", x"8e", x"94", 
        x"8f", x"91", x"96", x"88", x"7a", x"7b", x"78", x"77", x"79", x"78", x"77", x"75", x"7c", x"82", x"83", 
        x"86", x"81", x"7d", x"7c", x"ca", x"e8", x"e3", x"d9", x"ca", x"b2", x"9d", x"87", x"75", x"68", x"5f", 
        x"5f", x"66", x"63", x"62", x"62", x"5f", x"53", x"44", x"45", x"47", x"48", x"4a", x"44", x"38", x"2e", 
        x"29", x"1d", x"17", x"16", x"16", x"12", x"12", x"17", x"20", x"2b", x"3f", x"44", x"47", x"50", x"54", 
        x"2b", x"0a", x"17", x"4b", x"51", x"40", x"39", x"35", x"40", x"4f", x"58", x"5a", x"5f", x"64", x"66", 
        x"66", x"65", x"6a", x"75", x"80", x"89", x"8e", x"8c", x"8a", x"85", x"83", x"83", x"86", x"89", x"88", 
        x"86", x"87", x"88", x"86", x"84", x"8a", x"5c", x"1e", x"5c", x"79", x"73", x"77", x"7f", x"80", x"7d", 
        x"a6", x"a7", x"a6", x"a2", x"a3", x"a6", x"a6", x"a8", x"a8", x"a7", x"a6", x"a6", x"a5", x"a5", x"a6", 
        x"a7", x"a6", x"a5", x"a5", x"a5", x"a5", x"a5", x"a6", x"a5", x"a4", x"a4", x"a5", x"a6", x"a5", x"a4", 
        x"a5", x"a4", x"a4", x"a6", x"a6", x"a4", x"a5", x"a5", x"a7", x"a0", x"a0", x"a8", x"a9", x"a6", x"a5", 
        x"a6", x"a6", x"a6", x"a7", x"a7", x"a7", x"a8", x"a7", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a7", 
        x"a6", x"a6", x"a7", x"a8", x"a8", x"a8", x"a9", x"aa", x"a8", x"a7", x"a7", x"a8", x"a8", x"a8", x"a9", 
        x"a9", x"aa", x"a9", x"a9", x"a7", x"a8", x"a9", x"aa", x"a9", x"a9", x"a8", x"a8", x"a8", x"a8", x"a9", 
        x"a9", x"aa", x"aa", x"a9", x"a9", x"a9", x"a9", x"a9", x"aa", x"aa", x"aa", x"a8", x"aa", x"ab", x"a8", 
        x"a9", x"b5", x"a1", x"69", x"36", x"21", x"1c", x"1a", x"14", x"12", x"13", x"16", x"17", x"16", x"18", 
        x"1a", x"18", x"15", x"14", x"0d", x"15", x"2f", x"42", x"52", x"3d", x"5c", x"63", x"64", x"6d", x"6e", 
        x"71", x"72", x"69", x"58", x"52", x"53", x"50", x"54", x"51", x"53", x"53", x"51", x"4e", x"4e", x"4f", 
        x"4a", x"49", x"99", x"e1", x"d3", x"d5", x"d7", x"d6", x"db", x"d4", x"ce", x"d0", x"d2", x"d3", x"d4", 
        x"d1", x"d1", x"d3", x"d5", x"d6", x"d4", x"d3", x"d1", x"d1", x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", 
        x"d4", x"d5", x"d5", x"d3", x"d2", x"d3", x"d5", x"d2", x"d2", x"d3", x"d4", x"d5", x"d3", x"d2", x"d4", 
        x"d6", x"d6", x"d6", x"d7", x"d3", x"d0", x"d3", x"d4", x"d3", x"d4", x"de", x"d6", x"cd", x"b7", x"9b", 
        x"8d", x"9d", x"b9", x"d1", x"cf", x"c5", x"bc", x"b2", x"a8", x"9f", x"a2", x"a9", x"ae", x"b8", x"c3", 
        x"cd", x"d4", x"db", x"e3", x"e7", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", 
        x"ee", x"ef", x"ee", x"ef", x"ee", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"ee", x"f0", x"f3", x"e4", x"7a", 
        x"3f", x"45", x"39", x"2f", x"26", x"1d", x"13", x"0e", x"0e", x"0b", x"09", x"07", x"08", x"0b", x"0f", 
        x"13", x"19", x"1b", x"1e", x"25", x"32", x"48", x"5c", x"68", x"70", x"79", x"81", x"83", x"7f", x"7c", 
        x"79", x"82", x"91", x"9d", x"aa", x"bd", x"cc", x"da", x"e4", x"e7", x"ed", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f1", x"ef", x"ed", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f1", x"ec", x"ed", 
        x"f3", x"f4", x"f3", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f1", x"f2", x"f2", x"f3", x"f2", 
        x"f2", x"f1", x"f3", x"f4", x"f4", x"f4", x"f5", x"f4", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f0", x"f1", x"f3", x"f5", x"f5", x"f4", x"f0", x"ea", x"e8", x"e6", x"de", x"d1", 
        x"c5", x"b8", x"b4", x"b3", x"b6", x"c1", x"ce", x"d9", x"e2", x"e9", x"f0", x"f5", x"f6", x"f4", x"f3", 
        x"f8", x"f7", x"f5", x"f2", x"f2", x"f3", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f3", x"f1", x"f2", x"f1", x"ed", x"f0", x"f0", x"f2", x"f2", x"f2", x"f4", 
        x"f5", x"f5", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f4", x"f7", x"f0", x"f1", x"f8", x"f7", x"f5", x"f6", x"f7", 
        x"f6", x"f2", x"b5", x"4d", x"4f", x"94", x"da", x"d7", x"d6", x"d3", x"da", x"be", x"9e", x"a3", x"a1", 
        x"9f", x"9f", x"9c", x"99", x"99", x"98", x"99", x"9a", x"98", x"97", x"97", x"99", x"98", x"95", x"91", 
        x"91", x"92", x"93", x"93", x"92", x"93", x"8d", x"58", x"54", x"54", x"7f", x"89", x"8c", x"8d", x"91", 
        x"8d", x"8f", x"97", x"8d", x"7c", x"7a", x"77", x"77", x"79", x"78", x"76", x"73", x"79", x"7f", x"82", 
        x"85", x"84", x"84", x"77", x"96", x"8c", x"7a", x"6e", x"68", x"69", x"6b", x"6e", x"70", x"6f", x"6e", 
        x"70", x"72", x"62", x"48", x"39", x"32", x"2b", x"26", x"2b", x"27", x"1f", x"1a", x"15", x"12", x"14", 
        x"18", x"1a", x"23", x"30", x"37", x"3e", x"51", x"69", x"79", x"87", x"85", x"65", x"56", x"5c", x"5a", 
        x"2d", x"10", x"2d", x"61", x"5a", x"4d", x"3b", x"2b", x"2c", x"27", x"25", x"29", x"38", x"4b", x"58", 
        x"61", x"65", x"66", x"62", x"60", x"68", x"75", x"83", x"89", x"8d", x"8c", x"8a", x"88", x"87", x"86", 
        x"83", x"82", x"85", x"87", x"87", x"8b", x"67", x"1e", x"58", x"79", x"71", x"7a", x"80", x"80", x"7d", 
        x"a5", x"a6", x"a8", x"a4", x"a4", x"a8", x"a6", x"a7", x"a6", x"a4", x"a6", x"a7", x"a8", x"a6", x"a6", 
        x"a8", x"a6", x"a5", x"a7", x"a5", x"a5", x"a6", x"a5", x"a5", x"a5", x"a5", x"a6", x"a6", x"a6", x"a5", 
        x"a8", x"a3", x"a4", x"a5", x"a4", x"a6", x"a6", x"a5", x"aa", x"7d", x"74", x"a2", x"aa", x"a7", x"a7", 
        x"a8", x"a9", x"a9", x"a7", x"a6", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a7", 
        x"a7", x"a6", x"a7", x"a7", x"a7", x"a9", x"aa", x"aa", x"a9", x"a9", x"a8", x"a7", x"a9", x"a8", x"a9", 
        x"a9", x"a9", x"a9", x"aa", x"a9", x"a8", x"a8", x"a8", x"a9", x"a9", x"a9", x"a9", x"a9", x"aa", x"ab", 
        x"ab", x"aa", x"aa", x"a9", x"a9", x"a9", x"a9", x"aa", x"aa", x"aa", x"ab", x"aa", x"a6", x"a9", x"ae", 
        x"ab", x"a3", x"8a", x"41", x"1f", x"32", x"2f", x"1c", x"19", x"18", x"18", x"15", x"14", x"14", x"12", 
        x"11", x"14", x"12", x"0f", x"0a", x"10", x"33", x"44", x"54", x"49", x"5a", x"64", x"68", x"70", x"71", 
        x"72", x"71", x"6f", x"66", x"60", x"60", x"5d", x"5c", x"5e", x"60", x"65", x"69", x"6a", x"68", x"64", 
        x"5c", x"53", x"9e", x"e1", x"cf", x"d4", x"d6", x"d6", x"de", x"d6", x"ce", x"d0", x"d0", x"d0", x"d3", 
        x"d3", x"d2", x"d3", x"d4", x"d4", x"d3", x"d2", x"d0", x"d1", x"d2", x"d1", x"d5", x"d3", x"d3", x"d5", 
        x"d4", x"d3", x"d3", x"d3", x"d3", x"d4", x"d5", x"d4", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", 
        x"d5", x"d6", x"d6", x"d6", x"d4", x"d2", x"d2", x"d2", x"d3", x"d6", x"d6", x"a5", x"82", x"89", x"ae", 
        x"cd", x"d5", x"d7", x"e9", x"f0", x"ef", x"ef", x"ef", x"ec", x"e7", x"e0", x"d9", x"d4", x"c8", x"b7", 
        x"b2", x"a9", x"a3", x"a6", x"ac", x"bd", x"c4", x"c6", x"cd", x"d1", x"dc", x"e2", x"e3", x"eb", x"ec", 
        x"ed", x"ec", x"eb", x"ef", x"ef", x"ef", x"f0", x"ef", x"ed", x"ee", x"ef", x"ef", x"f0", x"f0", x"ee", 
        x"f0", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", 
        x"ee", x"f0", x"f0", x"ef", x"f1", x"f1", x"f1", x"f1", x"ee", x"ee", x"ef", x"ef", x"ef", x"f1", x"f2", 
        x"f1", x"ef", x"ee", x"ee", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"ee", x"ef", x"f1", x"e4", x"7b", 
        x"52", x"60", x"5e", x"5f", x"5c", x"56", x"53", x"50", x"49", x"3d", x"38", x"2e", x"26", x"1b", x"16", 
        x"10", x"0d", x"0e", x"12", x"11", x"0e", x"0f", x"10", x"0e", x"13", x"21", x"32", x"45", x"55", x"64", 
        x"6f", x"74", x"7d", x"81", x"7e", x"77", x"72", x"7a", x"84", x"8d", x"9f", x"b2", x"bf", x"cb", x"d5", 
        x"de", x"e4", x"e9", x"ed", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", 
        x"f1", x"f1", x"f2", x"f3", x"f1", x"f1", x"f4", x"f2", x"f1", x"f3", x"f3", x"f1", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"ef", x"f1", x"f2", x"f2", x"f2", x"f0", x"f1", x"f2", x"f3", x"f3", x"f2", x"f0", x"f2", 
        x"f3", x"f2", x"f1", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f2", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f0", x"ed", 
        x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f5", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f5", x"f5", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f0", x"ed", x"e7", x"dd", x"cd", x"be", x"b3", x"a8", x"b3", x"bf", x"cb", x"d6", x"de", x"e6", 
        x"ec", x"f0", x"f2", x"f0", x"f1", x"f2", x"f3", x"f1", x"f1", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", 
        x"f3", x"f1", x"f2", x"f3", x"f3", x"f2", x"f3", x"ef", x"ed", x"f1", x"f1", x"f2", x"f1", x"f0", x"f3", 
        x"f5", x"f4", x"f2", x"f2", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f6", x"f3", x"f1", x"f6", x"f6", x"f4", x"f6", x"f4", 
        x"f8", x"f3", x"bb", x"51", x"50", x"8e", x"d9", x"d5", x"d3", x"d6", x"d7", x"c0", x"a0", x"a5", x"a3", 
        x"9e", x"9d", x"9c", x"9c", x"9a", x"99", x"98", x"97", x"97", x"97", x"96", x"96", x"9d", x"99", x"91", 
        x"94", x"93", x"93", x"93", x"90", x"93", x"8d", x"59", x"53", x"53", x"7f", x"8a", x"8d", x"88", x"8d", 
        x"8d", x"8c", x"94", x"91", x"80", x"79", x"79", x"79", x"7a", x"7a", x"76", x"77", x"7b", x"83", x"83", 
        x"83", x"84", x"84", x"7f", x"77", x"72", x"74", x"75", x"76", x"71", x"73", x"75", x"6a", x"5f", x"59", 
        x"57", x"4f", x"44", x"2f", x"20", x"14", x"0a", x"0c", x"10", x"11", x"16", x"20", x"2d", x"3b", x"4a", 
        x"5a", x"6e", x"7d", x"87", x"8f", x"8c", x"81", x"81", x"81", x"87", x"80", x"5d", x"4d", x"50", x"53", 
        x"34", x"10", x"35", x"74", x"76", x"72", x"5b", x"46", x"42", x"37", x"2e", x"22", x"21", x"23", x"27", 
        x"30", x"3c", x"49", x"56", x"5f", x"62", x"5f", x"5e", x"6a", x"7e", x"89", x"8b", x"87", x"86", x"86", 
        x"88", x"83", x"86", x"87", x"85", x"8a", x"6e", x"1e", x"4e", x"74", x"6f", x"78", x"7f", x"82", x"7c", 
        x"a8", x"a7", x"a7", x"a2", x"a2", x"a7", x"a4", x"a5", x"a5", x"a5", x"a6", x"a8", x"a9", x"a7", x"a7", 
        x"a8", x"a8", x"a7", x"a8", x"a7", x"a7", x"a7", x"a5", x"a5", x"a6", x"a6", x"a6", x"a7", x"a6", x"a5", 
        x"a7", x"a5", x"a5", x"a7", x"a6", x"a7", x"a4", x"a7", x"a0", x"8d", x"80", x"9a", x"ac", x"aa", x"a7", 
        x"a7", x"a9", x"aa", x"a9", x"a8", x"a7", x"a8", x"a8", x"a8", x"a8", x"a9", x"a8", x"a7", x"a7", x"a7", 
        x"a7", x"a7", x"a7", x"a7", x"a7", x"a9", x"aa", x"a9", x"a9", x"a8", x"a8", x"a8", x"a8", x"a7", x"a8", 
        x"a8", x"a8", x"a8", x"a9", x"a9", x"a8", x"a8", x"a7", x"a8", x"a9", x"aa", x"a9", x"a9", x"a9", x"aa", 
        x"aa", x"aa", x"a9", x"a8", x"a8", x"a8", x"a9", x"a9", x"aa", x"ab", x"ac", x"ab", x"aa", x"a9", x"aa", 
        x"a9", x"ab", x"9c", x"5e", x"5f", x"7f", x"84", x"72", x"56", x"42", x"35", x"2d", x"27", x"22", x"1c", 
        x"19", x"19", x"14", x"11", x"0e", x"20", x"46", x"46", x"6a", x"6b", x"60", x"62", x"6e", x"73", x"71", 
        x"73", x"6d", x"68", x"61", x"60", x"62", x"5c", x"57", x"57", x"54", x"4f", x"4b", x"4b", x"51", x"58", 
        x"58", x"56", x"9f", x"e2", x"d2", x"d7", x"d8", x"d5", x"dd", x"d7", x"cf", x"d0", x"d0", x"d0", x"d1", 
        x"d2", x"d2", x"d3", x"d4", x"d4", x"d3", x"d2", x"cf", x"cf", x"d1", x"d2", x"d6", x"d5", x"d4", x"d5", 
        x"d4", x"d3", x"d3", x"d3", x"d4", x"d5", x"d5", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", 
        x"d5", x"d6", x"d6", x"d6", x"d4", x"d3", x"d3", x"d3", x"d5", x"d4", x"d4", x"c0", x"c0", x"cf", x"d7", 
        x"d4", x"ce", x"d4", x"e9", x"ee", x"eb", x"ec", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ec", x"e8", 
        x"ea", x"e6", x"e2", x"de", x"d7", x"d2", x"cc", x"bf", x"b6", x"ac", x"ae", x"af", x"b4", x"bd", x"c0", 
        x"c6", x"ca", x"ce", x"d5", x"da", x"e3", x"e5", x"e8", x"ee", x"ec", x"ed", x"ef", x"f2", x"f3", x"f2", 
        x"f3", x"f0", x"ef", x"f0", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", 
        x"ef", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"ee", x"ef", x"f0", x"f1", 
        x"f2", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"e3", x"7b", 
        x"52", x"5d", x"55", x"58", x"5a", x"5b", x"5c", x"5e", x"5f", x"61", x"60", x"5c", x"5a", x"53", x"4e", 
        x"41", x"33", x"2a", x"2e", x"27", x"1b", x"19", x"11", x"0e", x"1c", x"24", x"1f", x"19", x"1a", x"1b", 
        x"1b", x"1f", x"2e", x"3d", x"4b", x"55", x"5d", x"69", x"72", x"77", x"7b", x"7f", x"7f", x"7f", x"82", 
        x"87", x"95", x"a7", x"b4", x"be", x"c8", x"d2", x"da", x"e3", x"e8", x"ee", x"f4", x"f6", x"f1", x"f2", 
        x"f1", x"f2", x"f4", x"f4", x"f4", x"f5", x"f5", x"f3", x"f0", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f3", x"f4", 
        x"f4", x"f3", x"f3", x"f3", x"f2", x"f0", x"f2", x"f0", x"f0", x"f1", x"ee", x"ef", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ed", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f5", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f4", x"f4", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f2", x"f3", x"f3", x"f2", x"f0", x"ee", x"e5", x"df", x"d4", x"c8", x"be", x"ba", x"b9", 
        x"be", x"c5", x"cd", x"d5", x"db", x"e2", x"e8", x"ed", x"f1", x"f3", x"f5", x"f4", x"f3", x"f2", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f0", x"f2", x"f1", x"ee", x"f2", x"f2", x"f3", x"f2", x"f2", x"f4", 
        x"f5", x"f3", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f6", x"f3", x"f1", x"f5", x"f6", x"f5", x"f6", x"f5", 
        x"f8", x"f5", x"c0", x"54", x"53", x"8a", x"d7", x"d6", x"d3", x"d6", x"d7", x"c2", x"a0", x"a5", x"a3", 
        x"9e", x"9d", x"9c", x"9c", x"9b", x"99", x"98", x"97", x"96", x"96", x"96", x"94", x"9a", x"99", x"94", 
        x"95", x"94", x"94", x"94", x"90", x"94", x"90", x"5c", x"52", x"50", x"7c", x"87", x"8a", x"89", x"8d", 
        x"8b", x"8a", x"92", x"90", x"86", x"7e", x"7a", x"76", x"75", x"76", x"76", x"75", x"78", x"82", x"84", 
        x"85", x"85", x"85", x"85", x"82", x"85", x"87", x"83", x"7b", x"4f", x"30", x"29", x"28", x"1c", x"1e", 
        x"26", x"24", x"1e", x"18", x"1c", x"25", x"2f", x"39", x"43", x"50", x"5e", x"6d", x"7b", x"85", x"8c", 
        x"8d", x"8c", x"8e", x"89", x"89", x"89", x"83", x"87", x"88", x"85", x"7b", x"69", x"66", x"67", x"66", 
        x"42", x"13", x"2f", x"6f", x"7b", x"79", x"69", x"58", x"55", x"4f", x"4b", x"3e", x"35", x"2e", x"2a", 
        x"29", x"28", x"25", x"27", x"34", x"41", x"4d", x"5b", x"5b", x"60", x"6a", x"74", x"7d", x"83", x"82", 
        x"86", x"84", x"86", x"86", x"82", x"87", x"74", x"1c", x"4c", x"79", x"6b", x"74", x"7f", x"81", x"7c", 
        x"aa", x"a8", x"a7", x"9f", x"9e", x"a6", x"a2", x"a4", x"a6", x"a6", x"a7", x"a8", x"a8", x"a8", x"a6", 
        x"a4", x"a6", x"a7", x"a5", x"a6", x"a6", x"a5", x"a4", x"a5", x"a5", x"a5", x"a5", x"a6", x"a5", x"a5", 
        x"a8", x"a7", x"a7", x"a8", x"a9", x"a8", x"a6", x"a7", x"90", x"8b", x"a0", x"ac", x"ab", x"a7", x"a4", 
        x"a4", x"a7", x"a7", x"a6", x"a8", x"a7", x"a7", x"a8", x"a8", x"a8", x"a8", x"a9", x"a8", x"a6", x"a6", 
        x"a6", x"a7", x"a7", x"a7", x"a8", x"a9", x"a9", x"a8", x"a8", x"a8", x"a9", x"a9", x"a7", x"a7", x"a7", 
        x"a8", x"a8", x"a8", x"a9", x"a9", x"a8", x"a7", x"a7", x"a8", x"aa", x"ab", x"aa", x"a8", x"a8", x"a9", 
        x"aa", x"aa", x"a8", x"a8", x"a8", x"a8", x"a9", x"aa", x"ab", x"ab", x"aa", x"a9", x"ab", x"aa", x"aa", 
        x"aa", x"ae", x"a1", x"6c", x"85", x"a6", x"bb", x"c9", x"be", x"b6", x"ad", x"a1", x"94", x"86", x"78", 
        x"6c", x"64", x"57", x"51", x"54", x"68", x"79", x"52", x"71", x"69", x"60", x"6d", x"75", x"74", x"6f", 
        x"74", x"75", x"75", x"74", x"72", x"71", x"70", x"71", x"73", x"70", x"6f", x"6e", x"6b", x"69", x"67", 
        x"60", x"56", x"9a", x"de", x"d1", x"d6", x"d6", x"d1", x"db", x"d8", x"d0", x"d0", x"d1", x"d2", x"d0", 
        x"d2", x"d3", x"d3", x"d4", x"d3", x"d3", x"d1", x"d0", x"d0", x"d1", x"d3", x"d5", x"d4", x"d3", x"d3", 
        x"d3", x"d4", x"d5", x"d5", x"d5", x"d5", x"d4", x"d4", x"d5", x"d5", x"d5", x"d5", x"d5", x"d4", x"d4", 
        x"d5", x"d6", x"d6", x"d6", x"d4", x"d3", x"d1", x"d2", x"d5", x"d4", x"da", x"d5", x"d4", x"d5", x"d4", 
        x"d0", x"cd", x"d3", x"e9", x"f1", x"ed", x"ec", x"ec", x"ec", x"ee", x"ee", x"ef", x"ef", x"ee", x"ed", 
        x"e9", x"e9", x"ee", x"f0", x"ef", x"f0", x"f2", x"f0", x"f1", x"ea", x"e8", x"e2", x"d5", x"cf", x"c4", 
        x"bb", x"b2", x"ad", x"ac", x"ab", x"b7", x"b8", x"bd", x"cb", x"cb", x"d0", x"d5", x"d9", x"df", x"e6", 
        x"ec", x"ee", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ee", x"ed", x"ee", 
        x"ef", x"f1", x"f3", x"ef", x"f0", x"f2", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"f1", 
        x"f2", x"f3", x"f1", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f2", x"e6", x"7f", 
        x"52", x"5f", x"5b", x"5b", x"5c", x"5c", x"5b", x"5c", x"5d", x"5d", x"5c", x"5b", x"5b", x"5c", x"66", 
        x"5c", x"4f", x"45", x"47", x"45", x"3f", x"3a", x"32", x"46", x"55", x"52", x"44", x"3b", x"38", x"32", 
        x"2f", x"2e", x"29", x"1c", x"0f", x"09", x"08", x"14", x"25", x"33", x"41", x"4f", x"59", x"65", x"6c", 
        x"6f", x"78", x"7a", x"77", x"77", x"7d", x"81", x"8b", x"9e", x"ac", x"b5", x"c2", x"cd", x"d0", x"dc", 
        x"e3", x"eb", x"f1", x"f2", x"f1", x"f4", x"f5", x"f4", x"f4", x"f4", x"f3", x"f2", x"f4", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f0", x"f0", x"f1", x"f2", x"f4", x"f4", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f3", x"f3", x"f2", x"f2", x"f0", x"f0", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ed", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f3", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f1", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f2", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f5", x"f6", x"f6", x"f6", x"f4", x"f0", x"ea", 
        x"da", x"cc", x"bd", x"b1", x"af", x"b6", x"c3", x"d1", x"d7", x"d9", x"df", x"e6", x"ee", x"f2", x"f2", 
        x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f3", x"f3", x"ef", x"f3", x"f2", x"f2", x"f1", x"f1", x"f4", 
        x"f6", x"f4", x"f3", x"f3", x"f3", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f5", x"f3", x"f1", x"f5", x"f7", x"f5", x"f5", x"f6", 
        x"f6", x"f5", x"c5", x"58", x"57", x"85", x"d5", x"d7", x"d4", x"d5", x"d8", x"c6", x"a0", x"a5", x"a3", 
        x"9e", x"9c", x"9b", x"9a", x"9a", x"99", x"98", x"97", x"96", x"96", x"95", x"94", x"97", x"99", x"98", 
        x"95", x"93", x"93", x"94", x"90", x"93", x"92", x"60", x"51", x"52", x"7b", x"87", x"8a", x"8b", x"8e", 
        x"89", x"88", x"8f", x"90", x"8a", x"81", x"79", x"76", x"78", x"7a", x"7a", x"7a", x"7e", x"88", x"8a", 
        x"8a", x"89", x"83", x"7b", x"6f", x"62", x"56", x"47", x"3d", x"31", x"17", x"13", x"3c", x"43", x"52", 
        x"64", x"66", x"5f", x"57", x"5d", x"6c", x"7b", x"87", x"8f", x"93", x"95", x"93", x"91", x"91", x"91", 
        x"8e", x"8f", x"90", x"8a", x"8a", x"87", x"80", x"80", x"82", x"82", x"7b", x"75", x"79", x"7a", x"7e", 
        x"58", x"19", x"2c", x"6f", x"81", x"78", x"69", x"5b", x"5c", x"5a", x"5c", x"52", x"47", x"3c", x"31", 
        x"2f", x"39", x"38", x"2e", x"29", x"25", x"25", x"34", x"3c", x"48", x"54", x"59", x"5a", x"5c", x"63", 
        x"70", x"79", x"80", x"83", x"82", x"89", x"7a", x"1e", x"46", x"78", x"6d", x"78", x"80", x"7d", x"7c", 
        x"a7", x"a8", x"a7", x"9f", x"9a", x"a4", x"a3", x"a5", x"a7", x"a7", x"a7", x"a7", x"a7", x"a7", x"a6", 
        x"a4", x"a6", x"a8", x"a5", x"a7", x"a7", x"a5", x"a5", x"a6", x"a6", x"a6", x"a6", x"a7", x"a6", x"a5", 
        x"a6", x"a7", x"a6", x"a6", x"a6", x"a7", x"a6", x"a9", x"9f", x"85", x"95", x"98", x"9f", x"a6", x"a7", 
        x"a9", x"ab", x"a9", x"a5", x"a6", x"a5", x"a7", x"a8", x"a8", x"a8", x"a8", x"aa", x"a8", x"a6", x"a6", 
        x"a6", x"a6", x"a7", x"a7", x"a8", x"a9", x"a8", x"a8", x"a8", x"a8", x"a9", x"a9", x"a8", x"a8", x"a8", 
        x"a8", x"a9", x"a9", x"a9", x"a7", x"a7", x"a8", x"a8", x"a9", x"aa", x"aa", x"aa", x"a8", x"a7", x"a8", 
        x"aa", x"aa", x"a8", x"a8", x"a9", x"aa", x"a9", x"aa", x"aa", x"aa", x"ab", x"aa", x"a8", x"a8", x"a9", 
        x"a9", x"aa", x"9b", x"67", x"84", x"9f", x"ad", x"b7", x"bd", x"c1", x"c4", x"c7", x"c9", x"c9", x"c8", 
        x"c6", x"c5", x"c1", x"bd", x"b8", x"a3", x"91", x"54", x"75", x"79", x"84", x"85", x"6f", x"74", x"76", 
        x"74", x"77", x"78", x"74", x"73", x"76", x"74", x"72", x"74", x"73", x"73", x"74", x"75", x"75", x"75", 
        x"71", x"69", x"a3", x"e1", x"d1", x"d4", x"d4", x"d1", x"db", x"d9", x"d0", x"ce", x"d0", x"d3", x"d1", 
        x"d2", x"d3", x"d3", x"d3", x"d3", x"d2", x"d1", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", 
        x"d3", x"d3", x"d5", x"d5", x"d5", x"d4", x"d4", x"d3", x"d4", x"d4", x"d5", x"d4", x"d4", x"d3", x"d4", 
        x"d5", x"d6", x"d6", x"d5", x"d3", x"d2", x"d0", x"cf", x"d4", x"d5", x"d7", x"d2", x"d2", x"d3", x"d3", 
        x"d3", x"d1", x"d5", x"ea", x"f1", x"ec", x"ec", x"ee", x"f0", x"f0", x"ef", x"ed", x"eb", x"ef", x"f1", 
        x"ee", x"ef", x"f0", x"ed", x"ee", x"f0", x"ee", x"eb", x"ec", x"ed", x"f1", x"f1", x"f0", x"f1", x"f1", 
        x"f2", x"ef", x"eb", x"e7", x"dc", x"da", x"d0", x"c6", x"c3", x"b9", x"b5", x"b3", x"b2", x"b4", x"b6", 
        x"bb", x"bc", x"bc", x"c1", x"c8", x"d2", x"dd", x"e5", x"ea", x"ee", x"f0", x"f4", x"f4", x"f1", x"f1", 
        x"ef", x"ed", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f2", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"e6", x"81", 
        x"50", x"5f", x"5f", x"5d", x"5d", x"5d", x"5b", x"5c", x"5f", x"5d", x"5d", x"5d", x"5e", x"5f", x"65", 
        x"59", x"47", x"44", x"46", x"43", x"44", x"44", x"50", x"7d", x"76", x"5d", x"52", x"51", x"52", x"53", 
        x"58", x"5d", x"5c", x"4c", x"33", x"29", x"35", x"4d", x"56", x"48", x"3d", x"3a", x"33", x"28", x"22", 
        x"22", x"2e", x"3c", x"47", x"50", x"59", x"60", x"67", x"71", x"77", x"79", x"7c", x"7f", x"82", x"91", 
        x"99", x"a2", x"ad", x"b7", x"c2", x"cd", x"d7", x"e1", x"ec", x"f5", x"f6", x"f5", x"f5", x"f2", x"f0", 
        x"f1", x"f0", x"f1", x"f0", x"f1", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", 
        x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ed", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f5", x"f4", 
        x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f4", x"f2", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f4", x"f5", x"f4", x"f5", x"f6", x"f7", x"f7", x"f6", x"f5", x"f3", x"f5", x"f8", x"fa", x"f9", x"f6", 
        x"f5", x"f5", x"f6", x"f3", x"e8", x"dd", x"d6", x"cb", x"c4", x"bd", x"b9", x"bb", x"bf", x"c3", x"ca", 
        x"d3", x"de", x"e8", x"ef", x"f3", x"f5", x"f4", x"f3", x"ee", x"f2", x"f1", x"f1", x"f1", x"f3", x"f6", 
        x"f6", x"f3", x"f1", x"f3", x"f3", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f5", x"f3", x"f1", x"f5", x"f7", x"f6", x"f5", x"f7", 
        x"f4", x"f6", x"cb", x"5c", x"58", x"81", x"d3", x"d9", x"d4", x"d4", x"d8", x"c8", x"a0", x"a5", x"a3", 
        x"9e", x"9c", x"9a", x"99", x"9a", x"99", x"97", x"96", x"96", x"96", x"95", x"95", x"95", x"97", x"99", 
        x"95", x"92", x"93", x"93", x"90", x"92", x"94", x"64", x"4e", x"4e", x"77", x"87", x"8a", x"8b", x"8b", 
        x"8a", x"8b", x"8e", x"8c", x"90", x"8a", x"81", x"7c", x"7c", x"7e", x"7e", x"7b", x"75", x"6d", x"5b", 
        x"4d", x"44", x"3a", x"34", x"2f", x"2b", x"34", x"40", x"55", x"47", x"1e", x"22", x"76", x"86", x"89", 
        x"8a", x"8b", x"87", x"84", x"87", x"8c", x"8f", x"91", x"92", x"92", x"8f", x"8c", x"8b", x"8c", x"8e", 
        x"8e", x"90", x"8f", x"8c", x"8e", x"90", x"8e", x"8e", x"8a", x"8a", x"84", x"81", x"82", x"81", x"8a", 
        x"6e", x"1a", x"28", x"6c", x"7d", x"78", x"70", x"65", x"64", x"60", x"60", x"5a", x"51", x"48", x"3c", 
        x"35", x"3d", x"3d", x"37", x"37", x"37", x"35", x"30", x"2e", x"2c", x"2b", x"2c", x"33", x"3c", x"44", 
        x"4c", x"4f", x"56", x"61", x"6e", x"7c", x"76", x"21", x"3a", x"72", x"78", x"7b", x"7a", x"7a", x"7c", 
        x"a5", x"a8", x"a6", x"9f", x"99", x"a1", x"a5", x"a7", x"a7", x"a7", x"a7", x"a6", x"a6", x"a5", x"a6", 
        x"a5", x"a7", x"a8", x"a7", x"a8", x"a9", x"a6", x"a6", x"a6", x"a7", x"a7", x"a7", x"a7", x"a7", x"a5", 
        x"a5", x"a6", x"a5", x"a3", x"a4", x"a6", x"a7", x"aa", x"a8", x"94", x"80", x"7b", x"8c", x"a8", x"aa", 
        x"a8", x"a9", x"a9", x"a8", x"a7", x"a6", x"a7", x"a8", x"a8", x"a8", x"a8", x"a9", x"a8", x"a6", x"a6", 
        x"a7", x"a7", x"a7", x"a8", x"a8", x"a9", x"a8", x"a8", x"a8", x"a9", x"aa", x"a9", x"a9", x"a9", x"a9", 
        x"a9", x"aa", x"aa", x"aa", x"a6", x"a7", x"a8", x"aa", x"aa", x"a9", x"a9", x"aa", x"a8", x"a7", x"a8", 
        x"aa", x"aa", x"a9", x"aa", x"ab", x"aa", x"aa", x"a9", x"a8", x"a8", x"aa", x"ac", x"aa", x"a8", x"a8", 
        x"a8", x"ab", x"9e", x"6d", x"84", x"a1", x"a7", x"9e", x"a1", x"a2", x"a6", x"ac", x"b1", x"b3", x"b6", 
        x"b8", x"ba", x"bd", x"c3", x"ba", x"99", x"92", x"58", x"70", x"7b", x"83", x"86", x"74", x"78", x"7a", 
        x"76", x"78", x"7a", x"78", x"7a", x"7a", x"75", x"76", x"7a", x"79", x"79", x"78", x"78", x"78", x"77", 
        x"74", x"6d", x"a2", x"e2", x"d6", x"d6", x"d6", x"d3", x"dd", x"d9", x"cf", x"ce", x"d0", x"d3", x"d1", 
        x"d0", x"d0", x"d2", x"d2", x"d3", x"d4", x"d4", x"d5", x"d2", x"d0", x"d0", x"d0", x"d2", x"d3", x"d1", 
        x"d2", x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d3", x"d4", x"d5", x"d6", x"d5", x"d4", x"d3", x"d3", 
        x"d4", x"d5", x"d5", x"d4", x"d3", x"d3", x"d7", x"d1", x"d2", x"d6", x"d8", x"d3", x"d3", x"d4", x"d4", 
        x"d2", x"ce", x"d0", x"ea", x"f3", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ed", x"ef", x"f1", 
        x"ee", x"ef", x"ef", x"ec", x"ee", x"ef", x"ee", x"ed", x"ec", x"ed", x"ee", x"ef", x"ed", x"ec", x"ec", 
        x"ef", x"ee", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ec", x"e9", x"e3", x"df", x"d7", x"cd", 
        x"c7", x"c0", x"ba", x"b7", x"b3", x"b7", x"b9", x"b9", x"ba", x"bc", x"bf", x"c7", x"d0", x"d6", x"e1", 
        x"e7", x"e9", x"ef", x"f1", x"f2", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"ee", x"e7", x"87", 
        x"53", x"63", x"5e", x"5d", x"5d", x"5e", x"5f", x"5f", x"61", x"61", x"61", x"5e", x"5e", x"63", x"61", 
        x"59", x"4a", x"47", x"4e", x"49", x"44", x"45", x"51", x"65", x"5f", x"56", x"59", x"60", x"61", x"62", 
        x"62", x"62", x"62", x"65", x"64", x"65", x"70", x"7a", x"7c", x"7a", x"7d", x"7f", x"71", x"57", x"41", 
        x"2d", x"22", x"1d", x"19", x"12", x"11", x"18", x"26", x"32", x"3f", x"46", x"4c", x"56", x"61", x"6a", 
        x"70", x"76", x"7b", x"7f", x"85", x"8d", x"91", x"97", x"a2", x"ad", x"b7", x"c3", x"d1", x"da", x"e6", 
        x"ed", x"ef", x"f2", x"f2", x"f3", x"f5", x"f3", x"f3", x"f3", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f2", x"f3", x"f2", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ed", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f4", x"f3", x"f3", x"f2", x"f3", x"f3", x"f4", x"f4", x"f3", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f3", x"f4", x"f2", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f4", x"f6", x"f6", x"f6", x"f6", x"f3", x"f4", x"f8", x"fa", x"f7", x"f3", 
        x"f4", x"f3", x"f4", x"f4", x"f3", x"f2", x"f3", x"f2", x"ef", x"e9", x"e1", x"d7", x"cd", x"c4", x"c0", 
        x"be", x"be", x"bf", x"c3", x"cb", x"d1", x"db", x"e7", x"e7", x"f0", x"f3", x"f3", x"f2", x"f3", x"f2", 
        x"f3", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f5", x"f3", x"f1", x"f5", x"f7", x"f7", x"f7", x"f6", 
        x"f3", x"f6", x"cf", x"61", x"56", x"7d", x"d0", x"da", x"d4", x"d3", x"d8", x"ca", x"a1", x"a5", x"a3", 
        x"9e", x"9c", x"99", x"99", x"99", x"98", x"97", x"96", x"96", x"96", x"95", x"94", x"93", x"94", x"97", 
        x"97", x"94", x"94", x"94", x"92", x"91", x"96", x"69", x"4d", x"4f", x"75", x"87", x"8b", x"8a", x"8b", 
        x"8e", x"8f", x"90", x"90", x"90", x"87", x"77", x"68", x"5d", x"54", x"48", x"40", x"37", x"32", x"2f", 
        x"35", x"3f", x"4b", x"56", x"66", x"70", x"78", x"7d", x"8d", x"62", x"21", x"1f", x"7b", x"87", x"7f", 
        x"7b", x"7b", x"7c", x"7a", x"7a", x"7a", x"7a", x"7c", x"7f", x"83", x"84", x"88", x"8c", x"8b", x"8b", 
        x"8d", x"8d", x"8d", x"8a", x"8b", x"8a", x"86", x"86", x"89", x"88", x"82", x"83", x"85", x"84", x"8c", 
        x"77", x"20", x"3e", x"84", x"8b", x"7d", x"73", x"64", x"64", x"60", x"61", x"5f", x"55", x"49", x"40", 
        x"3b", x"41", x"43", x"41", x"40", x"3e", x"3b", x"3a", x"37", x"34", x"30", x"2a", x"24", x"22", x"22", 
        x"27", x"2b", x"2e", x"34", x"3b", x"40", x"45", x"23", x"3c", x"5b", x"6c", x"78", x"7c", x"7c", x"7d", 
        x"a6", x"a8", x"a2", x"a0", x"9a", x"9e", x"a6", x"a7", x"a7", x"a6", x"a6", x"a7", x"a8", x"a6", x"a4", 
        x"a4", x"a4", x"a5", x"a6", x"a6", x"a7", x"a6", x"a5", x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", x"a6", 
        x"a4", x"a6", x"a3", x"a2", x"a6", x"a7", x"ab", x"aa", x"ab", x"a1", x"7a", x"70", x"7b", x"a7", x"ae", 
        x"a8", x"a5", x"a7", x"a9", x"a7", x"a7", x"a8", x"a8", x"a8", x"a8", x"a9", x"a8", x"a8", x"a8", x"a8", 
        x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a8", x"a9", x"a9", x"aa", x"a9", x"a8", x"a9", x"a9", 
        x"a9", x"a9", x"aa", x"a9", x"a7", x"a7", x"a9", x"aa", x"aa", x"a9", x"a8", x"aa", x"a9", x"a8", x"a8", 
        x"a9", x"aa", x"aa", x"aa", x"ab", x"aa", x"aa", x"a9", x"a8", x"a8", x"a9", x"aa", x"ad", x"ad", x"ac", 
        x"a9", x"ad", x"a0", x"6c", x"83", x"a5", x"ac", x"a5", x"a2", x"9d", x"9d", x"9e", x"9d", x"9b", x"9c", 
        x"9c", x"9b", x"9c", x"9e", x"8d", x"6c", x"7c", x"55", x"6a", x"75", x"6c", x"77", x"78", x"76", x"78", 
        x"76", x"78", x"7d", x"78", x"75", x"78", x"79", x"78", x"79", x"79", x"7a", x"7a", x"7b", x"7a", x"7a", 
        x"76", x"6e", x"a1", x"e2", x"d6", x"d6", x"d5", x"d3", x"de", x"d7", x"ce", x"cf", x"d0", x"d1", x"d2", 
        x"cf", x"cf", x"d1", x"d2", x"d4", x"d6", x"d6", x"d5", x"d0", x"ce", x"d0", x"d0", x"d3", x"d4", x"d2", 
        x"d2", x"d2", x"d2", x"d3", x"d3", x"d4", x"d3", x"d2", x"d3", x"d4", x"d5", x"d4", x"d3", x"d2", x"d3", 
        x"d4", x"d5", x"d5", x"d4", x"d3", x"d2", x"d5", x"d1", x"d1", x"d3", x"d6", x"d2", x"d1", x"d1", x"d2", 
        x"d0", x"cd", x"cf", x"e9", x"f3", x"ee", x"ef", x"ee", x"ec", x"ec", x"ed", x"ef", x"ef", x"ef", x"f0", 
        x"ec", x"ed", x"ee", x"ef", x"f1", x"ed", x"ed", x"ed", x"eb", x"eb", x"ed", x"ee", x"ef", x"ee", x"ef", 
        x"f0", x"ed", x"ef", x"ee", x"ed", x"ea", x"ec", x"ef", x"ee", x"f0", x"ee", x"ee", x"f1", x"f1", x"f1", 
        x"f4", x"f2", x"ee", x"ea", x"e3", x"df", x"d8", x"ce", x"c5", x"c1", x"bd", x"b4", x"b3", x"ac", x"ad", 
        x"b0", x"b1", x"ba", x"c0", x"c9", x"ce", x"dc", x"e8", x"eb", x"f3", x"f4", x"f4", x"f5", x"f4", x"f3", 
        x"f2", x"f3", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"e9", x"8f", 
        x"5a", x"6c", x"6a", x"67", x"63", x"60", x"5e", x"5b", x"57", x"52", x"57", x"54", x"58", x"60", x"51", 
        x"52", x"52", x"4a", x"50", x"4b", x"47", x"49", x"51", x"57", x"5b", x"62", x"69", x"6c", x"6c", x"6d", 
        x"6f", x"6e", x"6b", x"6f", x"75", x"77", x"78", x"77", x"7e", x"83", x"78", x"5f", x"3f", x"2c", x"27", 
        x"24", x"21", x"22", x"1e", x"14", x"0b", x"09", x"06", x"05", x"07", x"0c", x"13", x"1a", x"1f", x"28", 
        x"2f", x"38", x"41", x"47", x"51", x"60", x"6b", x"74", x"7e", x"85", x"88", x"8b", x"8d", x"8f", x"98", 
        x"a2", x"ab", x"ba", x"ca", x"d9", x"e8", x"f1", x"f5", x"f7", x"f8", x"f6", x"f4", x"f2", x"ee", x"f0", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"ef", x"f1", x"f2", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ed", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f4", x"f3", x"f3", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f1", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f1", x"f2", x"f4", x"f7", x"f9", x"f8", x"f7", x"f5", x"f3", x"f3", x"f7", x"f8", x"f5", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f3", x"f5", x"f7", x"f6", x"f3", x"f1", x"ec", 
        x"e6", x"de", x"d5", x"cc", x"c4", x"be", x"bd", x"c3", x"bd", x"c2", x"ca", x"d5", x"df", x"ea", x"f1", 
        x"f4", x"f5", x"f4", x"f3", x"f1", x"ee", x"f3", x"f3", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f5", x"f3", x"f0", x"f5", x"f6", x"f6", x"f7", x"f5", 
        x"f3", x"f7", x"d5", x"69", x"53", x"78", x"cd", x"db", x"d4", x"d5", x"d8", x"cd", x"a3", x"a6", x"a3", 
        x"9d", x"9c", x"9a", x"9a", x"99", x"98", x"97", x"96", x"95", x"95", x"95", x"93", x"93", x"92", x"96", 
        x"9a", x"96", x"93", x"94", x"90", x"8d", x"93", x"69", x"4b", x"53", x"79", x"8f", x"97", x"98", x"95", 
        x"8b", x"7d", x"6f", x"5e", x"4f", x"3e", x"31", x"2e", x"30", x"33", x"3c", x"43", x"50", x"62", x"6e", 
        x"79", x"82", x"86", x"86", x"89", x"84", x"81", x"7e", x"87", x"62", x"23", x"1c", x"77", x"85", x"7d", 
        x"7e", x"7c", x"7a", x"7c", x"7d", x"7c", x"7c", x"7c", x"7c", x"7a", x"7b", x"7d", x"7f", x"7f", x"82", 
        x"86", x"89", x"8a", x"8c", x"8c", x"8a", x"87", x"85", x"87", x"87", x"83", x"83", x"80", x"81", x"8a", 
        x"79", x"24", x"4d", x"97", x"a3", x"94", x"8c", x"7a", x"71", x"63", x"5b", x"55", x"4c", x"41", x"3c", 
        x"38", x"3d", x"43", x"46", x"46", x"45", x"45", x"43", x"3f", x"3e", x"3c", x"37", x"30", x"2c", x"2a", 
        x"27", x"20", x"1b", x"1a", x"19", x"17", x"1c", x"24", x"45", x"4b", x"4e", x"61", x"75", x"7a", x"7d", 
        x"aa", x"a9", x"9f", x"9e", x"9c", x"9d", x"a6", x"a6", x"a5", x"a5", x"a7", x"a9", x"aa", x"a8", x"a6", 
        x"a6", x"a5", x"a5", x"a8", x"a7", x"a8", x"a7", x"a5", x"a6", x"a6", x"a6", x"a6", x"a7", x"a7", x"a6", 
        x"a4", x"a6", x"a4", x"a4", x"a9", x"a7", x"8b", x"78", x"a3", x"9b", x"72", x"5b", x"6c", x"89", x"9b", 
        x"a9", x"a9", x"a9", x"a9", x"a7", x"a8", x"a8", x"a8", x"a8", x"a9", x"a8", x"a8", x"a8", x"a9", x"a9", 
        x"a9", x"a9", x"a8", x"a8", x"a8", x"a8", x"a9", x"aa", x"aa", x"aa", x"aa", x"a9", x"a8", x"a8", x"a8", 
        x"a8", x"a9", x"a9", x"a8", x"a8", x"a8", x"a9", x"a9", x"a9", x"a9", x"a9", x"aa", x"aa", x"a9", x"a9", 
        x"a9", x"aa", x"ab", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"a9", x"a8", x"aa", x"ac", x"ac", 
        x"a9", x"ac", x"9f", x"6d", x"84", x"a2", x"a8", x"af", x"ab", x"aa", x"ad", x"aa", x"a6", x"a4", x"a7", 
        x"a6", x"a2", x"a0", x"a1", x"9a", x"74", x"76", x"55", x"66", x"76", x"69", x"72", x"7b", x"79", x"7b", 
        x"76", x"73", x"74", x"74", x"76", x"7b", x"7a", x"78", x"7a", x"7a", x"7a", x"7a", x"7a", x"79", x"79", 
        x"76", x"70", x"a1", x"e2", x"d6", x"d5", x"d5", x"d4", x"dd", x"d6", x"cf", x"d2", x"d1", x"cf", x"d1", 
        x"d2", x"d2", x"d3", x"d3", x"d3", x"d4", x"d3", x"d5", x"d0", x"cf", x"d0", x"d0", x"d3", x"d3", x"d0", 
        x"d2", x"d1", x"d1", x"d1", x"d2", x"d3", x"d3", x"d2", x"d3", x"d4", x"d5", x"d4", x"d3", x"d2", x"d3", 
        x"d4", x"d5", x"d5", x"d4", x"d3", x"d2", x"d3", x"d1", x"d2", x"d7", x"d6", x"cf", x"d2", x"d4", x"d3", 
        x"d4", x"d2", x"d0", x"e6", x"ef", x"ec", x"ed", x"ec", x"ec", x"ec", x"ec", x"ec", x"ed", x"ef", x"f1", 
        x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"ee", x"ed", x"ee", x"f0", x"ef", x"ee", x"ef", 
        x"f0", x"ec", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ee", x"ee", x"eb", x"ef", x"f2", x"ef", x"ec", 
        x"ef", x"ef", x"ee", x"ef", x"ef", x"f2", x"f2", x"f0", x"ee", x"ef", x"ee", x"e9", x"e8", x"e0", x"dc", 
        x"d6", x"ce", x"ce", x"c0", x"be", x"b3", x"b2", x"b7", x"b4", x"bc", x"b9", x"bc", x"c6", x"d0", x"da", 
        x"e5", x"ec", x"ef", x"f0", x"f2", x"f2", x"f1", x"f1", x"f2", x"f0", x"ef", x"ef", x"ef", x"e9", x"8c", 
        x"50", x"5f", x"5f", x"5f", x"5f", x"60", x"63", x"63", x"60", x"5c", x"59", x"52", x"62", x"71", x"4b", 
        x"42", x"51", x"54", x"57", x"4e", x"4b", x"4b", x"5d", x"6d", x"6e", x"6e", x"6f", x"70", x"71", x"73", 
        x"73", x"77", x"79", x"7a", x"7f", x"81", x"7d", x"69", x"55", x"3d", x"24", x"15", x"0b", x"16", x"25", 
        x"25", x"28", x"3a", x"45", x"41", x"40", x"45", x"44", x"41", x"41", x"45", x"50", x"53", x"4f", x"4b", 
        x"45", x"3d", x"32", x"26", x"21", x"1e", x"20", x"25", x"2b", x"33", x"40", x"50", x"5d", x"66", x"72", 
        x"7b", x"80", x"87", x"87", x"86", x"8b", x"8d", x"9a", x"a7", x"b8", x"c9", x"d8", x"e1", x"ea", x"ef", 
        x"f2", x"f4", x"f4", x"f3", x"f3", x"ef", x"ed", x"f0", x"f1", x"f0", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f0", x"ed", 
        x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f4", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f0", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f2", x"f3", x"f5", x"f7", x"f8", x"f7", x"f4", x"f2", x"f3", x"f7", x"f7", x"f4", x"f0", 
        x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f6", 
        x"f6", x"f4", x"f2", x"f1", x"ee", x"eb", x"e6", x"e3", x"d8", x"d5", x"cd", x"c5", x"c0", x"c1", x"c2", 
        x"c7", x"cc", x"d6", x"e1", x"eb", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f4", x"f3", x"f0", x"f4", x"f6", x"f5", x"f8", x"f5", 
        x"f5", x"f8", x"d9", x"72", x"52", x"74", x"c9", x"da", x"d5", x"d6", x"da", x"d0", x"a4", x"a6", x"a3", 
        x"9d", x"9c", x"9a", x"9a", x"9a", x"98", x"97", x"96", x"95", x"95", x"95", x"94", x"96", x"93", x"96", 
        x"9c", x"96", x"8e", x"94", x"96", x"94", x"9c", x"74", x"51", x"54", x"6e", x"70", x"5e", x"4d", x"3d", 
        x"33", x"2d", x"2d", x"35", x"47", x"57", x"5e", x"62", x"69", x"73", x"79", x"78", x"7a", x"83", x"86", 
        x"86", x"84", x"80", x"7c", x"7e", x"7d", x"7f", x"7e", x"86", x"67", x"29", x"1b", x"73", x"86", x"80", 
        x"80", x"7f", x"7f", x"7e", x"7d", x"7c", x"7e", x"7e", x"7d", x"7d", x"7e", x"7c", x"79", x"79", x"7b", 
        x"7d", x"7f", x"7f", x"80", x"81", x"84", x"89", x"8c", x"89", x"87", x"84", x"83", x"80", x"83", x"8a", 
        x"7e", x"28", x"46", x"90", x"aa", x"a4", x"a0", x"9a", x"99", x"8d", x"82", x"73", x"5a", x"41", x"36", 
        x"34", x"37", x"3e", x"41", x"41", x"43", x"46", x"45", x"45", x"46", x"44", x"41", x"40", x"40", x"3b", 
        x"32", x"26", x"20", x"23", x"27", x"25", x"19", x"20", x"4a", x"4f", x"45", x"4e", x"5a", x"6a", x"79", 
        x"a4", x"a8", x"a3", x"9b", x"9c", x"9a", x"a3", x"a2", x"a3", x"a6", x"a8", x"a7", x"a6", x"a6", x"a7", 
        x"a8", x"a8", x"a8", x"a8", x"a7", x"a6", x"a6", x"a5", x"a8", x"a9", x"a7", x"a5", x"a8", x"a7", x"a6", 
        x"a5", x"a5", x"a6", x"a7", x"a8", x"a2", x"8a", x"7e", x"94", x"a0", x"7a", x"58", x"65", x"78", x"7e", 
        x"a3", x"a7", x"a9", x"a9", x"a8", x"a9", x"a8", x"aa", x"aa", x"a9", x"a9", x"a8", x"aa", x"ab", x"ab", 
        x"aa", x"aa", x"a8", x"a8", x"a8", x"aa", x"aa", x"a9", x"aa", x"aa", x"aa", x"a9", x"a8", x"a9", x"aa", 
        x"aa", x"aa", x"aa", x"a9", x"aa", x"a9", x"ab", x"ab", x"aa", x"ac", x"ab", x"aa", x"aa", x"aa", x"ab", 
        x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"a9", x"a7", x"a9", x"ab", x"ac", 
        x"ab", x"ad", x"a1", x"70", x"84", x"a3", x"ab", x"ae", x"aa", x"a8", x"ab", x"ab", x"aa", x"a9", x"a9", 
        x"a9", x"a9", x"aa", x"ad", x"a7", x"81", x"79", x"53", x"67", x"7b", x"74", x"73", x"79", x"74", x"73", 
        x"76", x"81", x"91", x"a2", x"96", x"80", x"7b", x"79", x"79", x"7a", x"7a", x"79", x"7b", x"7d", x"7a", 
        x"77", x"70", x"a0", x"df", x"d5", x"d6", x"d6", x"d5", x"dc", x"d6", x"d0", x"d4", x"d3", x"d1", x"cf", 
        x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", x"d4", x"d4", x"d2", x"d1", x"cf", x"ce", x"d2", x"d3", x"d2", 
        x"d3", x"d3", x"d2", x"d2", x"d3", x"d3", x"d3", x"d3", x"d4", x"d5", x"d4", x"d3", x"d3", x"d3", x"d5", 
        x"d5", x"d8", x"d6", x"d4", x"d3", x"d1", x"d0", x"d3", x"d4", x"d6", x"d8", x"d1", x"d1", x"d4", x"d4", 
        x"d4", x"d3", x"d0", x"e6", x"f0", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ee", x"f0", 
        x"ef", x"ef", x"ee", x"ed", x"ed", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", 
        x"ee", x"ed", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f1", x"ef", x"ee", 
        x"f0", x"f0", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", 
        x"ef", x"ed", x"ee", x"eb", x"ea", x"e5", x"e1", x"de", x"d9", x"d6", x"c9", x"c2", x"bb", x"b3", x"b1", 
        x"b1", x"b9", x"bc", x"be", x"c7", x"cc", x"d5", x"de", x"e4", x"ec", x"ec", x"ef", x"ee", x"e6", x"93", 
        x"48", x"4b", x"4c", x"4d", x"53", x"54", x"57", x"5c", x"58", x"59", x"56", x"57", x"60", x"64", x"5c", 
        x"62", x"63", x"5c", x"5f", x"54", x"53", x"53", x"62", x"6e", x"6d", x"6e", x"6e", x"6b", x"6f", x"71", 
        x"6c", x"68", x"65", x"5e", x"53", x"42", x"30", x"1f", x"16", x"10", x"14", x"29", x"40", x"52", x"5c", 
        x"4d", x"3c", x"55", x"63", x"5d", x"62", x"61", x"61", x"5e", x"5d", x"5d", x"60", x"5f", x"5c", x"60", 
        x"62", x"60", x"5c", x"57", x"56", x"3a", x"12", x"0b", x"0e", x"0d", x"0f", x"14", x"19", x"1e", x"22", 
        x"28", x"34", x"43", x"53", x"62", x"6c", x"73", x"7e", x"80", x"88", x"89", x"89", x"8c", x"96", x"a4", 
        x"b1", x"bc", x"ce", x"d9", x"e2", x"e5", x"eb", x"ed", x"f0", x"f3", x"f1", x"f1", x"f1", x"f1", x"f3", 
        x"f2", x"f1", x"f0", x"f1", x"f0", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f2", 
        x"f3", x"f3", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"ef", x"ec", 
        x"f0", x"f2", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", 
        x"f0", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f6", x"f7", x"f8", x"f8", x"f5", x"f5", x"f5", x"f7", x"f6", x"f4", x"f3", 
        x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", 
        x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", x"f2", x"f3", x"ee", x"ee", x"ed", x"eb", x"e7", x"e4", x"da", 
        x"d2", x"c9", x"c0", x"bc", x"bb", x"c0", x"ca", x"d2", x"dd", x"e7", x"ed", x"f1", x"f2", x"f0", x"f1", 
        x"f2", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f4", x"f5", x"f2", x"f4", x"f6", x"f5", x"f6", x"f6", 
        x"f7", x"f6", x"d9", x"78", x"54", x"73", x"c5", x"d9", x"d4", x"d8", x"db", x"d2", x"a2", x"a2", x"a4", 
        x"9e", x"9d", x"9c", x"99", x"9a", x"99", x"96", x"95", x"97", x"98", x"97", x"94", x"94", x"94", x"95", 
        x"9d", x"9d", x"96", x"90", x"8b", x"80", x"6d", x"57", x"46", x"35", x"3f", x"37", x"36", x"3e", x"4c", 
        x"5c", x"68", x"6f", x"76", x"7a", x"8a", x"88", x"79", x"7a", x"7e", x"7c", x"7a", x"77", x"7e", x"82", 
        x"83", x"81", x"7f", x"7e", x"7f", x"7d", x"7f", x"7f", x"88", x"69", x"2a", x"18", x"6d", x"86", x"7e", 
        x"7e", x"80", x"80", x"7d", x"7c", x"7d", x"7e", x"7c", x"7a", x"7c", x"7e", x"7e", x"7d", x"7b", x"7b", 
        x"7c", x"7b", x"7b", x"7b", x"7b", x"7c", x"7e", x"7f", x"80", x"81", x"7e", x"80", x"80", x"84", x"87", 
        x"82", x"2d", x"3f", x"8e", x"a8", x"a2", x"9f", x"9b", x"9c", x"9b", x"95", x"92", x"86", x"71", x"65", 
        x"59", x"51", x"4c", x"48", x"40", x"3d", x"3f", x"40", x"43", x"44", x"43", x"43", x"45", x"46", x"42", 
        x"3b", x"31", x"29", x"2a", x"2e", x"2e", x"23", x"23", x"4c", x"59", x"46", x"4f", x"5a", x"63", x"76", 
        x"9f", x"a2", x"a6", x"9b", x"9b", x"a2", x"9b", x"90", x"9d", x"a5", x"a1", x"9f", x"a4", x"a8", x"a8", 
        x"a8", x"a9", x"a8", x"a5", x"a5", x"a7", x"a5", x"a2", x"a7", x"a6", x"a8", x"a8", x"a7", x"a6", x"a8", 
        x"a7", x"a6", x"a6", x"a7", x"a8", x"a5", x"a6", x"9b", x"7c", x"9e", x"8e", x"5f", x"78", x"9e", x"9a", 
        x"aa", x"a7", x"a6", x"a7", x"a8", x"a6", x"a7", x"a9", x"a8", x"a9", x"a6", x"a7", x"a8", x"a7", x"a7", 
        x"a8", x"a8", x"a8", x"a8", x"a9", x"ab", x"aa", x"a9", x"a9", x"aa", x"aa", x"a9", x"a8", x"a9", x"aa", 
        x"ab", x"ab", x"aa", x"aa", x"ac", x"aa", x"ac", x"ab", x"a9", x"ac", x"ab", x"aa", x"aa", x"aa", x"ab", 
        x"aa", x"aa", x"aa", x"a9", x"a9", x"aa", x"aa", x"aa", x"aa", x"ab", x"a9", x"a8", x"a9", x"ab", x"ac", 
        x"ab", x"ad", x"a2", x"72", x"83", x"a3", x"ab", x"ac", x"ab", x"a9", x"aa", x"a9", x"a9", x"a8", x"a8", 
        x"a8", x"a9", x"ac", x"ab", x"a4", x"85", x"7c", x"53", x"64", x"7b", x"78", x"71", x"77", x"81", x"94", 
        x"a2", x"a5", x"ab", x"b4", x"9d", x"7e", x"7d", x"7e", x"7c", x"7a", x"7a", x"7a", x"7d", x"7f", x"7a", 
        x"79", x"6f", x"a0", x"dd", x"d5", x"d8", x"d7", x"d6", x"dc", x"d7", x"cf", x"d3", x"d3", x"d1", x"d0", 
        x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", x"d4", x"d3", x"d3", x"d2", x"d0", x"cf", x"d2", x"d3", x"d1", 
        x"d3", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d4", x"d4", x"d3", x"d2", x"d3", x"d4", x"d6", 
        x"d5", x"d7", x"d6", x"d5", x"d4", x"d1", x"d0", x"d4", x"d4", x"d4", x"d8", x"d3", x"d1", x"d3", x"d2", 
        x"d2", x"d2", x"d0", x"e7", x"f1", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ed", x"ed", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f0", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"f0", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"ee", x"eb", x"e7", x"e4", 
        x"dd", x"dd", x"d5", x"cb", x"c7", x"bb", x"b4", x"af", x"ae", x"b3", x"b4", x"c3", x"cd", x"d6", x"c3", 
        x"a2", x"97", x"87", x"76", x"68", x"58", x"50", x"4e", x"4a", x"53", x"51", x"52", x"54", x"52", x"53", 
        x"59", x"58", x"5d", x"63", x"5b", x"59", x"56", x"66", x"74", x"67", x"58", x"4b", x"3b", x"36", x"2b", 
        x"23", x"1f", x"19", x"16", x"14", x"13", x"13", x"18", x"24", x"34", x"49", x"5a", x"64", x"61", x"61", 
        x"50", x"38", x"50", x"62", x"5b", x"60", x"5e", x"61", x"61", x"60", x"5f", x"5e", x"5d", x"5d", x"60", 
        x"62", x"62", x"62", x"60", x"65", x"4c", x"1a", x"11", x"29", x"31", x"27", x"20", x"14", x"0f", x"0e", 
        x"0c", x"0f", x"11", x"13", x"17", x"1a", x"1f", x"2d", x"38", x"4a", x"59", x"65", x"6f", x"7d", x"84", 
        x"86", x"82", x"81", x"7e", x"83", x"90", x"a1", x"b1", x"c4", x"d3", x"da", x"e5", x"ea", x"ed", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"f0", x"f3", x"f2", x"f1", x"f2", x"f3", x"f1", x"f2", x"f2", x"f1", x"f0", 
        x"f0", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", x"f0", x"ee", x"ee", 
        x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f3", 
        x"f3", x"f2", x"f4", x"f6", x"f7", x"f8", x"f8", x"f7", x"f5", x"f6", x"f6", x"f6", x"f5", x"f5", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f3", x"ee", x"ef", x"f4", x"f6", x"f5", x"f5", x"f2", 
        x"f0", x"ee", x"e9", x"e3", x"de", x"da", x"ca", x"bf", x"b4", x"b3", x"ba", x"c7", x"d1", x"dc", x"e1", 
        x"ea", x"ef", x"f1", x"f0", x"f1", x"ef", x"ef", x"f4", x"f6", x"f3", x"f3", x"f5", x"f5", x"f6", x"f7", 
        x"f6", x"f8", x"df", x"7d", x"50", x"6e", x"bf", x"da", x"d5", x"d5", x"d7", x"d1", x"a7", x"a3", x"a5", 
        x"9e", x"9e", x"9f", x"9c", x"9a", x"9a", x"98", x"98", x"9a", x"9b", x"9c", x"9b", x"98", x"93", x"86", 
        x"7a", x"6e", x"5d", x"50", x"42", x"31", x"2f", x"41", x"41", x"30", x"58", x"72", x"7d", x"85", x"88", 
        x"8b", x"8d", x"8b", x"84", x"79", x"84", x"84", x"76", x"76", x"7a", x"79", x"78", x"78", x"7f", x"81", 
        x"82", x"83", x"80", x"80", x"80", x"7d", x"7f", x"80", x"88", x"6e", x"2f", x"18", x"68", x"84", x"7c", 
        x"7d", x"7f", x"7f", x"7e", x"7d", x"7d", x"7c", x"7c", x"7b", x"7a", x"7d", x"7e", x"7e", x"7d", x"7c", 
        x"7d", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", x"7a", x"79", x"7b", x"76", x"78", x"78", x"7d", x"81", 
        x"81", x"31", x"3b", x"89", x"a8", x"a4", x"9f", x"9b", x"9b", x"99", x"93", x"94", x"90", x"82", x"80", 
        x"7f", x"78", x"71", x"6a", x"61", x"59", x"50", x"44", x"41", x"3f", x"3f", x"42", x"46", x"46", x"42", 
        x"3d", x"39", x"32", x"2c", x"2d", x"31", x"26", x"21", x"47", x"5d", x"4f", x"54", x"5d", x"5f", x"73", 
        x"9a", x"a5", x"a4", x"9a", x"9a", x"9e", x"9b", x"9e", x"a7", x"a2", x"9e", x"a1", x"a4", x"a7", x"a7", 
        x"a8", x"aa", x"a9", x"a5", x"a4", x"a6", x"a9", x"a9", x"a9", x"a4", x"a8", x"ab", x"a7", x"a6", x"a7", 
        x"a9", x"a7", x"a5", x"a7", x"a7", x"a6", x"a6", x"a6", x"9c", x"a4", x"a4", x"97", x"97", x"aa", x"a9", 
        x"a8", x"a7", x"a7", x"ab", x"ac", x"ab", x"ab", x"aa", x"a8", x"a9", x"a3", x"a2", x"a7", x"a9", x"a9", 
        x"a9", x"a9", x"aa", x"aa", x"ab", x"ab", x"aa", x"a9", x"a9", x"a9", x"aa", x"a9", x"a8", x"a8", x"a9", 
        x"aa", x"aa", x"a9", x"a9", x"ac", x"ab", x"ab", x"a9", x"a8", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", 
        x"aa", x"aa", x"aa", x"a9", x"a9", x"aa", x"aa", x"aa", x"aa", x"ab", x"aa", x"a9", x"ab", x"ab", x"ac", 
        x"aa", x"ad", x"a1", x"70", x"83", x"a3", x"ab", x"ab", x"ac", x"ab", x"ab", x"a9", x"a9", x"a9", x"a9", 
        x"a9", x"a9", x"ab", x"ac", x"a4", x"82", x"79", x"52", x"66", x"7a", x"76", x"7b", x"9c", x"ac", x"b0", 
        x"ae", x"ae", x"af", x"b1", x"9a", x"7f", x"7e", x"7e", x"7c", x"7b", x"7c", x"7b", x"7d", x"7f", x"7b", 
        x"7b", x"73", x"a2", x"e0", x"d7", x"d7", x"d5", x"d3", x"dc", x"d7", x"ce", x"d2", x"d1", x"d1", x"d2", 
        x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", x"d4", x"d4", x"d2", x"d3", x"d2", x"d0", x"d3", x"d3", x"d0", 
        x"d1", x"d3", x"d4", x"d3", x"d3", x"d5", x"d7", x"d5", x"d4", x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", 
        x"d4", x"d4", x"d6", x"d7", x"d4", x"d2", x"d3", x"d5", x"d4", x"d5", x"da", x"d4", x"d2", x"d3", x"d2", 
        x"d2", x"d1", x"cf", x"e5", x"ef", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ed", x"ed", x"ee", x"ef", x"ee", x"ed", x"ed", x"ed", x"ec", x"ed", x"ed", x"ee", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ed", x"ee", x"f0", x"f2", 
        x"f0", x"ef", x"f0", x"f0", x"f1", x"ef", x"ed", x"ea", x"e6", x"e4", x"d7", x"cf", x"c0", x"b9", x"bf", 
        x"c3", x"c4", x"ca", x"c4", x"c4", x"bf", x"b9", x"b0", x"a1", x"97", x"89", x"78", x"6d", x"63", x"5c", 
        x"58", x"4a", x"4f", x"52", x"55", x"59", x"5b", x"62", x"64", x"51", x"3f", x"34", x"27", x"28", x"30", 
        x"35", x"28", x"17", x"1a", x"32", x"46", x"4f", x"55", x"5d", x"60", x"5e", x"5d", x"5d", x"5b", x"5f", 
        x"58", x"3c", x"4c", x"62", x"5a", x"5f", x"60", x"61", x"62", x"62", x"61", x"61", x"62", x"63", x"62", 
        x"61", x"60", x"60", x"5f", x"63", x"52", x"1e", x"12", x"43", x"5e", x"5b", x"65", x"5e", x"56", x"4f", 
        x"44", x"38", x"2c", x"20", x"1a", x"17", x"14", x"13", x"0e", x"0c", x"0d", x"0f", x"10", x"18", x"2e", 
        x"3f", x"4e", x"5d", x"67", x"70", x"7b", x"7f", x"7e", x"7d", x"7b", x"7c", x"8b", x"94", x"9f", x"b2", 
        x"c2", x"ce", x"da", x"dd", x"e3", x"eb", x"ed", x"f1", x"f4", x"f3", x"f1", x"f1", x"f2", x"f3", x"f4", 
        x"f3", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f4", x"f2", x"ec", 
        x"f0", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f4", x"f7", x"f9", x"f9", x"f8", x"f6", x"f5", x"f5", x"f5", x"f5", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f0", x"f0", x"f2", x"f3", x"f1", x"f2", x"f2", 
        x"f2", x"f4", x"f3", x"f1", x"f0", x"f2", x"f3", x"f0", x"eb", x"e6", x"dd", x"ce", x"bf", x"ad", x"aa", 
        x"b6", x"c4", x"cd", x"d4", x"de", x"e6", x"ea", x"ef", x"f2", x"f1", x"f4", x"f8", x"f8", x"f6", x"f5", 
        x"f6", x"f9", x"e1", x"81", x"4f", x"6b", x"b9", x"db", x"d5", x"d3", x"d6", x"d2", x"a8", x"a2", x"a6", 
        x"a2", x"a1", x"9e", x"9b", x"9c", x"9c", x"9a", x"94", x"87", x"79", x"70", x"60", x"53", x"44", x"32", 
        x"32", x"41", x"4f", x"5a", x"6a", x"7c", x"86", x"7a", x"4c", x"39", x"6d", x"88", x"8c", x"8b", x"87", 
        x"86", x"87", x"88", x"84", x"74", x"7c", x"84", x"7c", x"79", x"7e", x"7c", x"78", x"79", x"80", x"80", 
        x"82", x"83", x"80", x"7f", x"7f", x"7d", x"80", x"81", x"88", x"72", x"34", x"19", x"62", x"83", x"7c", 
        x"7f", x"7e", x"7e", x"80", x"7f", x"7c", x"7b", x"7d", x"7d", x"79", x"7b", x"7d", x"7d", x"7d", x"7d", 
        x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7c", x"7b", x"7c", x"7e", x"76", x"79", x"74", x"76", x"7a", 
        x"7b", x"36", x"3f", x"81", x"a8", x"a8", x"a2", x"9d", x"9b", x"9a", x"95", x"93", x"8c", x"7f", x"7e", 
        x"7e", x"7e", x"7c", x"7c", x"7c", x"78", x"74", x"70", x"67", x"5c", x"57", x"51", x"49", x"44", x"3c", 
        x"37", x"38", x"36", x"2e", x"2e", x"36", x"2b", x"22", x"41", x"5d", x"58", x"59", x"5e", x"61", x"75", 
        x"97", x"9b", x"9f", x"a2", x"9d", x"96", x"8c", x"93", x"a0", x"a1", x"a3", x"a2", x"a1", x"a9", x"a9", 
        x"a8", x"a9", x"a9", x"a8", x"a8", x"a7", x"a8", x"a9", x"a8", x"a6", x"a6", x"a9", x"aa", x"a6", x"a6", 
        x"a9", x"a8", x"a5", x"a6", x"a8", x"a8", x"a9", x"a8", x"97", x"7f", x"8e", x"9c", x"a3", x"a7", x"ab", 
        x"ac", x"a9", x"a8", x"a8", x"a8", x"a9", x"ab", x"a9", x"a8", x"ac", x"a6", x"a4", x"aa", x"a8", x"a8", 
        x"a8", x"a9", x"aa", x"ab", x"ab", x"a9", x"a9", x"aa", x"aa", x"aa", x"a9", x"a8", x"a8", x"a9", x"a9", 
        x"a9", x"a9", x"a9", x"a9", x"ab", x"ab", x"ab", x"a9", x"a9", x"aa", x"ab", x"ab", x"ab", x"aa", x"aa", 
        x"aa", x"ab", x"ab", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"ab", x"ac", x"ab", x"ab", x"ab", x"ab", 
        x"aa", x"ac", x"9f", x"6d", x"82", x"a5", x"ad", x"ac", x"ac", x"ab", x"ab", x"a9", x"a8", x"a9", x"a9", 
        x"a9", x"a9", x"ac", x"ad", x"9f", x"81", x"81", x"57", x"67", x"7d", x"73", x"73", x"9e", x"ad", x"ab", 
        x"ac", x"ad", x"ac", x"b0", x"9c", x"82", x"81", x"7e", x"7c", x"7b", x"7d", x"7c", x"7e", x"7f", x"7c", 
        x"7c", x"72", x"a0", x"e0", x"d8", x"d8", x"d7", x"d5", x"dd", x"d7", x"ce", x"d1", x"d1", x"d1", x"d3", 
        x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", x"d4", x"d3", x"d2", x"d2", x"d1", x"d0", x"d4", x"d4", x"d0", 
        x"d0", x"d3", x"d4", x"d3", x"d3", x"d5", x"d7", x"d5", x"d3", x"d2", x"d3", x"d4", x"d3", x"d2", x"d3", 
        x"d4", x"d3", x"d6", x"d8", x"d4", x"d4", x"d6", x"d6", x"d5", x"d6", x"da", x"d4", x"d3", x"d6", x"d5", 
        x"d4", x"d2", x"cf", x"e4", x"ee", x"ec", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ee", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"f1", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f1", x"f1", 
        x"ef", x"ef", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"ed", x"ee", x"ef", x"f1", x"f0", x"ed", x"e5", 
        x"e5", x"e1", x"da", x"cf", x"c9", x"c5", x"c5", x"c6", x"c3", x"c9", x"c6", x"c0", x"bc", x"b7", x"af", 
        x"a7", x"9e", x"93", x"81", x"79", x"6c", x"66", x"5a", x"4f", x"58", x"5c", x"5a", x"50", x"4d", x"48", 
        x"4b", x"42", x"36", x"3a", x"4d", x"5d", x"61", x"5f", x"5d", x"5e", x"5d", x"5d", x"5e", x"5c", x"5d", 
        x"56", x"3b", x"48", x"60", x"58", x"5f", x"63", x"62", x"60", x"60", x"61", x"61", x"61", x"60", x"65", 
        x"63", x"61", x"61", x"62", x"65", x"54", x"23", x"11", x"41", x"5b", x"5e", x"6e", x"6b", x"6e", x"71", 
        x"70", x"6f", x"6b", x"62", x"5b", x"57", x"4f", x"48", x"3c", x"30", x"26", x"1f", x"18", x"1c", x"2c", 
        x"2c", x"23", x"22", x"1f", x"1c", x"27", x"33", x"45", x"59", x"61", x"63", x"70", x"79", x"7e", x"7f", 
        x"82", x"83", x"86", x"8a", x"9a", x"aa", x"b5", x"c0", x"cb", x"d3", x"dc", x"e6", x"ec", x"ef", x"f1", 
        x"f3", x"f3", x"f5", x"f5", x"f3", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f1", x"f1", x"ef", x"ea", 
        x"f0", x"f2", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", 
        x"f3", x"f3", x"f5", x"f7", x"f8", x"f8", x"f7", x"f6", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f0", x"ef", x"f0", x"f2", x"f0", x"f1", x"f1", 
        x"f1", x"f3", x"f2", x"f0", x"f0", x"f3", x"f4", x"f2", x"f1", x"f2", x"f3", x"f2", x"f0", x"ee", x"e8", 
        x"e1", x"d8", x"ca", x"ba", x"b6", x"ba", x"c2", x"cf", x"d8", x"dd", x"e3", x"e8", x"ee", x"f3", x"f6", 
        x"f8", x"f9", x"e2", x"88", x"4e", x"6b", x"b6", x"db", x"d6", x"d6", x"db", x"d7", x"ad", x"a3", x"a5", 
        x"9e", x"94", x"87", x"7f", x"73", x"67", x"59", x"4c", x"40", x"3d", x"3f", x"45", x"53", x"65", x"72", 
        x"81", x"8f", x"9b", x"9e", x"98", x"95", x"95", x"81", x"4a", x"3c", x"6d", x"87", x"8a", x"89", x"87", 
        x"88", x"8a", x"8a", x"84", x"73", x"78", x"83", x"7c", x"76", x"7d", x"81", x"78", x"77", x"80", x"83", 
        x"83", x"82", x"80", x"7f", x"7e", x"7e", x"81", x"81", x"86", x"74", x"36", x"18", x"5c", x"83", x"7e", 
        x"80", x"7f", x"7e", x"7f", x"7f", x"7d", x"7c", x"7d", x"7c", x"79", x"7b", x"7c", x"7c", x"7b", x"7c", 
        x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7b", x"79", x"7c", x"76", x"7d", x"78", x"7a", x"7d", 
        x"7f", x"49", x"51", x"85", x"aa", x"a7", x"a4", x"a1", x"9d", x"9b", x"98", x"94", x"8c", x"81", x"7f", 
        x"7f", x"7f", x"80", x"81", x"82", x"80", x"7e", x"7e", x"7a", x"7a", x"78", x"72", x"6a", x"65", x"5b", 
        x"4b", x"3e", x"35", x"2b", x"2b", x"32", x"2b", x"21", x"3d", x"5e", x"57", x"58", x"64", x"68", x"7b", 
        x"92", x"97", x"93", x"97", x"9c", x"90", x"94", x"a0", x"a2", x"9f", x"a3", x"a5", x"a5", x"a8", x"aa", 
        x"a9", x"a7", x"a7", x"a9", x"aa", x"a9", x"a7", x"a7", x"a7", x"a9", x"a5", x"a6", x"aa", x"a8", x"a7", 
        x"a8", x"a8", x"a7", x"a7", x"a8", x"a8", x"a9", x"9f", x"82", x"6c", x"7d", x"90", x"9f", x"a7", x"aa", 
        x"aa", x"a6", x"a8", x"a8", x"a8", x"a9", x"ab", x"a9", x"a8", x"ac", x"a7", x"a5", x"a7", x"a5", x"a6", 
        x"a8", x"aa", x"ab", x"ac", x"aa", x"a9", x"aa", x"ab", x"ab", x"aa", x"a9", x"a8", x"a9", x"a9", x"aa", 
        x"aa", x"aa", x"aa", x"aa", x"aa", x"ab", x"aa", x"aa", x"ab", x"ab", x"ac", x"ac", x"ab", x"ab", x"ab", 
        x"ab", x"ab", x"ac", x"ab", x"aa", x"ab", x"ab", x"ab", x"ab", x"ac", x"ad", x"ac", x"ad", x"ac", x"ac", 
        x"ab", x"ad", x"a1", x"6e", x"82", x"a4", x"ac", x"ac", x"ac", x"ac", x"ac", x"aa", x"a9", x"a9", x"aa", 
        x"aa", x"aa", x"ad", x"ac", x"a1", x"9b", x"a0", x"63", x"65", x"79", x"74", x"76", x"a2", x"ae", x"ae", 
        x"ad", x"ac", x"ac", x"b0", x"9c", x"81", x"80", x"80", x"7e", x"7b", x"7d", x"7c", x"7e", x"7f", x"7c", 
        x"7c", x"73", x"9f", x"e1", x"d8", x"d7", x"d6", x"d5", x"dc", x"d7", x"ce", x"d0", x"d0", x"d1", x"d4", 
        x"d4", x"d4", x"d4", x"d3", x"d3", x"d3", x"d4", x"d4", x"d2", x"d2", x"d1", x"d0", x"d4", x"d5", x"d1", 
        x"d0", x"d3", x"d5", x"d4", x"d3", x"d4", x"d6", x"d3", x"d3", x"d3", x"d3", x"d3", x"d2", x"d1", x"d2", 
        x"d4", x"d4", x"d6", x"d8", x"d5", x"d5", x"d6", x"d5", x"d4", x"d6", x"d9", x"d3", x"d3", x"d6", x"d5", 
        x"d4", x"d3", x"d0", x"e6", x"ef", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ed", x"ee", x"ef", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"f0", x"f3", x"f2", x"ee", 
        x"ee", x"ef", x"f1", x"ef", x"ef", x"ed", x"ed", x"ee", x"ed", x"ee", x"f1", x"f0", x"ef", x"ee", x"e7", 
        x"f1", x"f2", x"ef", x"ee", x"f0", x"ef", x"ec", x"e8", x"e2", x"de", x"d8", x"ce", x"c8", x"c5", x"c6", 
        x"c5", x"c6", x"c8", x"c2", x"c4", x"bd", x"b9", x"ac", x"9e", x"95", x"87", x"7c", x"70", x"6c", x"68", 
        x"66", x"61", x"5c", x"57", x"53", x"54", x"57", x"5b", x"5c", x"5f", x"63", x"63", x"65", x"64", x"67", 
        x"64", x"43", x"48", x"5f", x"5f", x"60", x"60", x"60", x"5e", x"5c", x"5d", x"5f", x"5f", x"5e", x"5f", 
        x"61", x"62", x"63", x"65", x"68", x"5b", x"2c", x"16", x"41", x"5c", x"62", x"70", x"6b", x"6e", x"6e", 
        x"6c", x"6c", x"6d", x"6c", x"6e", x"71", x"71", x"73", x"73", x"6d", x"64", x"57", x"4a", x"48", x"58", 
        x"5c", x"57", x"52", x"49", x"3e", x"37", x"2f", x"28", x"25", x"20", x"1d", x"24", x"2d", x"3e", x"4e", 
        x"5c", x"5f", x"61", x"68", x"73", x"7a", x"7e", x"82", x"85", x"8b", x"98", x"a6", x"b0", x"b9", x"c3", 
        x"cf", x"d7", x"e1", x"e5", x"ec", x"ef", x"f2", x"f3", x"f4", x"f4", x"f3", x"f2", x"f1", x"ee", x"ed", 
        x"f2", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f3", x"f4", x"f5", x"f6", x"f7", x"f7", x"f7", x"f6", x"f3", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f3", x"f0", x"f0", x"f1", x"f2", x"f0", x"f1", x"f0", 
        x"f0", x"f2", x"f2", x"f1", x"f1", x"f4", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f0", x"f1", 
        x"f2", x"f1", x"ef", x"ec", x"e8", x"df", x"d7", x"d0", x"c8", x"c1", x"c3", x"ca", x"d2", x"da", x"e1", 
        x"e4", x"e8", x"dc", x"8d", x"50", x"72", x"b7", x"dd", x"d8", x"d2", x"c6", x"b6", x"8d", x"79", x"6c", 
        x"5b", x"4d", x"46", x"45", x"41", x"45", x"51", x"60", x"70", x"7f", x"8c", x"94", x"9a", x"9e", x"9a", 
        x"95", x"95", x"98", x"99", x"91", x"90", x"95", x"83", x"4c", x"3f", x"66", x"86", x"89", x"8a", x"88", 
        x"87", x"88", x"87", x"83", x"75", x"78", x"81", x"7c", x"78", x"7e", x"85", x"7a", x"76", x"81", x"87", 
        x"86", x"82", x"80", x"7f", x"7f", x"7e", x"80", x"80", x"85", x"77", x"39", x"19", x"57", x"84", x"7e", 
        x"7e", x"7f", x"7f", x"7e", x"7e", x"7e", x"7e", x"7d", x"7c", x"7c", x"7c", x"7c", x"7b", x"7b", x"7b", 
        x"7d", x"7c", x"7d", x"7c", x"7c", x"7c", x"7b", x"7a", x"7a", x"7c", x"76", x"7d", x"77", x"78", x"7b", 
        x"7d", x"4e", x"56", x"85", x"aa", x"a9", x"a6", x"a5", x"9e", x"9c", x"99", x"95", x"8f", x"84", x"7f", 
        x"7c", x"7e", x"81", x"82", x"81", x"7f", x"7e", x"80", x"81", x"83", x"82", x"7e", x"7d", x"7d", x"77", 
        x"6e", x"66", x"5f", x"54", x"46", x"3c", x"35", x"27", x"39", x"5d", x"55", x"59", x"6c", x"6e", x"7e", 
        x"bb", x"b5", x"a3", x"94", x"9c", x"8d", x"93", x"98", x"88", x"89", x"97", x"9f", x"a0", x"a7", x"ab", 
        x"aa", x"a9", x"a8", x"a8", x"a8", x"a7", x"a7", x"a8", x"a8", x"a8", x"a8", x"a9", x"a9", x"ae", x"a8", 
        x"a7", x"a8", x"a9", x"a7", x"a7", x"a9", x"a6", x"97", x"9e", x"98", x"8b", x"9f", x"ac", x"ab", x"aa", 
        x"a9", x"a6", x"a8", x"aa", x"a8", x"a7", x"a9", x"a8", x"a5", x"a9", x"a9", x"a5", x"a6", x"a7", x"a9", 
        x"ab", x"ab", x"ab", x"ab", x"aa", x"aa", x"ab", x"ac", x"ab", x"a9", x"aa", x"aa", x"ab", x"aa", x"aa", 
        x"aa", x"ab", x"ac", x"ab", x"a9", x"ac", x"ab", x"ab", x"ad", x"ab", x"ab", x"ac", x"ac", x"ac", x"ac", 
        x"ac", x"ac", x"ac", x"ab", x"ab", x"ab", x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", 
        x"aa", x"ae", x"a2", x"70", x"82", x"a2", x"aa", x"ac", x"ad", x"ac", x"ac", x"aa", x"aa", x"a9", x"a9", 
        x"a9", x"aa", x"aa", x"a9", x"a5", x"af", x"ae", x"63", x"63", x"7c", x"76", x"78", x"a5", x"af", x"ad", 
        x"ac", x"aa", x"ab", x"b0", x"9a", x"7d", x"7e", x"7d", x"7c", x"7b", x"7c", x"7b", x"7e", x"80", x"7c", 
        x"7c", x"73", x"9e", x"e0", x"d7", x"d5", x"d7", x"d5", x"db", x"d6", x"cf", x"d1", x"d0", x"d2", x"d4", 
        x"d4", x"d4", x"d4", x"d3", x"d3", x"d3", x"d4", x"d3", x"d1", x"d2", x"d1", x"d0", x"d4", x"d5", x"d1", 
        x"d0", x"d3", x"d5", x"d5", x"d4", x"d4", x"d4", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", x"d1", x"d1", 
        x"d3", x"d6", x"d6", x"d6", x"d6", x"d6", x"d4", x"d4", x"d4", x"d5", x"d6", x"d0", x"d3", x"d5", x"d2", 
        x"d3", x"d3", x"d0", x"e8", x"f2", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"ee", x"ef", x"ef", x"f0", x"ef", x"ef", x"ee", x"ed", x"ef", x"f1", x"ee", x"ea", 
        x"ed", x"ef", x"ee", x"ed", x"ef", x"f0", x"ef", x"f0", x"f0", x"ee", x"ee", x"ec", x"f1", x"ed", x"e4", 
        x"ed", x"ee", x"ed", x"ee", x"ef", x"f0", x"f0", x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f2", x"f0", 
        x"ec", x"e1", x"de", x"d3", x"d1", x"cf", x"ca", x"c4", x"c2", x"cc", x"cd", x"cb", x"c5", x"bc", x"af", 
        x"a8", x"9f", x"92", x"83", x"77", x"6e", x"66", x"62", x"5d", x"5a", x"57", x"52", x"56", x"5c", x"60", 
        x"5f", x"50", x"58", x"66", x"69", x"6b", x"6c", x"68", x"66", x"63", x"61", x"60", x"5f", x"5f", x"5c", 
        x"5e", x"60", x"5f", x"60", x"63", x"5e", x"2f", x"15", x"41", x"5f", x"66", x"72", x"6e", x"73", x"73", 
        x"70", x"6f", x"6f", x"6d", x"6e", x"6f", x"6e", x"6e", x"6e", x"6f", x"6e", x"65", x"5e", x"59", x"5f", 
        x"5e", x"5f", x"5d", x"5d", x"60", x"64", x"60", x"5c", x"59", x"50", x"44", x"3b", x"31", x"2a", x"13", 
        x"09", x"12", x"22", x"25", x"2f", x"3c", x"49", x"57", x"61", x"63", x"6a", x"73", x"7a", x"7f", x"83", 
        x"8c", x"94", x"a1", x"a8", x"b1", x"b9", x"c3", x"cc", x"d7", x"e3", x"eb", x"ef", x"f6", x"f0", x"ed", 
        x"ef", x"f5", x"f3", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f4", x"f3", 
        x"f3", x"f4", x"f5", x"f6", x"f7", x"f7", x"f7", x"f5", x"f3", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f4", x"f1", x"f1", x"f1", x"f2", x"f1", x"f3", x"f2", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f4", x"f2", x"f1", x"f1", x"f1", x"f0", x"f2", x"f3", x"f1", x"f3", 
        x"f1", x"ee", x"ef", x"f2", x"ef", x"f2", x"f5", x"f6", x"f5", x"ec", x"e4", x"de", x"d5", x"cf", x"ce", 
        x"cd", x"cc", x"c3", x"85", x"4f", x"6e", x"8d", x"95", x"80", x"72", x"63", x"5a", x"48", x"41", x"45", 
        x"4a", x"58", x"70", x"84", x"97", x"9c", x"a0", x"a1", x"a0", x"9d", x"99", x"94", x"94", x"96", x"93", 
        x"91", x"92", x"94", x"9a", x"94", x"90", x"93", x"86", x"4f", x"44", x"64", x"86", x"85", x"85", x"87", 
        x"89", x"87", x"86", x"84", x"75", x"76", x"7c", x"7b", x"78", x"7b", x"87", x"7f", x"76", x"81", x"89", 
        x"86", x"83", x"81", x"80", x"80", x"7e", x"7f", x"7d", x"83", x"79", x"3c", x"19", x"50", x"82", x"7d", 
        x"7c", x"7f", x"80", x"7e", x"7e", x"7f", x"7f", x"7d", x"7c", x"7d", x"7e", x"7d", x"7c", x"7b", x"7c", 
        x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", x"7b", x"7e", x"7d", x"79", x"7c", x"77", x"77", x"7c", 
        x"7f", x"50", x"53", x"84", x"a9", x"a9", x"a4", x"a3", x"9d", x"9e", x"9d", x"99", x"93", x"83", x"7a", 
        x"7b", x"7c", x"7d", x"7f", x"80", x"81", x"81", x"7f", x"81", x"81", x"7f", x"7f", x"84", x"88", x"88", 
        x"84", x"82", x"83", x"81", x"7a", x"72", x"64", x"44", x"35", x"58", x"55", x"54", x"66", x"6e", x"7c", 
        x"d2", x"c7", x"c7", x"ba", x"c1", x"b1", x"ac", x"a3", x"8d", x"92", x"99", x"98", x"97", x"98", x"9d", 
        x"a1", x"a7", x"a8", x"a7", x"a6", x"a8", x"a9", x"a9", x"ac", x"a8", x"ac", x"a6", x"90", x"a1", x"a9", 
        x"a6", x"a7", x"aa", x"a8", x"a7", x"a9", x"a8", x"a4", x"ab", x"a7", x"95", x"97", x"a0", x"a5", x"a8", 
        x"ab", x"a9", x"a7", x"ab", x"ab", x"a9", x"a8", x"a8", x"a4", x"a7", x"ab", x"a6", x"a4", x"a6", x"a9", 
        x"ab", x"ac", x"ab", x"aa", x"a9", x"ac", x"ac", x"ab", x"a9", x"a9", x"ac", x"ad", x"ac", x"ab", x"aa", 
        x"aa", x"ab", x"ac", x"ac", x"aa", x"ad", x"ac", x"ad", x"ad", x"a9", x"a9", x"ab", x"ab", x"ac", x"ac", 
        x"ac", x"ac", x"ab", x"ab", x"ab", x"ac", x"ac", x"ac", x"ac", x"ad", x"ad", x"ad", x"ac", x"ac", x"ac", 
        x"ab", x"af", x"a3", x"70", x"82", x"a3", x"ac", x"ad", x"ac", x"ab", x"ab", x"ab", x"aa", x"a9", x"a8", 
        x"a9", x"ab", x"aa", x"a9", x"a3", x"ab", x"ab", x"63", x"62", x"7c", x"76", x"73", x"a3", x"ae", x"ab", 
        x"ab", x"aa", x"ac", x"af", x"98", x"7e", x"82", x"7f", x"7c", x"7b", x"7b", x"7a", x"7e", x"80", x"7c", 
        x"7b", x"71", x"9b", x"df", x"d6", x"d5", x"d7", x"d6", x"da", x"d6", x"cf", x"d2", x"d0", x"d2", x"d4", 
        x"d4", x"d4", x"d4", x"d3", x"d3", x"d3", x"d4", x"d2", x"cf", x"d1", x"d2", x"d1", x"d4", x"d3", x"d0", 
        x"d2", x"d3", x"d4", x"d5", x"d4", x"d3", x"d2", x"d3", x"d3", x"d3", x"d2", x"d1", x"d2", x"d3", x"d1", 
        x"d2", x"d7", x"d6", x"d4", x"d6", x"d6", x"d5", x"d5", x"d6", x"d7", x"d7", x"d1", x"d5", x"d5", x"d2", 
        x"d2", x"d2", x"cf", x"e6", x"f0", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", 
        x"ef", x"f0", x"ee", x"ee", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"f0", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"ed", 
        x"f1", x"ef", x"ec", x"ed", x"ef", x"f1", x"ee", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"f0", x"e7", 
        x"ed", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ee", x"ee", x"f0", x"f0", x"ef", 
        x"ef", x"f0", x"ef", x"f2", x"f1", x"ed", x"ee", x"eb", x"e6", x"e4", x"df", x"de", x"da", x"d2", x"cf", 
        x"d2", x"d0", x"cc", x"c7", x"c4", x"be", x"b4", x"ad", x"a6", x"9b", x"92", x"87", x"81", x"79", x"6f", 
        x"61", x"57", x"56", x"50", x"50", x"54", x"59", x"5b", x"61", x"68", x"6a", x"69", x"6a", x"6c", x"6a", 
        x"65", x"62", x"61", x"62", x"62", x"60", x"30", x"11", x"40", x"64", x"66", x"70", x"70", x"73", x"73", 
        x"71", x"72", x"72", x"72", x"73", x"74", x"72", x"71", x"6f", x"70", x"6d", x"60", x"5a", x"58", x"5c", 
        x"59", x"5a", x"5a", x"5b", x"5a", x"5b", x"59", x"5b", x"5d", x"5f", x"60", x"5d", x"5f", x"57", x"29", 
        x"18", x"30", x"53", x"49", x"3d", x"31", x"24", x"1c", x"1b", x"1b", x"22", x"2e", x"3d", x"43", x"49", 
        x"50", x"59", x"6a", x"74", x"81", x"89", x"91", x"96", x"9a", x"a1", x"a9", x"b5", x"b9", x"c6", x"e6", 
        x"f3", x"f5", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f4", x"f3", 
        x"f3", x"f3", x"f5", x"f7", x"f8", x"f7", x"f6", x"f4", x"f3", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f5", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"ef", 
        x"f0", x"f2", x"f2", x"f0", x"ef", x"f1", x"f1", x"f1", x"f2", x"f4", x"f5", x"f3", x"f0", x"f0", x"f2", 
        x"f0", x"ef", x"f0", x"f3", x"f0", x"f1", x"f1", x"f0", x"f2", x"f2", x"f5", x"f6", x"f7", x"f4", x"f0", 
        x"ed", x"e6", x"d6", x"93", x"40", x"43", x"56", x"5d", x"53", x"5a", x"6c", x"82", x"87", x"93", x"a6", 
        x"a7", x"a3", x"a1", x"a0", x"9d", x"9b", x"98", x"96", x"96", x"97", x"95", x"95", x"92", x"93", x"92", 
        x"92", x"92", x"92", x"96", x"96", x"92", x"92", x"8b", x"50", x"41", x"60", x"84", x"86", x"86", x"87", 
        x"89", x"8b", x"8b", x"87", x"75", x"73", x"79", x"7d", x"7b", x"79", x"86", x"85", x"79", x"80", x"88", 
        x"85", x"87", x"82", x"81", x"82", x"7f", x"7e", x"7b", x"81", x"79", x"3c", x"16", x"4a", x"81", x"7e", 
        x"7e", x"80", x"80", x"80", x"7f", x"7e", x"7d", x"7c", x"7c", x"7c", x"7d", x"7c", x"7c", x"7c", x"7e", 
        x"7f", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7c", x"7c", x"7a", x"7a", x"7d", x"7a", x"76", x"7b", 
        x"81", x"51", x"51", x"84", x"a7", x"ab", x"a7", x"a5", x"9e", x"9f", x"9c", x"99", x"95", x"82", x"73", 
        x"76", x"78", x"77", x"76", x"79", x"78", x"78", x"83", x"88", x"88", x"87", x"87", x"88", x"88", x"8a", 
        x"89", x"8a", x"8c", x"8c", x"88", x"85", x"82", x"5c", x"32", x"5f", x"73", x"69", x"71", x"73", x"7a", 
        x"b9", x"c1", x"d0", x"c6", x"d4", x"d1", x"d4", x"cd", x"ca", x"c3", x"c3", x"c2", x"b8", x"af", x"a8", 
        x"9e", x"9e", x"8f", x"96", x"9e", x"a2", x"a6", x"a8", x"ad", x"9e", x"9a", x"8a", x"6e", x"87", x"a8", 
        x"a7", x"a7", x"a9", x"ab", x"aa", x"a7", x"a9", x"a7", x"ac", x"a8", x"91", x"8a", x"9e", x"a9", x"a9", 
        x"a8", x"a8", x"a9", x"a7", x"aa", x"aa", x"aa", x"aa", x"a9", x"a2", x"a6", x"a1", x"a1", x"a4", x"a6", 
        x"a9", x"aa", x"aa", x"a9", x"a9", x"aa", x"ab", x"aa", x"aa", x"aa", x"aa", x"ac", x"ac", x"aa", x"ab", 
        x"ac", x"ab", x"aa", x"ac", x"ab", x"ab", x"aa", x"ac", x"ae", x"ab", x"a9", x"aa", x"ab", x"ac", x"ad", 
        x"ad", x"ac", x"ab", x"ab", x"ac", x"ad", x"ad", x"ad", x"ad", x"ad", x"ad", x"ad", x"ac", x"ab", x"aa", 
        x"aa", x"ad", x"a4", x"6f", x"80", x"a4", x"ac", x"ad", x"ac", x"ab", x"ab", x"ac", x"ab", x"aa", x"a9", 
        x"aa", x"ab", x"ab", x"ad", x"a5", x"ad", x"ab", x"64", x"61", x"7e", x"7a", x"76", x"a3", x"ae", x"ac", 
        x"ad", x"ac", x"ae", x"af", x"9a", x"80", x"81", x"7f", x"7e", x"7b", x"79", x"79", x"7d", x"7f", x"7b", 
        x"7a", x"75", x"9b", x"de", x"d8", x"d5", x"d6", x"d5", x"d9", x"d7", x"cf", x"d2", x"d1", x"d0", x"d1", 
        x"d2", x"d2", x"d4", x"d4", x"d4", x"d4", x"d4", x"d3", x"d1", x"d3", x"d2", x"d2", x"d3", x"d3", x"d1", 
        x"d0", x"d1", x"d4", x"d5", x"d5", x"d3", x"d0", x"d2", x"d4", x"d3", x"d3", x"d3", x"d5", x"d3", x"d0", 
        x"d3", x"d8", x"d7", x"d6", x"d8", x"d6", x"d5", x"d5", x"d5", x"d6", x"d9", x"d3", x"d5", x"d7", x"d3", 
        x"d1", x"d0", x"d0", x"e5", x"f0", x"ed", x"ed", x"ed", x"ec", x"ed", x"ee", x"ed", x"ed", x"ee", x"ef", 
        x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", 
        x"f0", x"ef", x"ed", x"ed", x"ee", x"f0", x"ee", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"f0", x"e7", 
        x"ed", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ee", x"ef", x"ef", x"ee", 
        x"ef", x"f0", x"ee", x"f1", x"ef", x"ed", x"f1", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"ee", x"eb", 
        x"e9", x"e7", x"e3", x"df", x"dc", x"da", x"d7", x"d5", x"d2", x"ce", x"cb", x"c7", x"c3", x"bc", x"b4", 
        x"a8", x"9d", x"93", x"87", x"80", x"7a", x"76", x"68", x"5f", x"5a", x"53", x"52", x"52", x"58", x"5e", 
        x"5f", x"61", x"66", x"6a", x"6a", x"6d", x"48", x"2b", x"4d", x"6a", x"6f", x"81", x"84", x"80", x"7c", 
        x"79", x"76", x"75", x"76", x"75", x"75", x"73", x"74", x"73", x"73", x"73", x"65", x"63", x"5a", x"5c", 
        x"5a", x"5a", x"5a", x"5c", x"5d", x"5a", x"58", x"5b", x"5e", x"5d", x"5d", x"5d", x"63", x"5d", x"2a", 
        x"1c", x"2d", x"4a", x"45", x"3e", x"37", x"36", x"38", x"35", x"31", x"35", x"3f", x"44", x"39", x"2c", 
        x"25", x"27", x"2e", x"34", x"3f", x"46", x"52", x"5b", x"63", x"6b", x"68", x"63", x"58", x"98", x"e0", 
        x"f5", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", 
        x"f4", x"f3", x"f5", x"f7", x"f8", x"f6", x"f3", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f5", x"f2", x"f0", x"f1", x"f2", x"f0", x"f2", x"f0", 
        x"f1", x"f2", x"f1", x"f0", x"f0", x"f2", x"f0", x"f0", x"f0", x"f2", x"f3", x"f3", x"f1", x"ef", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"ef", x"f0", x"f1", x"f2", x"f5", x"f5", x"f6", x"f5", 
        x"f6", x"f7", x"ee", x"a9", x"3c", x"3a", x"7d", x"bd", x"bd", x"b7", x"b0", x"ac", x"90", x"81", x"89", 
        x"8c", x"89", x"8c", x"94", x"97", x"9c", x"9c", x"9c", x"9a", x"97", x"95", x"97", x"95", x"92", x"91", 
        x"91", x"92", x"92", x"95", x"98", x"94", x"93", x"8f", x"53", x"44", x"5d", x"84", x"89", x"88", x"85", 
        x"86", x"89", x"89", x"83", x"73", x"72", x"75", x"7a", x"79", x"7a", x"85", x"88", x"7e", x"7e", x"84", 
        x"84", x"87", x"82", x"7f", x"7f", x"7f", x"80", x"7d", x"81", x"7b", x"49", x"21", x"3f", x"81", x"80", 
        x"80", x"80", x"80", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7c", x"7d", x"7c", x"7c", x"7e", x"7e", 
        x"7e", x"7e", x"7f", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7c", x"77", x"7d", x"7b", x"74", x"79", 
        x"81", x"59", x"4c", x"7c", x"a5", x"aa", x"a6", x"a7", x"a0", x"a1", x"9e", x"9b", x"98", x"89", x"79", 
        x"7a", x"7b", x"7a", x"74", x"74", x"71", x"6e", x"87", x"90", x"8c", x"8c", x"8b", x"8c", x"89", x"89", 
        x"89", x"88", x"88", x"8a", x"8b", x"89", x"8b", x"70", x"35", x"5f", x"81", x"7a", x"83", x"84", x"7f", 
        x"d6", x"d4", x"d1", x"ce", x"af", x"9c", x"bc", x"ba", x"cb", x"d2", x"df", x"e0", x"e7", x"e8", x"e3", 
        x"da", x"d2", x"bd", x"b3", x"a6", x"9c", x"97", x"90", x"95", x"8d", x"76", x"73", x"7c", x"8f", x"ab", 
        x"a9", x"a8", x"a6", x"9e", x"a4", x"a9", x"a7", x"a7", x"a5", x"99", x"88", x"99", x"b0", x"ad", x"ab", 
        x"b3", x"a9", x"a5", x"a9", x"a7", x"a8", x"ab", x"a4", x"98", x"8e", x"9e", x"a0", x"9e", x"9e", x"9f", 
        x"a1", x"aa", x"ab", x"aa", x"ad", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"ac", 
        x"ad", x"ac", x"aa", x"ab", x"ad", x"ac", x"ab", x"ad", x"af", x"af", x"ad", x"ac", x"ac", x"ac", x"ad", 
        x"ad", x"ac", x"ac", x"ac", x"ad", x"ad", x"ad", x"ad", x"ad", x"ad", x"ad", x"ae", x"ab", x"ac", x"a9", 
        x"ab", x"ad", x"a5", x"72", x"80", x"a4", x"ac", x"ac", x"ac", x"ad", x"ac", x"ac", x"ab", x"ab", x"ab", 
        x"ab", x"ab", x"ab", x"ae", x"a5", x"ad", x"aa", x"64", x"63", x"7f", x"79", x"77", x"a2", x"ac", x"a9", 
        x"ac", x"ad", x"ad", x"af", x"9e", x"81", x"7e", x"7e", x"7f", x"7b", x"7a", x"7a", x"7d", x"7e", x"7c", 
        x"79", x"77", x"9a", x"dd", x"da", x"d6", x"d6", x"d5", x"da", x"d7", x"ce", x"d2", x"d2", x"d0", x"d0", 
        x"d3", x"d3", x"d2", x"d1", x"d0", x"d1", x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", x"d4", x"d4", x"d2", 
        x"cf", x"d0", x"d4", x"d4", x"d5", x"d3", x"d0", x"d3", x"d5", x"d4", x"d3", x"d4", x"d4", x"d1", x"d0", 
        x"d5", x"d7", x"d6", x"d7", x"d7", x"d6", x"d6", x"d6", x"d5", x"d7", x"da", x"d3", x"d1", x"d4", x"d3", 
        x"d2", x"d0", x"cf", x"e4", x"f1", x"ed", x"ee", x"ec", x"ec", x"ee", x"ee", x"ed", x"ed", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ee", x"ee", x"f1", x"f0", x"e5", 
        x"ec", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f2", x"ef", x"ec", x"eb", x"ec", x"ea", x"e7", x"e4", x"e2", x"e1", x"dd", 
        x"d2", x"d0", x"ce", x"cc", x"c8", x"c3", x"bf", x"b5", x"ad", x"ac", x"a3", x"99", x"89", x"81", x"6f", 
        x"65", x"58", x"4b", x"46", x"45", x"4d", x"5b", x"54", x"60", x"6c", x"6a", x"71", x"78", x"7a", x"7a", 
        x"7e", x"81", x"82", x"81", x"7e", x"7f", x"7c", x"7a", x"77", x"73", x"73", x"64", x"61", x"5d", x"5b", 
        x"5b", x"5b", x"5d", x"5d", x"5d", x"5a", x"59", x"5c", x"60", x"5f", x"60", x"60", x"59", x"4c", x"1d", 
        x"12", x"19", x"30", x"3a", x"4c", x"56", x"5b", x"64", x"67", x"69", x"6d", x"70", x"6e", x"69", x"64", 
        x"60", x"5c", x"57", x"4e", x"4a", x"4a", x"37", x"20", x"19", x"20", x"48", x"65", x"87", x"c9", x"e5", 
        x"f0", x"f4", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"f0", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f5", 
        x"f5", x"f3", x"f6", x"f8", x"f8", x"f5", x"f2", x"f0", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f6", x"f2", x"ef", x"f2", x"f3", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"f0", x"ef", x"f1", x"f0", x"f2", x"f6", x"f5", x"f5", x"f5", 
        x"f5", x"f5", x"ef", x"ac", x"41", x"4b", x"95", x"db", x"d9", x"d7", x"d4", x"d2", x"b0", x"91", x"92", 
        x"8c", x"7a", x"6e", x"6c", x"68", x"71", x"7a", x"84", x"90", x"97", x"9f", x"9f", x"9c", x"9a", x"97", 
        x"94", x"90", x"8e", x"92", x"98", x"94", x"93", x"90", x"55", x"43", x"59", x"83", x"8b", x"8b", x"87", 
        x"86", x"85", x"87", x"86", x"75", x"72", x"70", x"74", x"77", x"7a", x"82", x"86", x"81", x"7e", x"84", 
        x"85", x"88", x"82", x"7f", x"7e", x"7f", x"82", x"7f", x"81", x"81", x"58", x"35", x"3b", x"80", x"81", 
        x"7f", x"81", x"81", x"7e", x"7d", x"7e", x"7e", x"7d", x"7c", x"7c", x"7d", x"7c", x"7c", x"7d", x"7e", 
        x"7d", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7e", x"7e", x"76", x"7d", x"7d", x"76", x"7a", 
        x"7f", x"5e", x"46", x"78", x"a6", x"b0", x"ab", x"a5", x"a0", x"a3", x"9d", x"9e", x"99", x"89", x"78", 
        x"75", x"77", x"78", x"72", x"74", x"74", x"71", x"8c", x"96", x"8e", x"8b", x"89", x"8b", x"8a", x"8a", 
        x"8d", x"8b", x"89", x"8b", x"8b", x"87", x"8c", x"7b", x"38", x"5a", x"7e", x"7c", x"89", x"8f", x"88", 
        x"cc", x"c5", x"ca", x"cf", x"aa", x"91", x"a9", x"c1", x"d0", x"e0", x"e9", x"e9", x"ef", x"ea", x"e8", 
        x"e9", x"e4", x"e9", x"e6", x"e6", x"df", x"d5", x"c4", x"bb", x"ad", x"8b", x"80", x"90", x"8d", x"89", 
        x"8f", x"a7", x"a8", x"9f", x"93", x"8f", x"a3", x"ad", x"ab", x"9b", x"88", x"9f", x"a8", x"94", x"80", 
        x"96", x"9f", x"a8", x"aa", x"aa", x"aa", x"aa", x"a9", x"a5", x"9a", x"9d", x"9c", x"a1", x"a7", x"a6", 
        x"a4", x"a7", x"a9", x"a7", x"a9", x"ab", x"ab", x"aa", x"a9", x"a9", x"aa", x"aa", x"ab", x"ab", x"ac", 
        x"ab", x"ac", x"ab", x"aa", x"ac", x"ac", x"ac", x"ad", x"ae", x"ad", x"ad", x"ac", x"ac", x"ab", x"ab", 
        x"ab", x"ac", x"ac", x"ac", x"ad", x"ac", x"ac", x"ab", x"ab", x"ab", x"ac", x"ae", x"ab", x"ac", x"aa", 
        x"ac", x"ae", x"a5", x"74", x"80", x"a4", x"ab", x"ab", x"ac", x"ab", x"ac", x"ac", x"ab", x"ab", x"ab", 
        x"ab", x"ab", x"ac", x"ae", x"a4", x"ac", x"aa", x"65", x"64", x"7c", x"75", x"74", x"a1", x"ac", x"a8", 
        x"ab", x"ac", x"ad", x"b0", x"9f", x"81", x"7f", x"7f", x"7f", x"7b", x"7c", x"7d", x"7d", x"7d", x"7c", 
        x"7a", x"76", x"9a", x"dd", x"d8", x"d6", x"d6", x"d5", x"db", x"d8", x"ce", x"d1", x"d2", x"d1", x"d1", 
        x"d4", x"d5", x"d4", x"d2", x"d1", x"d1", x"d4", x"d2", x"d2", x"d3", x"d2", x"d2", x"d4", x"d4", x"d1", 
        x"ce", x"d0", x"d4", x"d2", x"d2", x"d4", x"d2", x"d4", x"d5", x"d4", x"d3", x"d4", x"d3", x"d1", x"d3", 
        x"d6", x"d7", x"d5", x"d4", x"d4", x"d4", x"d5", x"d5", x"d5", x"d7", x"dc", x"d4", x"d1", x"d3", x"d4", 
        x"d4", x"d2", x"ce", x"e3", x"f2", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ee", x"ef", x"f1", x"f1", x"e6", 
        x"ed", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ee", x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f2", x"f2", x"f1", x"ef", x"ee", 
        x"ed", x"ec", x"eb", x"ea", x"e8", x"e6", x"e3", x"dc", x"d5", x"d4", x"d0", x"d0", x"cb", x"ca", x"bc", 
        x"ba", x"b5", x"aa", x"9f", x"93", x"8c", x"80", x"70", x"65", x"5c", x"4f", x"44", x"4a", x"55", x"57", 
        x"5d", x"66", x"68", x"67", x"67", x"6c", x"6d", x"78", x"7e", x"7c", x"7d", x"78", x"70", x"62", x"61", 
        x"60", x"5f", x"5f", x"5e", x"5b", x"59", x"5b", x"5c", x"55", x"4c", x"48", x"42", x"37", x"3b", x"46", 
        x"53", x"5d", x"67", x"6a", x"6e", x"6d", x"68", x"67", x"68", x"69", x"67", x"65", x"67", x"68", x"6a", 
        x"6c", x"6d", x"6d", x"6e", x"6f", x"70", x"6a", x"48", x"25", x"18", x"5c", x"ae", x"d7", x"e2", x"df", 
        x"ef", x"f5", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f4", x"f5", x"f5", 
        x"f3", x"f3", x"f6", x"f8", x"f6", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f5", x"f2", x"ef", x"f3", x"f4", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"ef", x"f1", x"f0", x"f2", x"f6", x"f5", x"f4", x"f6", 
        x"f6", x"f5", x"f0", x"af", x"46", x"53", x"92", x"d8", x"d1", x"d3", x"d8", x"d8", x"b8", x"9b", x"a5", 
        x"a3", x"99", x"95", x"94", x"91", x"8c", x"7f", x"75", x"6f", x"6c", x"6f", x"7a", x"81", x"87", x"8f", 
        x"96", x"98", x"97", x"95", x"96", x"96", x"97", x"93", x"58", x"42", x"57", x"83", x"8a", x"8b", x"87", 
        x"86", x"86", x"89", x"89", x"78", x"73", x"72", x"73", x"75", x"78", x"82", x"86", x"84", x"84", x"86", 
        x"85", x"86", x"83", x"81", x"7f", x"80", x"82", x"7f", x"80", x"7e", x"56", x"42", x"3a", x"7b", x"81", 
        x"80", x"81", x"81", x"7f", x"7e", x"7e", x"7d", x"7c", x"7c", x"7c", x"7c", x"7c", x"7d", x"7b", x"7c", 
        x"7c", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7d", x"7c", x"75", x"7c", x"7d", x"78", x"7a", 
        x"80", x"62", x"46", x"76", x"a4", x"af", x"aa", x"a8", x"a4", x"a4", x"9f", x"9f", x"9b", x"8c", x"78", 
        x"77", x"79", x"7c", x"76", x"74", x"73", x"72", x"8c", x"97", x"91", x"8f", x"8e", x"8e", x"8d", x"8d", 
        x"8e", x"8c", x"8b", x"8b", x"8b", x"8b", x"8d", x"7d", x"37", x"4f", x"72", x"6c", x"74", x"7e", x"7b", 
        x"9e", x"aa", x"c1", x"cc", x"c6", x"94", x"a1", x"a3", x"a2", x"c5", x"da", x"f0", x"ec", x"df", x"e1", 
        x"e1", x"d7", x"e5", x"df", x"e8", x"e5", x"eb", x"ef", x"eb", x"e7", x"de", x"cf", x"ce", x"b9", x"82", 
        x"6c", x"83", x"9d", x"9d", x"9b", x"8d", x"9e", x"a1", x"a7", x"a8", x"8d", x"95", x"96", x"84", x"57", 
        x"54", x"79", x"a9", x"aa", x"ac", x"ab", x"aa", x"ad", x"ad", x"9f", x"93", x"8a", x"92", x"99", x"a0", 
        x"ab", x"a8", x"ab", x"ae", x"aa", x"ab", x"ab", x"aa", x"a9", x"a9", x"a9", x"a9", x"aa", x"ad", x"ab", 
        x"aa", x"ab", x"ad", x"aa", x"aa", x"aa", x"aa", x"aa", x"aa", x"ab", x"ac", x"ac", x"ac", x"ab", x"ab", 
        x"ab", x"ab", x"ac", x"ac", x"ac", x"ac", x"ac", x"ab", x"aa", x"aa", x"ac", x"ae", x"aa", x"ac", x"ab", 
        x"ad", x"ae", x"a5", x"75", x"7f", x"a3", x"aa", x"ac", x"ac", x"ab", x"ac", x"ac", x"ab", x"ab", x"ab", 
        x"ab", x"ab", x"ad", x"ae", x"a6", x"aa", x"ab", x"66", x"63", x"7a", x"73", x"74", x"a1", x"ac", x"a8", 
        x"ab", x"ac", x"ad", x"b1", x"a0", x"82", x"80", x"80", x"7f", x"7c", x"7d", x"7e", x"7e", x"7e", x"7c", 
        x"7b", x"75", x"99", x"dd", x"d8", x"d5", x"d5", x"d5", x"dc", x"d9", x"cf", x"d1", x"d0", x"d0", x"d2", 
        x"d1", x"d1", x"d4", x"d5", x"d4", x"d4", x"d4", x"d3", x"d2", x"d3", x"d2", x"d3", x"d4", x"d4", x"d1", 
        x"ce", x"d1", x"d3", x"d0", x"d0", x"d4", x"d3", x"d2", x"d4", x"d3", x"d3", x"d5", x"d5", x"d3", x"d3", 
        x"d6", x"d7", x"d5", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", x"d6", x"db", x"d4", x"d1", x"d3", x"d4", 
        x"d4", x"d1", x"cf", x"e3", x"f3", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"e7", 
        x"ee", x"f2", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ef", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", 
        x"ed", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"ef", x"f0", x"ed", x"ec", x"e9", x"e7", x"dd", 
        x"da", x"d5", x"cd", x"ca", x"ca", x"cb", x"c7", x"c6", x"bb", x"b3", x"a9", x"9a", x"92", x"83", x"6f", 
        x"63", x"5a", x"51", x"4b", x"4b", x"4e", x"4f", x"55", x"5a", x"59", x"61", x"6c", x"69", x"69", x"63", 
        x"57", x"4b", x"45", x"44", x"41", x"3e", x"3f", x"40", x"3b", x"3b", x"45", x"51", x"5e", x"64", x"6e", 
        x"6d", x"67", x"63", x"62", x"63", x"64", x"65", x"65", x"67", x"69", x"69", x"69", x"67", x"67", x"69", 
        x"69", x"68", x"6b", x"71", x"76", x"76", x"76", x"6a", x"52", x"48", x"9a", x"df", x"df", x"da", x"e0", 
        x"f0", x"f0", x"f1", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f4", x"f6", x"f7", x"f6", 
        x"f3", x"f3", x"f6", x"f7", x"f5", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f0", x"ee", x"f2", x"f4", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"ef", x"f1", x"f0", x"f2", x"f6", x"f5", x"f2", x"f4", 
        x"f6", x"f3", x"f2", x"b7", x"48", x"4c", x"83", x"d9", x"d6", x"cf", x"d6", x"d2", x"b3", x"93", x"9d", 
        x"9a", x"95", x"9a", x"9a", x"98", x"99", x"98", x"98", x"97", x"92", x"8d", x"81", x"74", x"68", x"62", 
        x"6a", x"77", x"82", x"8d", x"94", x"96", x"96", x"92", x"5c", x"46", x"55", x"7c", x"85", x"8b", x"89", 
        x"87", x"84", x"87", x"87", x"78", x"74", x"75", x"76", x"77", x"79", x"81", x"85", x"86", x"89", x"8b", 
        x"87", x"88", x"84", x"81", x"82", x"82", x"82", x"7e", x"7d", x"7f", x"56", x"50", x"3d", x"77", x"7e", 
        x"7d", x"7f", x"7f", x"7f", x"7e", x"7e", x"7d", x"7c", x"7c", x"7b", x"7b", x"7d", x"7e", x"7c", x"7c", 
        x"7e", x"7d", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7b", x"75", x"7c", x"7e", x"79", x"7a", 
        x"80", x"69", x"45", x"72", x"a0", x"ae", x"a9", x"a6", x"9f", x"a1", x"a2", x"a0", x"9b", x"8e", x"79", 
        x"7a", x"7a", x"7b", x"73", x"70", x"71", x"75", x"8c", x"99", x"94", x"92", x"8f", x"8f", x"8d", x"8e", 
        x"8d", x"8d", x"8c", x"8a", x"8b", x"8e", x"90", x"85", x"41", x"50", x"7a", x"77", x"7d", x"80", x"7a", 
        x"90", x"87", x"93", x"95", x"b0", x"a3", x"86", x"8c", x"a3", x"d0", x"dc", x"e8", x"e3", x"e6", x"e8", 
        x"ec", x"df", x"e0", x"d3", x"e3", x"e3", x"e7", x"ea", x"e8", x"eb", x"ea", x"eb", x"f0", x"ee", x"db", 
        x"b3", x"aa", x"b7", x"b1", x"b0", x"a5", x"96", x"88", x"83", x"94", x"8d", x"92", x"8b", x"73", x"7e", 
        x"8a", x"93", x"a7", x"a8", x"a9", x"aa", x"ab", x"ab", x"a1", x"8e", x"8a", x"95", x"9d", x"99", x"9d", 
        x"aa", x"a3", x"a3", x"aa", x"aa", x"ab", x"ab", x"ac", x"ab", x"aa", x"aa", x"a9", x"ab", x"ad", x"ab", 
        x"aa", x"ab", x"ad", x"ab", x"ab", x"ab", x"aa", x"aa", x"ab", x"ac", x"ad", x"ad", x"ac", x"ac", x"ab", 
        x"ab", x"ac", x"ad", x"ad", x"ad", x"ac", x"ac", x"ab", x"aa", x"aa", x"ac", x"ad", x"aa", x"ac", x"ac", 
        x"ad", x"ad", x"a5", x"75", x"7e", x"a0", x"aa", x"ad", x"ad", x"ac", x"ac", x"ac", x"ab", x"ab", x"ab", 
        x"ab", x"ab", x"ae", x"af", x"a8", x"aa", x"ab", x"66", x"60", x"7a", x"73", x"74", x"a2", x"ae", x"aa", 
        x"ac", x"ad", x"ad", x"b1", x"a2", x"82", x"81", x"80", x"7e", x"7d", x"7c", x"7d", x"7f", x"7f", x"7d", 
        x"7a", x"74", x"99", x"dd", x"d8", x"d4", x"d5", x"d5", x"da", x"da", x"d1", x"d1", x"cf", x"cf", x"d2", 
        x"ce", x"cd", x"d2", x"d4", x"d5", x"d3", x"d3", x"d1", x"d2", x"d3", x"d3", x"d3", x"d4", x"d3", x"d0", 
        x"cf", x"d1", x"d3", x"cf", x"cf", x"d4", x"d3", x"d2", x"d3", x"d3", x"d3", x"d4", x"d4", x"d2", x"d2", 
        x"d4", x"d6", x"d6", x"d3", x"d3", x"d4", x"d5", x"d5", x"d4", x"d5", x"da", x"d4", x"d3", x"d6", x"d4", 
        x"d2", x"d0", x"d1", x"e5", x"f2", x"ed", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"e8", 
        x"ee", x"f2", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f3", x"f2", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f3", x"f0", x"f1", x"f1", x"f0", x"ee", 
        x"ef", x"f0", x"ed", x"ea", x"e8", x"e4", x"df", x"db", x"d0", x"ca", x"cb", x"cc", x"ce", x"ca", x"c7", 
        x"bf", x"b8", x"af", x"a0", x"93", x"86", x"77", x"68", x"5d", x"54", x"53", x"56", x"4b", x"60", x"5c", 
        x"54", x"53", x"54", x"57", x"53", x"4c", x"4a", x"52", x"56", x"5b", x"62", x"69", x"64", x"5a", x"62", 
        x"65", x"64", x"63", x"63", x"63", x"65", x"69", x"6b", x"69", x"67", x"69", x"6c", x"6b", x"6b", x"6c", 
        x"6c", x"6b", x"6d", x"71", x"73", x"74", x"89", x"7e", x"54", x"4e", x"a2", x"e5", x"df", x"de", x"e2", 
        x"ef", x"f4", x"f3", x"f3", x"f2", x"f1", x"f2", x"f4", x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f4", x"f3", x"f2", x"f4", x"f7", x"f9", x"f6", 
        x"f3", x"f3", x"f6", x"f6", x"f3", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f2", x"f1", x"ef", x"ed", x"f1", x"f2", x"ef", x"f0", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"ef", x"f1", x"f0", x"f2", x"f6", x"f6", x"f3", x"f4", 
        x"f4", x"f2", x"f3", x"bf", x"4e", x"4c", x"72", x"c6", x"d7", x"d1", x"d4", x"d4", x"b9", x"93", x"9b", 
        x"97", x"95", x"98", x"98", x"96", x"94", x"95", x"97", x"98", x"98", x"96", x"96", x"96", x"96", x"93", 
        x"8c", x"80", x"73", x"68", x"68", x"72", x"7c", x"7f", x"57", x"47", x"56", x"7d", x"88", x"8e", x"8d", 
        x"8b", x"87", x"8b", x"8a", x"7b", x"74", x"76", x"76", x"77", x"7b", x"80", x"85", x"86", x"8a", x"8d", 
        x"88", x"86", x"86", x"82", x"82", x"81", x"80", x"7e", x"7e", x"82", x"59", x"5a", x"44", x"79", x"80", 
        x"7e", x"80", x"7f", x"7f", x"7e", x"7e", x"7d", x"7c", x"7b", x"7a", x"7b", x"7d", x"7e", x"7d", x"7e", 
        x"81", x"7f", x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7b", x"7a", x"75", x"7b", x"7d", x"7a", x"79", 
        x"7f", x"6d", x"41", x"6f", x"9f", x"b6", x"b8", x"b9", x"b4", x"a9", x"9e", x"9f", x"99", x"8b", x"76", 
        x"76", x"79", x"7b", x"75", x"71", x"70", x"73", x"89", x"98", x"95", x"93", x"90", x"91", x"8f", x"90", 
        x"8e", x"8d", x"8d", x"8a", x"8b", x"8f", x"8f", x"88", x"44", x"4a", x"7a", x"7a", x"7f", x"8c", x"8a", 
        x"c0", x"bd", x"b4", x"b4", x"bf", x"b5", x"9a", x"a1", x"b0", x"ba", x"c2", x"c9", x"cd", x"c9", x"d1", 
        x"d1", x"c3", x"da", x"e5", x"e7", x"e7", x"e7", x"e8", x"e9", x"ee", x"e8", x"e9", x"e9", x"e7", x"e8", 
        x"e0", x"e2", x"e2", x"e0", x"e0", x"e2", x"df", x"d0", x"b7", x"a9", x"9a", x"87", x"69", x"6d", x"71", 
        x"8b", x"9d", x"a7", x"a1", x"a8", x"aa", x"ab", x"a8", x"a2", x"9b", x"95", x"96", x"97", x"a2", x"9f", 
        x"97", x"96", x"a1", x"a9", x"ab", x"aa", x"ab", x"ac", x"ab", x"ab", x"aa", x"aa", x"ab", x"ab", x"aa", 
        x"aa", x"ab", x"ab", x"ab", x"ab", x"a9", x"a8", x"a8", x"a9", x"aa", x"ab", x"ac", x"ac", x"ac", x"ac", 
        x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ab", x"ab", x"aa", x"ab", x"ad", x"ab", x"ad", x"ab", 
        x"ac", x"ad", x"a6", x"77", x"7e", x"9f", x"a9", x"ad", x"ae", x"ac", x"ac", x"ac", x"ab", x"ab", x"ab", 
        x"ab", x"ab", x"ad", x"ae", x"a9", x"aa", x"ad", x"68", x"60", x"7b", x"75", x"76", x"a4", x"af", x"ab", 
        x"ad", x"ae", x"ac", x"b1", x"a3", x"82", x"81", x"80", x"7e", x"7d", x"7c", x"7b", x"7d", x"7f", x"7d", 
        x"7b", x"74", x"9a", x"de", x"d9", x"d5", x"d5", x"d6", x"da", x"d9", x"d0", x"d1", x"d0", x"d0", x"d2", 
        x"d2", x"d2", x"d2", x"d4", x"d5", x"d3", x"d2", x"d0", x"d1", x"d3", x"d3", x"d3", x"d4", x"d3", x"d1", 
        x"d1", x"d2", x"d4", x"cf", x"cf", x"d3", x"d3", x"d3", x"d5", x"d4", x"d2", x"d3", x"d2", x"d0", x"d1", 
        x"d2", x"d5", x"d5", x"d3", x"d1", x"d3", x"d5", x"d5", x"d4", x"d5", x"d9", x"d3", x"d4", x"d7", x"d4", 
        x"d2", x"d1", x"d1", x"e6", x"f2", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f0", x"f0", x"e8", 
        x"ef", x"f1", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ef", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f2", x"f0", x"f0", x"f2", x"f2", x"f5", 
        x"f4", x"f3", x"f1", x"ef", x"f1", x"f1", x"f2", x"f3", x"f3", x"f5", x"f1", x"ee", x"eb", x"e3", x"dd", 
        x"d3", x"cf", x"d0", x"d5", x"d9", x"d7", x"d4", x"cd", x"c7", x"bc", x"ac", x"a0", x"87", x"79", x"69", 
        x"58", x"57", x"59", x"5c", x"5b", x"5e", x"5a", x"63", x"69", x"6e", x"69", x"62", x"65", x"61", x"63", 
        x"6d", x"6d", x"6b", x"68", x"68", x"6a", x"68", x"67", x"66", x"68", x"6b", x"6d", x"6b", x"6b", x"6c", 
        x"6f", x"73", x"76", x"76", x"75", x"8e", x"ba", x"99", x"51", x"4e", x"9b", x"e5", x"e0", x"db", x"e0", 
        x"ef", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f3", x"f3", x"f5", x"f8", x"f8", x"f6", 
        x"f3", x"f3", x"f5", x"f4", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f2", x"f2", x"f0", x"ed", x"f1", x"f1", x"ee", x"ef", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"ee", x"f0", x"ef", x"f1", x"f0", x"f2", x"f6", x"f8", x"f6", x"f6", 
        x"f2", x"f1", x"f4", x"c5", x"52", x"4c", x"6d", x"af", x"d1", x"db", x"d4", x"d8", x"bd", x"93", x"99", 
        x"96", x"95", x"97", x"96", x"9a", x"96", x"96", x"95", x"94", x"95", x"94", x"91", x"90", x"90", x"92", 
        x"95", x"96", x"96", x"9b", x"95", x"89", x"7c", x"75", x"51", x"41", x"49", x"6a", x"7a", x"81", x"84", 
        x"87", x"86", x"89", x"8a", x"7c", x"75", x"78", x"76", x"75", x"78", x"7e", x"83", x"84", x"88", x"8d", 
        x"89", x"86", x"89", x"83", x"81", x"7f", x"7e", x"7f", x"80", x"80", x"5c", x"59", x"46", x"79", x"81", 
        x"7f", x"7e", x"7b", x"7d", x"7e", x"7e", x"7e", x"7e", x"7e", x"7d", x"7f", x"7f", x"7d", x"7c", x"7c", 
        x"7e", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7b", x"7a", x"75", x"7b", x"7c", x"7b", x"76", 
        x"7e", x"73", x"40", x"6c", x"9e", x"c0", x"c9", x"d3", x"d5", x"c9", x"b4", x"a2", x"98", x"90", x"7b", 
        x"7b", x"7e", x"7c", x"75", x"70", x"6c", x"6f", x"86", x"96", x"94", x"94", x"92", x"93", x"92", x"93", 
        x"90", x"8f", x"8f", x"8d", x"8c", x"8e", x"8d", x"8c", x"48", x"45", x"7b", x"7e", x"81", x"8a", x"89", 
        x"91", x"9a", x"c7", x"eb", x"e1", x"cd", x"d3", x"e1", x"d0", x"a3", x"9e", x"aa", x"a2", x"9a", x"99", 
        x"9f", x"b4", x"c8", x"db", x"dc", x"de", x"df", x"e7", x"e9", x"ec", x"e9", x"e9", x"e9", x"e8", x"eb", 
        x"e5", x"e2", x"e6", x"e8", x"e3", x"ea", x"e8", x"d4", x"dc", x"e3", x"c4", x"9c", x"8d", x"82", x"74", 
        x"92", x"a2", x"a7", x"99", x"9e", x"9e", x"9f", x"a2", x"a5", x"a9", x"a0", x"92", x"95", x"a7", x"9e", 
        x"91", x"90", x"9f", x"a7", x"a9", x"aa", x"ab", x"aa", x"ab", x"aa", x"ab", x"ac", x"ab", x"aa", x"aa", 
        x"ab", x"aa", x"aa", x"ac", x"ac", x"a9", x"a7", x"a8", x"aa", x"ab", x"ab", x"ab", x"ab", x"ac", x"ad", 
        x"ad", x"ac", x"ab", x"ab", x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ab", x"ad", x"aa", 
        x"aa", x"ac", x"a6", x"79", x"7e", x"9f", x"a8", x"ad", x"ad", x"ab", x"ac", x"ac", x"ab", x"ab", x"ab", 
        x"ab", x"ab", x"ab", x"ac", x"a9", x"ab", x"af", x"6a", x"60", x"7c", x"76", x"76", x"a3", x"ae", x"ab", 
        x"ad", x"ad", x"ab", x"b1", x"a3", x"82", x"81", x"81", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", 
        x"7c", x"75", x"9a", x"df", x"d9", x"d5", x"d6", x"d7", x"da", x"d8", x"ce", x"d2", x"d2", x"d1", x"d0", 
        x"d3", x"d3", x"d2", x"d3", x"d5", x"d4", x"d1", x"cf", x"d1", x"d3", x"d3", x"d4", x"d4", x"d3", x"d1", 
        x"d2", x"d3", x"d5", x"d1", x"d0", x"d2", x"d1", x"d2", x"d4", x"d3", x"d2", x"d3", x"d3", x"d1", x"d2", 
        x"d2", x"d4", x"d4", x"d1", x"d1", x"d4", x"d3", x"d4", x"d5", x"d4", x"d5", x"ce", x"cf", x"d4", x"d4", 
        x"d4", x"d2", x"d0", x"e5", x"f3", x"ee", x"ee", x"ed", x"ed", x"ee", x"ee", x"ed", x"ed", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f0", x"ef", x"e9", 
        x"ef", x"f1", x"ef", x"ef", x"f0", x"f0", x"f1", x"f2", x"f2", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f1", x"ee", x"ef", x"f2", x"f2", x"f2", 
        x"ef", x"f0", x"f2", x"ef", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f2", x"f2", x"f2", 
        x"ef", x"ef", x"ec", x"e7", x"e9", x"e7", x"e0", x"dd", x"dc", x"da", x"d8", x"dc", x"d7", x"d8", x"d1", 
        x"c6", x"be", x"ad", x"a0", x"95", x"89", x"7a", x"71", x"64", x"61", x"5f", x"5a", x"58", x"54", x"4f", 
        x"5b", x"5e", x"62", x"67", x"6a", x"6c", x"70", x"6f", x"6e", x"70", x"6d", x"6d", x"71", x"72", x"72", 
        x"76", x"79", x"78", x"79", x"94", x"b2", x"c4", x"9e", x"54", x"4b", x"92", x"e3", x"e1", x"dd", x"e1", 
        x"ed", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", 
        x"f0", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f6", x"f8", x"f8", x"f6", 
        x"f4", x"f4", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f2", x"f3", x"f4", x"f3", x"f4", x"f1", x"f0", x"f3", x"f3", x"ef", x"ef", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"f0", x"ef", x"f1", x"f0", x"f2", x"f6", x"f6", x"f6", x"f6", 
        x"f1", x"f3", x"f7", x"cb", x"56", x"4c", x"76", x"a8", x"bb", x"d6", x"d5", x"d6", x"c0", x"95", x"9c", 
        x"9b", x"9a", x"96", x"95", x"99", x"96", x"96", x"95", x"94", x"99", x"99", x"93", x"92", x"92", x"92", 
        x"91", x"90", x"8f", x"91", x"8d", x"90", x"94", x"94", x"6a", x"45", x"47", x"6c", x"71", x"6c", x"68", 
        x"6c", x"6f", x"73", x"77", x"6c", x"69", x"72", x"75", x"79", x"7e", x"81", x"87", x"86", x"89", x"8f", 
        x"8c", x"87", x"87", x"81", x"83", x"82", x"80", x"80", x"7e", x"80", x"63", x"57", x"45", x"77", x"82", 
        x"7f", x"7d", x"7b", x"7e", x"7f", x"7e", x"7d", x"7e", x"7d", x"7c", x"7f", x"7e", x"7c", x"7c", x"7d", 
        x"7e", x"7d", x"7d", x"7d", x"7d", x"7c", x"7c", x"7c", x"7c", x"7a", x"76", x"7b", x"7c", x"7b", x"75", 
        x"7c", x"78", x"43", x"6e", x"9d", x"be", x"c6", x"ca", x"cf", x"d6", x"d5", x"bb", x"9f", x"91", x"7b", 
        x"77", x"7a", x"78", x"77", x"7a", x"7b", x"7c", x"8a", x"99", x"97", x"94", x"91", x"92", x"91", x"92", 
        x"90", x"90", x"91", x"91", x"93", x"93", x"90", x"91", x"4e", x"43", x"7b", x"7c", x"7b", x"7b", x"7b", 
        x"55", x"7d", x"a7", x"cb", x"cb", x"a8", x"ba", x"e7", x"e6", x"d1", x"d8", x"da", x"c1", x"bb", x"bc", 
        x"bc", x"ba", x"b2", x"b5", x"c5", x"c5", x"c3", x"ce", x"d4", x"e1", x"e9", x"ed", x"ea", x"ec", x"ec", 
        x"e8", x"d7", x"e0", x"dd", x"b5", x"c5", x"ca", x"ab", x"af", x"d9", x"c1", x"9b", x"a9", x"7e", x"91", 
        x"b7", x"ad", x"b4", x"c3", x"ba", x"ad", x"a5", x"9f", x"a2", x"99", x"86", x"88", x"95", x"aa", x"a5", 
        x"a4", x"9f", x"a4", x"aa", x"ac", x"aa", x"a9", x"ac", x"ab", x"aa", x"ab", x"ac", x"ac", x"aa", x"aa", 
        x"ab", x"ab", x"ab", x"ac", x"ad", x"ac", x"ab", x"ac", x"ad", x"ad", x"ad", x"ac", x"ac", x"ac", x"ac", 
        x"ac", x"ac", x"ab", x"ab", x"ac", x"ac", x"ac", x"ab", x"ab", x"ac", x"ac", x"ab", x"ab", x"ad", x"ab", 
        x"aa", x"ac", x"a7", x"79", x"7f", x"a1", x"a9", x"ac", x"ac", x"ab", x"ab", x"ac", x"ac", x"ab", x"aa", 
        x"aa", x"ab", x"ab", x"ac", x"a9", x"ab", x"af", x"6a", x"61", x"7c", x"76", x"75", x"a0", x"ae", x"ac", 
        x"ac", x"ae", x"ac", x"b1", x"a4", x"82", x"81", x"80", x"7d", x"7c", x"7c", x"7b", x"7d", x"7c", x"7c", 
        x"7e", x"75", x"99", x"dd", x"d8", x"d5", x"d7", x"d6", x"d9", x"d7", x"cd", x"d2", x"d4", x"d2", x"d0", 
        x"d2", x"d1", x"d0", x"d3", x"d5", x"d4", x"d1", x"cf", x"d0", x"d3", x"d4", x"d5", x"d4", x"d2", x"d1", 
        x"d1", x"d4", x"d6", x"d2", x"d1", x"d1", x"d1", x"d1", x"d2", x"d4", x"d4", x"d3", x"d3", x"d2", x"d4", 
        x"d3", x"d5", x"d5", x"d2", x"d2", x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"cd", x"cd", x"d3", x"d3", 
        x"d5", x"d2", x"d1", x"e3", x"f4", x"ee", x"ed", x"ec", x"ed", x"ee", x"ee", x"ee", x"ed", x"ef", x"ef", 
        x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f2", x"f2", x"f0", x"ea", 
        x"ee", x"f1", x"ef", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"f0", x"f0", x"ef", x"ee", x"ed", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ef", x"f1", x"f1", x"f2", x"f3", x"f0", x"ee", x"ee", x"f0", x"f1", x"f3", 
        x"f0", x"f1", x"f2", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"ef", x"f1", x"ef", x"ed", x"f1", x"f4", x"f3", x"f2", x"f3", x"f3", x"f1", x"ee", x"e9", x"ea", x"e8", 
        x"e3", x"e3", x"e1", x"e4", x"e8", x"e3", x"db", x"d5", x"c6", x"b8", x"a8", x"95", x"88", x"7c", x"68", 
        x"62", x"5a", x"58", x"59", x"54", x"51", x"57", x"5c", x"62", x"6c", x"6f", x"70", x"75", x"7a", x"81", 
        x"83", x"82", x"8a", x"a0", x"c4", x"c5", x"c8", x"a5", x"58", x"4c", x"8e", x"e2", x"e2", x"e0", x"e0", 
        x"ed", x"f8", x"f2", x"f1", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f6", x"f8", x"f9", x"f7", 
        x"f5", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f0", x"f3", x"f3", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"f0", x"f0", x"f0", x"f0", x"f2", x"f5", x"f6", x"f5", x"f3", 
        x"f2", x"f6", x"f8", x"cf", x"5d", x"4b", x"7a", x"b8", x"a7", x"cc", x"d6", x"d3", x"c2", x"94", x"9a", 
        x"99", x"98", x"97", x"95", x"97", x"97", x"97", x"96", x"96", x"97", x"98", x"97", x"94", x"92", x"90", 
        x"90", x"8f", x"8d", x"90", x"8c", x"8d", x"90", x"93", x"68", x"3f", x"4a", x"7a", x"8d", x"8e", x"89", 
        x"83", x"77", x"6f", x"68", x"5b", x"54", x"5a", x"5e", x"62", x"68", x"70", x"7c", x"84", x"8c", x"95", 
        x"92", x"8a", x"87", x"82", x"82", x"83", x"7f", x"7e", x"7d", x"7e", x"67", x"56", x"44", x"78", x"85", 
        x"81", x"81", x"80", x"80", x"7f", x"7f", x"7d", x"7c", x"7a", x"7a", x"7f", x"7d", x"7b", x"7c", x"7e", 
        x"7f", x"7c", x"7d", x"7e", x"7c", x"7c", x"7c", x"7c", x"7c", x"7b", x"78", x"7a", x"7b", x"7b", x"76", 
        x"7d", x"78", x"42", x"6d", x"9d", x"bb", x"c2", x"c8", x"ca", x"d1", x"d7", x"d4", x"b5", x"92", x"79", 
        x"7c", x"80", x"7f", x"7e", x"7d", x"7b", x"7a", x"89", x"9a", x"95", x"95", x"95", x"94", x"92", x"94", 
        x"92", x"91", x"8e", x"8a", x"89", x"85", x"80", x"86", x"4c", x"3f", x"7b", x"80", x"80", x"7d", x"7b", 
        x"75", x"8a", x"6c", x"75", x"86", x"72", x"7a", x"a0", x"ba", x"cb", x"e1", x"eb", x"e3", x"d5", x"e7", 
        x"ec", x"ec", x"e1", x"c7", x"d5", x"d6", x"d0", x"ca", x"bf", x"b0", x"9f", x"be", x"d1", x"da", x"e4", 
        x"e6", x"e2", x"e9", x"dd", x"b3", x"a4", x"97", x"95", x"9f", x"c2", x"bf", x"7e", x"89", x"7d", x"82", 
        x"91", x"a2", x"b5", x"ee", x"f0", x"e7", x"e3", x"d0", x"d3", x"c5", x"ad", x"a4", x"93", x"87", x"7c", 
        x"88", x"92", x"9d", x"a4", x"ac", x"ac", x"ab", x"af", x"ad", x"ab", x"ad", x"ad", x"ad", x"ac", x"ab", 
        x"ab", x"ab", x"ab", x"ab", x"ad", x"ac", x"ab", x"aa", x"ac", x"ae", x"af", x"ab", x"ab", x"ac", x"ad", 
        x"ac", x"ac", x"ac", x"ac", x"ac", x"ac", x"ab", x"aa", x"aa", x"ac", x"ac", x"ac", x"ac", x"ad", x"ac", 
        x"ab", x"ad", x"a7", x"79", x"7e", x"a5", x"aa", x"ad", x"ad", x"ac", x"aa", x"ac", x"ac", x"ab", x"a9", 
        x"aa", x"ac", x"ad", x"ad", x"a8", x"ab", x"ac", x"67", x"61", x"7c", x"75", x"74", x"9c", x"ae", x"ad", 
        x"ac", x"ae", x"ae", x"b0", x"a2", x"7e", x"80", x"81", x"80", x"7b", x"7b", x"7a", x"7d", x"7d", x"7b", 
        x"7d", x"74", x"97", x"dd", x"da", x"d6", x"d8", x"d4", x"d7", x"d5", x"cd", x"d1", x"d1", x"d1", x"d0", 
        x"d2", x"d2", x"d1", x"d3", x"d4", x"d5", x"d4", x"d1", x"d0", x"d1", x"d3", x"d5", x"d4", x"d1", x"cf", 
        x"d0", x"d2", x"d3", x"d3", x"d4", x"d2", x"d2", x"d0", x"d1", x"d7", x"d6", x"d1", x"d2", x"d2", x"d2", 
        x"d4", x"d5", x"d5", x"d5", x"d4", x"d2", x"d4", x"d1", x"d2", x"d5", x"d6", x"d2", x"d2", x"d6", x"d4", 
        x"d4", x"d2", x"d2", x"e2", x"f5", x"ed", x"ed", x"ed", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f0", x"ef", x"ed", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f3", x"f2", x"eb", 
        x"eb", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"f2", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"ee", x"ee", x"f0", x"ed", x"ea", x"eb", x"ed", x"ec", x"e9", x"e8", x"e5", x"dd", 
        x"d3", x"ca", x"bf", x"b0", x"a3", x"97", x"8a", x"7d", x"70", x"65", x"5b", x"52", x"49", x"48", x"52", 
        x"57", x"5d", x"73", x"91", x"9a", x"a8", x"b8", x"a8", x"6b", x"59", x"8c", x"e1", x"e3", x"e2", x"e1", 
        x"eb", x"f4", x"f2", x"f0", x"f3", x"f1", x"f1", x"f1", x"f3", x"f3", x"f1", x"f1", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", 
        x"f2", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f5", x"f5", x"f6", x"f7", x"f9", x"f7", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f4", x"f4", x"f3", x"f1", x"f1", x"f0", x"f3", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"ef", x"f0", x"f2", x"f3", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f2", x"f4", x"f7", x"f5", x"f1", 
        x"f6", x"f7", x"f7", x"d2", x"64", x"4a", x"6f", x"ce", x"ae", x"ad", x"d9", x"d6", x"c6", x"96", x"9d", 
        x"9d", x"96", x"9a", x"97", x"93", x"96", x"93", x"93", x"95", x"95", x"98", x"98", x"93", x"90", x"90", 
        x"92", x"92", x"8f", x"8e", x"8e", x"8e", x"8b", x"92", x"6a", x"41", x"4a", x"6e", x"82", x"85", x"87", 
        x"8a", x"8b", x"8d", x"8b", x"7d", x"70", x"6d", x"68", x"63", x"5f", x"59", x"57", x"58", x"5e", x"6f", 
        x"78", x"7c", x"84", x"88", x"8c", x"90", x"8a", x"84", x"7f", x"81", x"69", x"50", x"40", x"76", x"86", 
        x"7c", x"7e", x"80", x"7d", x"7e", x"7f", x"7f", x"7e", x"7a", x"7b", x"80", x"7d", x"7c", x"7c", x"7b", 
        x"7d", x"79", x"79", x"7b", x"7e", x"7e", x"7d", x"7b", x"7a", x"7a", x"79", x"7a", x"78", x"7b", x"77", 
        x"7c", x"7c", x"45", x"68", x"98", x"b9", x"c3", x"ca", x"cc", x"d4", x"d2", x"da", x"d4", x"a5", x"7b", 
        x"7e", x"7e", x"7a", x"7b", x"7a", x"7b", x"7b", x"87", x"99", x"94", x"95", x"93", x"94", x"93", x"95", 
        x"96", x"94", x"86", x"79", x"7d", x"80", x"7f", x"82", x"57", x"3c", x"66", x"6c", x"64", x"55", x"56", 
        x"7b", x"8b", x"81", x"7a", x"8e", x"75", x"6d", x"8a", x"90", x"8a", x"8c", x"95", x"9c", x"9e", x"ba", 
        x"c3", x"da", x"e0", x"df", x"df", x"e8", x"ea", x"e9", x"dd", x"ac", x"75", x"a4", x"d1", x"ca", x"b4", 
        x"c6", x"d0", x"c7", x"c8", x"c0", x"c1", x"a8", x"9d", x"a8", x"bf", x"ba", x"92", x"9c", x"96", x"9d", 
        x"9b", x"b3", x"ba", x"de", x"d9", x"da", x"e1", x"e1", x"ed", x"ed", x"e3", x"b9", x"86", x"80", x"83", 
        x"96", x"99", x"97", x"9d", x"9e", x"99", x"9a", x"a3", x"a6", x"a7", x"ab", x"ad", x"ae", x"ac", x"a9", 
        x"a9", x"aa", x"ab", x"ab", x"aa", x"a9", x"aa", x"ab", x"ae", x"ad", x"ab", x"ab", x"ac", x"ac", x"ac", 
        x"ab", x"ab", x"ac", x"ad", x"ac", x"ac", x"ac", x"ac", x"ad", x"ad", x"ac", x"ab", x"ac", x"ac", x"ad", 
        x"ac", x"ae", x"a8", x"79", x"7e", x"a4", x"ab", x"ad", x"ad", x"ac", x"ab", x"ab", x"ab", x"aa", x"aa", 
        x"ab", x"ac", x"ab", x"ac", x"a8", x"ab", x"ad", x"66", x"60", x"7d", x"77", x"75", x"9c", x"ad", x"ad", 
        x"ac", x"af", x"af", x"b1", x"a4", x"7f", x"7d", x"7d", x"7e", x"7c", x"7d", x"7b", x"7c", x"7d", x"7c", 
        x"7d", x"73", x"98", x"dc", x"d8", x"d5", x"d6", x"d5", x"d9", x"d5", x"cf", x"d3", x"d1", x"d2", x"d2", 
        x"d3", x"d2", x"d3", x"d3", x"d3", x"d3", x"d3", x"d1", x"cf", x"d0", x"d1", x"d3", x"d2", x"d1", x"d1", 
        x"d1", x"d0", x"d2", x"d4", x"d7", x"d2", x"d1", x"d2", x"d1", x"d6", x"d4", x"d2", x"d2", x"d3", x"d3", 
        x"d4", x"d4", x"d4", x"d3", x"d2", x"d1", x"d3", x"d2", x"d3", x"d4", x"d6", x"d4", x"d2", x"d7", x"d6", 
        x"d6", x"d3", x"d3", x"e3", x"f5", x"ed", x"ed", x"ed", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"ea", 
        x"eb", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", 
        x"ef", x"ee", x"ed", x"e7", x"e4", x"e3", x"dd", x"d5", x"ca", x"bc", x"ae", x"a3", x"96", x"8a", x"7f", 
        x"76", x"6b", x"63", x"5a", x"4d", x"4d", x"52", x"60", x"5c", x"5a", x"84", x"df", x"e7", x"e1", x"df", 
        x"ea", x"f3", x"f2", x"ef", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f3", x"f2", x"f3", x"f1", x"f1", 
        x"f3", x"f2", x"f3", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f3", x"f3", x"f2", x"f2", 
        x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f5", x"f6", x"f5", x"f6", x"f7", x"f8", x"f6", 
        x"f5", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f0", x"f3", x"ef", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f2", x"f4", x"f4", x"f3", x"f2", 
        x"f6", x"f6", x"f8", x"d6", x"6a", x"4b", x"68", x"d0", x"ca", x"94", x"cc", x"da", x"c6", x"96", x"9b", 
        x"9d", x"97", x"96", x"98", x"95", x"97", x"95", x"94", x"95", x"94", x"96", x"95", x"92", x"90", x"90", 
        x"91", x"91", x"90", x"8f", x"8e", x"8e", x"8d", x"93", x"70", x"48", x"50", x"72", x"83", x"85", x"86", 
        x"86", x"84", x"85", x"87", x"7e", x"75", x"77", x"77", x"75", x"74", x"73", x"70", x"6d", x"70", x"73", 
        x"67", x"5c", x"63", x"66", x"68", x"71", x"77", x"7c", x"80", x"87", x"6f", x"50", x"40", x"71", x"87", 
        x"7d", x"7c", x"7d", x"7d", x"7d", x"7e", x"7e", x"7d", x"7c", x"7f", x"80", x"7d", x"7c", x"7d", x"7c", 
        x"7d", x"7d", x"7b", x"7b", x"7d", x"7f", x"7f", x"7b", x"79", x"79", x"79", x"7b", x"7a", x"7c", x"76", 
        x"79", x"7e", x"49", x"62", x"95", x"b9", x"c4", x"c8", x"cd", x"d2", x"d3", x"d5", x"db", x"be", x"80", 
        x"7b", x"7d", x"7b", x"7d", x"7b", x"7b", x"7a", x"86", x"98", x"93", x"99", x"9a", x"9a", x"9c", x"9b", 
        x"9a", x"99", x"87", x"70", x"6b", x"69", x"65", x"5b", x"40", x"2d", x"54", x"62", x"62", x"5d", x"63", 
        x"77", x"70", x"81", x"a3", x"ab", x"8f", x"8b", x"a9", x"a0", x"8d", x"7f", x"7c", x"7c", x"85", x"77", 
        x"7a", x"96", x"96", x"98", x"94", x"b9", x"d9", x"eb", x"f2", x"e1", x"ce", x"dc", x"dc", x"be", x"a7", 
        x"d0", x"d1", x"9f", x"ac", x"be", x"aa", x"9a", x"a8", x"ac", x"b0", x"ab", x"ad", x"a0", x"93", x"c2", 
        x"af", x"ac", x"bb", x"be", x"b8", x"bd", x"d5", x"c4", x"cf", x"e9", x"f1", x"c8", x"95", x"8a", x"9e", 
        x"c8", x"db", x"db", x"d4", x"c9", x"c0", x"b3", x"a5", x"9b", x"97", x"9a", x"9a", x"9e", x"a3", x"aa", 
        x"af", x"b1", x"ad", x"ab", x"ad", x"ac", x"ab", x"ab", x"ac", x"ad", x"ad", x"aa", x"ab", x"ab", x"aa", 
        x"a9", x"a9", x"ab", x"ae", x"ae", x"ab", x"ab", x"ac", x"ad", x"ac", x"ab", x"ab", x"ab", x"ac", x"ad", 
        x"ac", x"af", x"a9", x"7a", x"7d", x"a4", x"ab", x"ad", x"ae", x"ad", x"ad", x"ab", x"aa", x"aa", x"ab", 
        x"ac", x"ac", x"aa", x"ab", x"a9", x"ac", x"ad", x"65", x"5d", x"7d", x"78", x"75", x"9c", x"ad", x"ad", 
        x"ad", x"b0", x"ae", x"ae", x"a3", x"81", x"7f", x"7d", x"7b", x"7a", x"7f", x"80", x"7e", x"7f", x"80", 
        x"80", x"78", x"9b", x"dd", x"d7", x"d7", x"d5", x"d3", x"db", x"d8", x"d1", x"d4", x"d2", x"d1", x"d4", 
        x"d4", x"d3", x"d4", x"d3", x"d2", x"d2", x"d3", x"d2", x"d0", x"cf", x"d0", x"d1", x"d1", x"d1", x"d3", 
        x"d4", x"d1", x"d1", x"d4", x"d6", x"d0", x"ce", x"d2", x"d0", x"d4", x"d3", x"d1", x"d3", x"d4", x"d5", 
        x"d5", x"d4", x"d3", x"d2", x"d2", x"d1", x"d2", x"d3", x"d4", x"d3", x"d6", x"d5", x"d2", x"d7", x"d6", 
        x"d6", x"d3", x"d3", x"e2", x"f4", x"ed", x"ed", x"ed", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"ea", 
        x"ea", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ef", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"ee", x"f1", x"f3", x"f2", x"f0", x"f0", x"f2", x"f2", x"f3", x"f3", 
        x"f0", x"f1", x"f1", x"ee", x"ef", x"f1", x"f0", x"ee", x"ed", x"eb", x"e7", x"e4", x"e4", x"e1", x"db", 
        x"d7", x"d1", x"c1", x"b0", x"a4", x"96", x"84", x"7b", x"75", x"65", x"80", x"db", x"e7", x"e2", x"e2", 
        x"ed", x"f6", x"f3", x"f0", x"f2", x"f0", x"f2", x"f4", x"f4", x"f2", x"ef", x"ee", x"f2", x"f1", x"f2", 
        x"f3", x"f0", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f1", x"f4", x"f4", x"f4", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f5", x"f6", x"f5", x"f6", x"f7", x"f8", x"f6", 
        x"f4", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"ef", x"ef", x"f0", x"f2", x"f1", 
        x"f1", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f0", x"f3", x"ee", x"f1", x"f3", x"f3", x"f2", x"f2", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f4", x"f3", x"f2", x"f3", 
        x"f5", x"f5", x"f8", x"da", x"6e", x"4a", x"67", x"cf", x"db", x"a5", x"ae", x"e0", x"c9", x"98", x"9a", 
        x"9c", x"9a", x"98", x"97", x"95", x"97", x"97", x"96", x"96", x"95", x"96", x"93", x"91", x"90", x"90", 
        x"91", x"91", x"91", x"8f", x"8d", x"8e", x"8c", x"90", x"71", x"46", x"50", x"74", x"85", x"87", x"8b", 
        x"89", x"88", x"89", x"89", x"81", x"77", x"76", x"77", x"75", x"73", x"77", x"77", x"78", x"84", x"93", 
        x"8c", x"81", x"86", x"82", x"71", x"62", x"5b", x"55", x"50", x"5e", x"58", x"4b", x"49", x"6f", x"89", 
        x"83", x"80", x"7e", x"7e", x"7e", x"7d", x"7d", x"7d", x"7d", x"7b", x"7c", x"7b", x"7e", x"7f", x"7d", 
        x"7c", x"7c", x"7b", x"79", x"7a", x"7b", x"7d", x"7c", x"79", x"78", x"78", x"7b", x"7c", x"7d", x"76", 
        x"7a", x"7e", x"49", x"5f", x"97", x"b8", x"c2", x"c7", x"cc", x"cf", x"d6", x"d3", x"dc", x"ca", x"84", 
        x"78", x"7b", x"7b", x"7e", x"7f", x"81", x"82", x"8e", x"a2", x"9c", x"9f", x"97", x"84", x"7b", x"73", 
        x"67", x"62", x"5b", x"55", x"5e", x"64", x"69", x"6b", x"51", x"39", x"6d", x"7e", x"7f", x"79", x"75", 
        x"89", x"6e", x"86", x"9c", x"9c", x"8b", x"91", x"aa", x"a7", x"9a", x"97", x"99", x"93", x"93", x"7f", 
        x"7f", x"7c", x"75", x"6b", x"63", x"6c", x"69", x"74", x"90", x"a9", x"b2", x"b3", x"bd", x"c8", x"d1", 
        x"e3", x"d9", x"8f", x"94", x"cc", x"9c", x"7d", x"9d", x"b3", x"96", x"9e", x"a0", x"93", x"6c", x"b3", 
        x"cf", x"c3", x"ba", x"aa", x"b6", x"a9", x"c9", x"bc", x"db", x"ec", x"e4", x"e2", x"c3", x"c8", x"d2", 
        x"da", x"dc", x"cc", x"d8", x"ea", x"eb", x"ea", x"e8", x"e0", x"d6", x"cb", x"bc", x"ac", x"a5", x"9d", 
        x"9b", x"9d", x"a2", x"a5", x"a8", x"ab", x"ac", x"ab", x"aa", x"ab", x"ad", x"ae", x"ae", x"ae", x"ac", 
        x"ab", x"aa", x"ac", x"ad", x"ab", x"a9", x"a9", x"ac", x"ac", x"ab", x"ab", x"ab", x"ab", x"ac", x"ad", 
        x"ac", x"af", x"aa", x"7b", x"7c", x"a4", x"ac", x"ae", x"ae", x"ae", x"ae", x"ac", x"aa", x"aa", x"ac", 
        x"ad", x"ac", x"ab", x"ac", x"aa", x"ad", x"ad", x"64", x"5b", x"7b", x"76", x"74", x"9c", x"ae", x"ae", 
        x"af", x"b1", x"ae", x"af", x"a4", x"82", x"81", x"7e", x"7f", x"7f", x"7e", x"7d", x"80", x"86", x"86", 
        x"80", x"6d", x"97", x"e0", x"d6", x"d7", x"d5", x"d4", x"d9", x"d9", x"cc", x"d0", x"d1", x"c9", x"cf", 
        x"d3", x"d3", x"d4", x"d3", x"d2", x"d1", x"d3", x"d3", x"d2", x"d0", x"d0", x"d1", x"d3", x"d2", x"d4", 
        x"d4", x"d4", x"d4", x"d4", x"d4", x"d0", x"d1", x"d3", x"d1", x"d4", x"d3", x"d1", x"d3", x"d4", x"d6", 
        x"d6", x"d5", x"d4", x"d3", x"d3", x"d2", x"d1", x"d4", x"d5", x"d3", x"d7", x"d6", x"d1", x"d6", x"d5", 
        x"d5", x"d2", x"d1", x"e1", x"f3", x"ed", x"ed", x"ed", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ea", 
        x"ea", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"f1", 
        x"ef", x"f0", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"ee", x"ec", x"ed", x"f1", x"f2", x"ef", 
        x"ee", x"ee", x"eb", x"e7", x"e3", x"dd", x"d8", x"d1", x"d1", x"c7", x"ca", x"df", x"e4", x"e5", x"d9", 
        x"d6", x"e7", x"ea", x"ea", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f3", x"f2", 
        x"f2", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f3", x"f6", x"f7", x"f7", x"f7", x"f8", x"f8", x"f6", 
        x"f4", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"ee", x"f1", x"f3", x"f3", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f1", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f6", x"f9", x"dc", x"71", x"48", x"63", x"c9", x"de", x"cf", x"a0", x"c9", x"cf", x"9d", x"9b", 
        x"9b", x"98", x"99", x"96", x"95", x"96", x"98", x"97", x"95", x"96", x"96", x"93", x"92", x"91", x"91", 
        x"90", x"90", x"91", x"8f", x"8d", x"8f", x"8d", x"8f", x"73", x"43", x"4e", x"76", x"87", x"86", x"88", 
        x"87", x"87", x"87", x"86", x"7e", x"73", x"71", x"73", x"74", x"72", x"74", x"75", x"72", x"7a", x"90", 
        x"92", x"87", x"8c", x"92", x"8b", x"85", x"82", x"7c", x"74", x"6d", x"60", x"4d", x"48", x"58", x"6d", 
        x"66", x"70", x"79", x"7d", x"80", x"80", x"7f", x"7d", x"7e", x"7f", x"7c", x"7c", x"7c", x"7d", x"7c", 
        x"7b", x"7d", x"7e", x"7e", x"7d", x"7c", x"7c", x"7c", x"7c", x"7a", x"78", x"7a", x"7a", x"7b", x"74", 
        x"77", x"7c", x"4f", x"5b", x"93", x"b6", x"c4", x"ca", x"d0", x"d3", x"d4", x"d2", x"db", x"cb", x"8d", 
        x"7e", x"81", x"80", x"7e", x"78", x"75", x"6e", x"69", x"70", x"68", x"57", x"5a", x"71", x"7c", x"84", 
        x"88", x"91", x"8d", x"7f", x"7c", x"7b", x"7e", x"83", x"5b", x"31", x"6d", x"80", x"7f", x"7d", x"75", 
        x"7f", x"86", x"a4", x"9d", x"9f", x"96", x"8f", x"a9", x"aa", x"a8", x"a6", x"a0", x"aa", x"a7", x"94", 
        x"8e", x"85", x"83", x"6d", x"79", x"88", x"5d", x"33", x"49", x"63", x"49", x"4e", x"6a", x"8a", x"9b", 
        x"b4", x"c5", x"bf", x"a6", x"b9", x"c8", x"99", x"af", x"d7", x"c8", x"cb", x"ca", x"b0", x"a1", x"b2", 
        x"bf", x"9b", x"90", x"a8", x"b6", x"c0", x"cd", x"bd", x"e3", x"d8", x"c1", x"cc", x"b1", x"bb", x"d0", 
        x"d5", x"cd", x"c0", x"d2", x"e8", x"eb", x"ea", x"eb", x"e9", x"eb", x"ed", x"ea", x"e9", x"e5", x"db", 
        x"cf", x"bf", x"ad", x"a0", x"95", x"99", x"a0", x"a3", x"a4", x"a6", x"a9", x"ac", x"ad", x"ae", x"ae", 
        x"ae", x"ae", x"ad", x"ab", x"a9", x"a8", x"a9", x"ab", x"ac", x"ad", x"ac", x"ab", x"ac", x"ac", x"ad", 
        x"ac", x"af", x"a9", x"7b", x"7b", x"a3", x"ab", x"ad", x"ad", x"ae", x"ae", x"ac", x"ab", x"ab", x"ac", 
        x"ad", x"ac", x"ab", x"ad", x"aa", x"ad", x"ad", x"65", x"5c", x"7a", x"75", x"73", x"9c", x"ae", x"af", 
        x"ae", x"af", x"ae", x"b2", x"a5", x"80", x"83", x"82", x"82", x"81", x"83", x"85", x"7f", x"70", x"5e", 
        x"47", x"2c", x"71", x"da", x"d7", x"d6", x"d3", x"d2", x"d6", x"d7", x"ca", x"cf", x"d1", x"cc", x"d2", 
        x"d4", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", x"d4", x"d3", x"d3", 
        x"d1", x"d4", x"d4", x"d3", x"d4", x"d2", x"d5", x"d4", x"d0", x"d3", x"d3", x"d2", x"d3", x"d3", x"d6", 
        x"d6", x"d6", x"d5", x"d4", x"d3", x"d3", x"d2", x"d4", x"d6", x"d4", x"d8", x"d6", x"d2", x"d5", x"d4", 
        x"d4", x"d2", x"d1", x"e1", x"f3", x"ed", x"ed", x"ed", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"ee", x"ef", x"f0", x"eb", 
        x"eb", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", x"f0", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"ef", x"f0", x"f2", x"f2", x"f1", x"f1", x"f0", x"ef", x"f0", x"f2", x"f3", x"f1", x"ef", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"ea", x"eb", x"e7", x"e0", x"de", x"db", x"d8", x"c6", 
        x"b7", x"bf", x"bd", x"bf", x"cb", x"d2", x"d6", x"da", x"e4", x"ec", x"ee", x"f0", x"f0", x"f1", x"f3", 
        x"f4", x"f6", x"f5", x"f4", x"f4", x"f3", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f4", x"f5", 
        x"f5", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", x"f4", x"f7", x"f8", x"f7", x"f7", x"f8", x"f8", x"f6", 
        x"f4", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"f0", x"f2", 
        x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"ed", x"f0", x"f3", x"f2", x"f0", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"f1", x"f3", x"f5", x"f5", x"f5", 
        x"f4", x"f7", x"f8", x"df", x"78", x"4b", x"5f", x"c4", x"dd", x"da", x"b0", x"a4", x"ca", x"a2", x"9a", 
        x"9c", x"95", x"97", x"97", x"98", x"98", x"98", x"96", x"93", x"94", x"94", x"93", x"92", x"91", x"91", 
        x"90", x"90", x"91", x"8f", x"8d", x"90", x"8e", x"91", x"7a", x"45", x"4e", x"76", x"8a", x"86", x"86", 
        x"84", x"84", x"84", x"85", x"7e", x"71", x"6f", x"72", x"75", x"73", x"73", x"76", x"75", x"78", x"8c", 
        x"91", x"84", x"85", x"8e", x"87", x"7f", x"80", x"81", x"82", x"81", x"74", x"51", x"4b", x"59", x"71", 
        x"62", x"5b", x"53", x"55", x"5b", x"63", x"6e", x"76", x"7b", x"7c", x"7b", x"7d", x"7d", x"7e", x"80", 
        x"80", x"7c", x"7a", x"79", x"79", x"7a", x"7b", x"7a", x"7c", x"7b", x"79", x"79", x"78", x"78", x"72", 
        x"76", x"7b", x"52", x"55", x"90", x"b9", x"c6", x"cb", x"d1", x"d4", x"d2", x"cd", x"c7", x"b2", x"7e", 
        x"67", x"60", x"55", x"50", x"50", x"58", x"5d", x"69", x"85", x"a0", x"7d", x"72", x"9b", x"9b", x"96", 
        x"98", x"9c", x"90", x"80", x"7e", x"7e", x"7f", x"82", x"63", x"34", x"65", x"7a", x"74", x"72", x"68", 
        x"8c", x"9e", x"a4", x"91", x"99", x"92", x"8a", x"aa", x"b0", x"ab", x"a1", x"a8", x"b3", x"a7", x"97", 
        x"8f", x"86", x"84", x"7c", x"84", x"8d", x"6d", x"3f", x"59", x"82", x"61", x"62", x"5a", x"73", x"67", 
        x"51", x"4a", x"99", x"c5", x"a4", x"99", x"a0", x"a1", x"bf", x"ba", x"b2", x"ab", x"a3", x"86", x"81", 
        x"93", x"8d", x"9c", x"a2", x"87", x"a3", x"b5", x"a1", x"b5", x"bc", x"b5", x"af", x"9d", x"cc", x"e6", 
        x"df", x"d2", x"c6", x"d7", x"e4", x"eb", x"ed", x"ed", x"e9", x"eb", x"ee", x"eb", x"ec", x"ec", x"ec", 
        x"ec", x"ea", x"e5", x"e1", x"d8", x"cf", x"c3", x"b7", x"ac", x"a4", x"a0", x"a2", x"a2", x"a1", x"a3", 
        x"a7", x"a9", x"aa", x"ab", x"ac", x"ab", x"ab", x"ab", x"ab", x"ac", x"ac", x"ac", x"ac", x"ad", x"ac", 
        x"ab", x"ae", x"a9", x"7c", x"7a", x"a2", x"ac", x"ad", x"ac", x"ad", x"ad", x"ac", x"ac", x"ac", x"ac", 
        x"ad", x"ac", x"ab", x"ac", x"aa", x"ad", x"ae", x"67", x"5f", x"7b", x"75", x"74", x"9d", x"ae", x"ad", 
        x"ac", x"ae", x"ae", x"b2", x"a6", x"86", x"8b", x"84", x"7e", x"76", x"68", x"56", x"3e", x"2e", x"29", 
        x"24", x"1f", x"6e", x"e1", x"d8", x"d4", x"d5", x"d6", x"d8", x"d5", x"cc", x"d0", x"d1", x"d5", x"d5", 
        x"d3", x"d1", x"d1", x"d1", x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d4", x"d4", x"d3", x"d2", 
        x"d1", x"d3", x"d4", x"d5", x"d6", x"d4", x"d5", x"d4", x"d0", x"d4", x"d4", x"d3", x"d4", x"d3", x"d3", 
        x"d4", x"d5", x"d5", x"d4", x"d3", x"d2", x"d2", x"d4", x"d6", x"d5", x"d9", x"d6", x"d2", x"d5", x"d4", 
        x"d4", x"d2", x"d2", x"e2", x"f4", x"ed", x"ed", x"ed", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", x"f2", x"ef", x"ef", x"f1", x"ec", 
        x"ec", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"ef", x"f0", x"f3", x"f1", x"f0", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", 
        x"f1", x"f2", x"f2", x"f3", x"f2", x"f3", x"f3", x"f0", x"f1", x"f3", x"f1", x"f0", x"ee", x"ef", x"eb", 
        x"e4", x"e5", x"de", x"d0", x"cd", x"c5", x"c0", x"be", x"c1", x"c3", x"c6", x"cd", x"cc", x"d3", x"da", 
        x"de", x"e6", x"e5", x"e9", x"ee", x"f1", x"f2", x"f2", x"f2", x"f3", x"f5", x"f4", x"f3", x"f4", x"f4", 
        x"f3", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f2", x"f2", x"f3", x"f4", x"f4", 
        x"f2", x"f1", x"f3", x"f4", x"f3", x"f1", x"f2", x"f4", x"f7", x"f8", x"f7", x"f7", x"f8", x"f8", x"f6", 
        x"f3", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f3", 
        x"f3", x"f1", x"f1", x"f0", x"f0", x"ef", x"f2", x"f4", x"f3", x"ed", x"f0", x"f2", x"f1", x"ef", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", x"f0", x"f2", x"f4", x"f5", x"f5", 
        x"f5", x"f6", x"f7", x"e2", x"7f", x"4c", x"5e", x"c0", x"db", x"d5", x"ca", x"9f", x"b8", x"a6", x"99", 
        x"9c", x"97", x"98", x"98", x"97", x"95", x"97", x"96", x"93", x"96", x"97", x"95", x"93", x"92", x"91", 
        x"91", x"91", x"90", x"90", x"8f", x"8f", x"8e", x"91", x"7e", x"47", x"4b", x"73", x"8c", x"87", x"87", 
        x"86", x"86", x"84", x"86", x"80", x"73", x"6f", x"72", x"74", x"72", x"72", x"74", x"75", x"75", x"85", 
        x"90", x"87", x"84", x"91", x"8d", x"83", x"81", x"7d", x"7d", x"81", x"79", x"4d", x"48", x"60", x"8b", 
        x"7f", x"7e", x"7a", x"77", x"73", x"6e", x"64", x"5b", x"59", x"5e", x"63", x"6c", x"6f", x"73", x"79", 
        x"7d", x"7c", x"7e", x"7e", x"7d", x"7c", x"7b", x"7b", x"7a", x"7b", x"7c", x"7e", x"7d", x"7f", x"7a", 
        x"7e", x"7f", x"59", x"55", x"89", x"aa", x"b3", x"b1", x"a9", x"9f", x"97", x"91", x"92", x"8e", x"6d", 
        x"62", x"6e", x"77", x"7e", x"80", x"81", x"7e", x"80", x"95", x"a9", x"82", x"6c", x"9a", x"9b", x"99", 
        x"9a", x"9b", x"8f", x"7e", x"79", x"73", x"71", x"6b", x"56", x"2c", x"48", x"5c", x"5a", x"5e", x"62", 
        x"b0", x"a6", x"97", x"94", x"8f", x"7b", x"89", x"ab", x"a9", x"a5", x"a4", x"ad", x"ab", x"a4", x"98", 
        x"94", x"88", x"88", x"8e", x"80", x"6b", x"6b", x"54", x"62", x"79", x"44", x"3a", x"4c", x"94", x"72", 
        x"55", x"5b", x"a3", x"d7", x"ad", x"78", x"7e", x"6f", x"6f", x"81", x"93", x"75", x"6e", x"6b", x"6f", 
        x"73", x"7d", x"9b", x"a9", x"9f", x"cc", x"d4", x"a2", x"86", x"98", x"b9", x"a8", x"98", x"bc", x"cc", 
        x"cf", x"cd", x"ca", x"cc", x"d2", x"e8", x"eb", x"ef", x"eb", x"ec", x"ee", x"e8", x"eb", x"ec", x"eb", 
        x"ec", x"ec", x"ec", x"ec", x"ef", x"ef", x"ee", x"ee", x"eb", x"e4", x"db", x"c9", x"ba", x"ad", x"a3", 
        x"a0", x"a2", x"a3", x"a4", x"a5", x"a6", x"a8", x"aa", x"ab", x"ac", x"ac", x"ad", x"ad", x"ac", x"ac", 
        x"ab", x"ae", x"a9", x"7b", x"7a", x"a1", x"ab", x"ad", x"ac", x"ad", x"ab", x"ac", x"ac", x"ad", x"ac", 
        x"ac", x"ad", x"ac", x"ac", x"a8", x"ac", x"ae", x"68", x"60", x"7c", x"78", x"74", x"9c", x"ae", x"ac", 
        x"af", x"b3", x"b5", x"b7", x"a9", x"80", x"71", x"5b", x"45", x"2e", x"26", x"23", x"23", x"22", x"1e", 
        x"14", x"0e", x"63", x"dc", x"d6", x"d4", x"d7", x"d5", x"da", x"d6", x"cd", x"ce", x"ce", x"d4", x"d1", 
        x"d1", x"d1", x"d1", x"d1", x"d3", x"d4", x"d3", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d3", x"d4", 
        x"d3", x"d3", x"d4", x"d5", x"d6", x"d3", x"d3", x"d3", x"d0", x"d4", x"d4", x"d3", x"d4", x"d2", x"d1", 
        x"d3", x"d5", x"d5", x"d4", x"d3", x"d2", x"d3", x"d3", x"d5", x"d5", x"d8", x"d5", x"d1", x"d6", x"d5", 
        x"d6", x"d4", x"d2", x"e1", x"f5", x"ee", x"ed", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"ee", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ed", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"f1", x"f2", x"ef", x"ef", x"f1", x"ed", 
        x"ec", x"f2", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"f1", x"f2", x"f2", x"f2", x"f0", x"ee", x"ec", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"ef", x"f0", x"f1", x"f2", x"f2", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", 
        x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"f1", x"f3", x"f2", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", 
        x"f1", x"f2", x"f3", x"f2", x"f2", x"f3", x"f1", x"ef", x"ef", x"f1", x"f2", x"f1", x"ef", x"f1", x"f3", 
        x"f2", x"f1", x"f0", x"ef", x"f3", x"f2", x"f0", x"f4", x"f1", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", 
        x"ee", x"ef", x"f1", x"f5", x"f5", x"f1", x"f1", x"f1", x"ee", x"e7", x"dc", x"d6", x"c9", x"c1", x"bb", 
        x"b9", x"bf", x"c0", x"c6", x"ca", x"d2", x"d7", x"db", x"df", x"e2", x"e8", x"e9", x"ec", x"ef", x"f1", 
        x"f1", x"f1", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f1", x"f1", x"f1", x"f2", x"f3", 
        x"f1", x"f1", x"f3", x"f5", x"f4", x"f2", x"f3", x"f4", x"f6", x"f7", x"f7", x"f8", x"f8", x"f7", x"f6", 
        x"f4", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", x"f2", x"f0", x"f0", x"ef", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f3", 
        x"f3", x"f1", x"f1", x"f1", x"f0", x"f1", x"f4", x"f4", x"f3", x"ee", x"ef", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f3", x"f4", x"f4", x"f6", 
        x"f7", x"f6", x"f6", x"e5", x"84", x"4b", x"5c", x"bd", x"d9", x"d5", x"da", x"bc", x"a6", x"a3", x"9a", 
        x"9c", x"9b", x"9a", x"98", x"98", x"98", x"99", x"95", x"93", x"95", x"95", x"95", x"93", x"91", x"91", 
        x"91", x"91", x"8f", x"90", x"8f", x"8e", x"8c", x"90", x"7f", x"46", x"46", x"6d", x"8c", x"87", x"88", 
        x"86", x"85", x"84", x"85", x"81", x"74", x"71", x"73", x"74", x"73", x"73", x"73", x"75", x"74", x"81", 
        x"8e", x"8a", x"85", x"91", x"91", x"86", x"81", x"80", x"82", x"80", x"7d", x"51", x"4a", x"5e", x"89", 
        x"7c", x"7d", x"7e", x"7f", x"82", x"85", x"86", x"84", x"7f", x"78", x"74", x"6e", x"62", x"5c", x"5b", 
        x"5b", x"5e", x"65", x"6a", x"6f", x"71", x"76", x"7b", x"78", x"78", x"78", x"7e", x"7d", x"7a", x"71", 
        x"70", x"6e", x"4e", x"40", x"61", x"78", x"83", x"8b", x"9e", x"b2", x"c5", x"d3", x"dc", x"d8", x"a3", 
        x"80", x"84", x"81", x"80", x"7e", x"7e", x"7e", x"80", x"91", x"9a", x"82", x"6d", x"8e", x"8f", x"8b", 
        x"84", x"7c", x"68", x"55", x"58", x"5a", x"5c", x"66", x"5e", x"38", x"5f", x"84", x"86", x"80", x"7b", 
        x"b8", x"b7", x"af", x"af", x"9f", x"87", x"96", x"ac", x"9a", x"94", x"a9", x"aa", x"a8", x"a0", x"96", 
        x"8d", x"87", x"8e", x"81", x"80", x"58", x"60", x"55", x"60", x"7e", x"70", x"58", x"66", x"8b", x"77", 
        x"7a", x"83", x"9e", x"b4", x"a4", x"92", x"a4", x"92", x"89", x"7c", x"74", x"5f", x"6a", x"68", x"7c", 
        x"81", x"6a", x"84", x"ba", x"a9", x"ae", x"cf", x"ab", x"98", x"b2", x"ca", x"a8", x"a3", x"bf", x"c5", 
        x"d1", x"cc", x"d0", x"cb", x"cc", x"d2", x"d3", x"dc", x"dc", x"e2", x"e9", x"ea", x"ef", x"f1", x"ec", 
        x"eb", x"ee", x"ee", x"ea", x"ec", x"ed", x"ea", x"eb", x"eb", x"ee", x"f0", x"f0", x"ef", x"ec", x"e5", 
        x"da", x"cc", x"bf", x"b3", x"ac", x"a5", x"9e", x"9d", x"a1", x"a2", x"a5", x"ab", x"af", x"ae", x"ae", 
        x"ae", x"ae", x"a8", x"7c", x"7c", x"a0", x"a9", x"ac", x"ad", x"ac", x"aa", x"ac", x"ac", x"ac", x"ac", 
        x"ac", x"ad", x"ae", x"ae", x"a6", x"ad", x"ad", x"66", x"5c", x"7a", x"77", x"72", x"9e", x"bb", x"b6", 
        x"b5", x"a9", x"95", x"7a", x"64", x"3e", x"2e", x"25", x"25", x"22", x"1e", x"14", x"0d", x"07", x"04", 
        x"02", x"07", x"63", x"dd", x"d6", x"d4", x"d7", x"d3", x"d7", x"d9", x"cd", x"cf", x"cf", x"d3", x"d1", 
        x"d0", x"d2", x"d2", x"d1", x"d2", x"d3", x"d2", x"d2", x"d4", x"d4", x"d4", x"d3", x"d3", x"d5", x"d5", 
        x"d3", x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d2", x"d1", x"d4", x"d3", x"d2", x"d4", x"d2", x"d1", 
        x"d3", x"d5", x"d5", x"d3", x"d3", x"d2", x"d2", x"d3", x"d5", x"d4", x"d7", x"d5", x"d0", x"d6", x"d6", 
        x"d7", x"d5", x"d1", x"df", x"f3", x"ee", x"ee", x"ee", x"ee", x"f1", x"ef", x"ed", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ee", x"ed", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ed", 
        x"ec", x"f3", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"ef", x"ef", x"f0", x"f1", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"ea", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f2", 
        x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f3", x"f1", x"ee", x"ed", x"f0", x"f0", x"ef", x"f2", x"f2", x"f0", 
        x"f0", x"f1", x"ef", x"ec", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f1", x"f1", x"ef", 
        x"ee", x"f2", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f2", x"ef", 
        x"eb", x"e8", x"e2", x"dc", x"d4", x"cd", x"cb", x"c6", x"c6", x"c4", x"c9", x"c7", x"c6", x"ca", x"cd", 
        x"d4", x"d7", x"de", x"e4", x"ea", x"f0", x"f3", x"f4", x"f4", x"f4", x"f3", x"f1", x"f1", x"f1", x"f1", 
        x"ef", x"f1", x"f3", x"f5", x"f6", x"f5", x"f4", x"f4", x"f5", x"f5", x"f7", x"f6", x"f5", x"f5", x"f5", 
        x"f5", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f4", x"f3", x"f3", x"f0", x"f2", x"f1", 
        x"f2", x"f1", x"f0", x"f1", x"f2", x"f2", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f0", x"ef", x"f2", x"f5", x"f4", x"f2", x"ef", x"ef", x"f2", x"f1", x"f2", x"f1", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"ef", x"f0", x"f4", x"f7", x"f7", x"f6", 
        x"f9", x"f7", x"f6", x"e9", x"8c", x"4f", x"56", x"b7", x"db", x"d5", x"d6", x"d7", x"ac", x"97", x"9d", 
        x"9b", x"98", x"99", x"99", x"97", x"9a", x"9c", x"95", x"96", x"95", x"92", x"93", x"91", x"8f", x"8f", 
        x"91", x"91", x"8f", x"8d", x"8e", x"8e", x"8c", x"91", x"81", x"48", x"44", x"68", x"8c", x"88", x"88", 
        x"83", x"82", x"84", x"86", x"80", x"73", x"73", x"71", x"73", x"74", x"72", x"72", x"73", x"74", x"80", 
        x"8a", x"8a", x"87", x"8c", x"92", x"8e", x"84", x"81", x"83", x"81", x"7e", x"4e", x"4b", x"58", x"86", 
        x"7e", x"7e", x"7d", x"7c", x"7c", x"7d", x"7d", x"7b", x"7b", x"7e", x"80", x"81", x"82", x"84", x"83", 
        x"7f", x"79", x"75", x"69", x"62", x"5d", x"57", x"59", x"5b", x"52", x"45", x"52", x"5b", x"57", x"4d", 
        x"4f", x"53", x"48", x"48", x"7c", x"ad", x"c6", x"ca", x"d1", x"d4", x"d7", x"d9", x"dd", x"db", x"a3", 
        x"7b", x"7e", x"78", x"75", x"71", x"6d", x"68", x"68", x"76", x"82", x"6e", x"4c", x"6d", x"77", x"7c", 
        x"7f", x"90", x"8c", x"7b", x"7d", x"81", x"82", x"83", x"71", x"3b", x"56", x"7c", x"80", x"80", x"7a", 
        x"6f", x"81", x"81", x"88", x"8e", x"7e", x"84", x"a8", x"a3", x"a5", x"b3", x"ac", x"a7", x"a4", x"8f", 
        x"78", x"83", x"79", x"5f", x"77", x"6a", x"60", x"5f", x"6c", x"83", x"82", x"74", x"6f", x"80", x"ae", 
        x"c6", x"a2", x"a0", x"9c", x"85", x"89", x"a9", x"91", x"9c", x"96", x"85", x"76", x"73", x"58", x"69", 
        x"79", x"6a", x"76", x"8b", x"7e", x"79", x"9c", x"9d", x"96", x"9b", x"98", x"81", x"8b", x"a6", x"a9", 
        x"d1", x"e0", x"e6", x"d5", x"d1", x"d9", x"d9", x"d6", x"d1", x"d3", x"d6", x"d9", x"db", x"de", x"e2", 
        x"e4", x"eb", x"ec", x"eb", x"e7", x"ec", x"ec", x"ee", x"ec", x"ea", x"ed", x"ea", x"eb", x"ee", x"f0", 
        x"f0", x"ef", x"ed", x"e9", x"e3", x"d8", x"c8", x"bc", x"b3", x"a9", x"a6", x"a6", x"a5", x"a2", x"a3", 
        x"a7", x"ac", x"a9", x"80", x"7f", x"a2", x"ab", x"af", x"ad", x"ac", x"ae", x"ac", x"ab", x"ac", x"ad", 
        x"ac", x"aa", x"ad", x"ae", x"a9", x"af", x"ae", x"61", x"5e", x"7e", x"7c", x"79", x"95", x"a0", x"8a", 
        x"73", x"5e", x"49", x"37", x"31", x"26", x"22", x"1b", x"15", x"08", x"03", x"04", x"03", x"04", x"05", 
        x"09", x"14", x"60", x"dc", x"d7", x"d5", x"d7", x"d5", x"d8", x"da", x"cf", x"d0", x"d0", x"d2", x"d2", 
        x"d0", x"d1", x"d2", x"d1", x"d2", x"d3", x"d2", x"d1", x"d2", x"d4", x"d5", x"d4", x"d4", x"d4", x"d5", 
        x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"d4", x"d2", x"d2", x"d4", x"d3", x"d2", x"d4", x"d1", x"d1", 
        x"d1", x"d2", x"d3", x"d4", x"d3", x"d3", x"d0", x"d3", x"d6", x"d3", x"d4", x"d3", x"d0", x"d6", x"d5", 
        x"d6", x"d5", x"d2", x"df", x"f3", x"ed", x"ed", x"ee", x"ee", x"f1", x"f0", x"ef", x"ee", x"eb", x"ed", 
        x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"ee", x"ee", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ed", 
        x"ec", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", 
        x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f0", x"f0", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", 
        x"f1", x"f2", x"f1", x"ee", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f0", x"f1", x"f1", x"ef", 
        x"ee", x"f2", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", 
        x"f1", x"f2", x"f3", x"f4", x"f1", x"f2", x"f3", x"ee", x"ec", x"e5", x"e2", x"da", x"cf", x"c9", x"c3", 
        x"c2", x"c0", x"c5", x"c7", x"c8", x"cb", x"cf", x"d3", x"d7", x"df", x"e2", x"e6", x"ea", x"ef", x"f1", 
        x"f2", x"f2", x"f2", x"f4", x"f5", x"f6", x"f5", x"f3", x"f7", x"f7", x"f6", x"f5", x"f5", x"f5", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f3", x"f2", x"f3", x"f2", 
        x"f1", x"f0", x"ef", x"f0", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f3", 
        x"f2", x"f2", x"f1", x"f0", x"f1", x"f3", x"f5", x"f4", x"f2", x"ef", x"ef", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"ee", x"ef", x"f3", x"f7", x"f7", x"f6", 
        x"f7", x"f5", x"f5", x"eb", x"90", x"4f", x"52", x"b1", x"db", x"d6", x"d3", x"d9", x"c3", x"9e", x"99", 
        x"9b", x"9b", x"98", x"97", x"99", x"9b", x"9b", x"96", x"96", x"94", x"92", x"93", x"92", x"91", x"91", 
        x"92", x"91", x"90", x"8f", x"90", x"8f", x"8c", x"90", x"82", x"4b", x"45", x"66", x"8c", x"89", x"89", 
        x"84", x"83", x"84", x"85", x"80", x"73", x"71", x"70", x"72", x"73", x"72", x"6f", x"70", x"73", x"7f", 
        x"87", x"86", x"87", x"85", x"8d", x"94", x"8b", x"82", x"80", x"81", x"82", x"4e", x"4d", x"54", x"86", 
        x"7d", x"7e", x"7e", x"7d", x"7d", x"7f", x"80", x"7f", x"80", x"82", x"7f", x"7d", x"7c", x"79", x"78", 
        x"77", x"6f", x"70", x"66", x"57", x"5e", x"5b", x"59", x"5e", x"59", x"4e", x"57", x"5e", x"61", x"63", 
        x"6d", x"6b", x"5a", x"52", x"7f", x"ab", x"c3", x"c9", x"cd", x"cd", x"cd", x"cb", x"c8", x"c0", x"8c", 
        x"66", x"66", x"60", x"5d", x"5c", x"59", x"59", x"62", x"77", x"8e", x"85", x"55", x"8b", x"9d", x"9d", 
        x"9b", x"9f", x"98", x"82", x"7c", x"7c", x"80", x"82", x"75", x"42", x"51", x"79", x"7d", x"79", x"6c", 
        x"61", x"66", x"52", x"44", x"4b", x"4a", x"43", x"68", x"7e", x"9f", x"a9", x"b2", x"bc", x"b2", x"93", 
        x"86", x"92", x"74", x"56", x"64", x"78", x"69", x"68", x"79", x"8c", x"88", x"84", x"83", x"8c", x"b2", 
        x"d0", x"c1", x"9e", x"a5", x"86", x"7d", x"a0", x"80", x"9f", x"b0", x"97", x"61", x"5f", x"61", x"51", 
        x"79", x"77", x"90", x"7d", x"6f", x"6a", x"6e", x"5c", x"4d", x"5e", x"61", x"60", x"6a", x"82", x"7f", 
        x"a3", x"cb", x"e6", x"e8", x"e7", x"f4", x"ef", x"e6", x"e7", x"e4", x"e1", x"dc", x"da", x"d3", x"cf", 
        x"c8", x"c7", x"c3", x"c1", x"be", x"db", x"e8", x"ee", x"f0", x"ef", x"ef", x"e9", x"e9", x"ec", x"ed", 
        x"ec", x"ec", x"ec", x"ed", x"ef", x"f1", x"f2", x"f0", x"e9", x"df", x"d7", x"ce", x"c4", x"b5", x"aa", 
        x"a3", x"9e", x"9c", x"79", x"79", x"a4", x"ae", x"b2", x"b1", x"b1", x"af", x"ae", x"af", x"ad", x"ab", 
        x"ad", x"ad", x"ab", x"ac", x"a8", x"b1", x"b0", x"6b", x"5f", x"72", x"67", x"56", x"4f", x"4d", x"42", 
        x"37", x"31", x"2a", x"25", x"1d", x"11", x"06", x"02", x"03", x"04", x"03", x"03", x"0a", x"22", x"37", 
        x"4e", x"4c", x"69", x"da", x"d9", x"d7", x"d6", x"d7", x"d8", x"da", x"d0", x"d0", x"cf", x"d1", x"d3", 
        x"d0", x"d1", x"d2", x"d1", x"d2", x"d4", x"d2", x"d1", x"d2", x"d4", x"d5", x"d4", x"d4", x"d4", x"d4", 
        x"d2", x"d4", x"d5", x"d5", x"d5", x"d4", x"d3", x"d2", x"d2", x"d5", x"d4", x"d3", x"d4", x"d1", x"d1", 
        x"d1", x"d1", x"d2", x"d4", x"d5", x"d4", x"d0", x"d2", x"d6", x"d4", x"d4", x"d3", x"d0", x"d6", x"d4", 
        x"d6", x"d5", x"d2", x"df", x"f3", x"ef", x"ef", x"ee", x"ee", x"f0", x"ef", x"ee", x"ed", x"eb", x"ed", 
        x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f1", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", 
        x"f1", x"ef", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"ed", 
        x"ec", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f1", 
        x"f0", x"f0", x"f0", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f3", x"f4", x"f2", x"f0", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", 
        x"ee", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f2", x"f0", x"f1", x"f2", x"f2", x"f3", x"f2", x"f5", x"f4", x"f2", x"f2", x"ef", 
        x"ec", x"e8", x"e5", x"e0", x"d8", x"d0", x"cb", x"c6", x"c5", x"c7", x"c6", x"c3", x"c3", x"c8", x"cc", 
        x"cf", x"d7", x"dd", x"e4", x"ec", x"f2", x"f4", x"f5", x"f8", x"f9", x"f7", x"f6", x"f6", x"f5", x"f0", 
        x"ef", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f3", x"f2", x"f1", x"f3", x"f3", x"f2", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"ef", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f5", x"f6", x"f4", x"f2", x"ef", x"ef", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"f2", x"f6", x"f8", x"f6", 
        x"f6", x"f4", x"f5", x"ed", x"95", x"4f", x"4f", x"ad", x"db", x"d7", x"d2", x"d9", x"d5", x"a8", x"98", 
        x"9c", x"9b", x"98", x"97", x"9a", x"99", x"99", x"97", x"96", x"94", x"95", x"94", x"93", x"92", x"93", 
        x"92", x"91", x"90", x"8f", x"90", x"91", x"8c", x"8e", x"83", x"4d", x"46", x"65", x"8a", x"89", x"8a", 
        x"86", x"85", x"84", x"83", x"80", x"72", x"6f", x"6f", x"71", x"73", x"75", x"6f", x"6e", x"70", x"7a", 
        x"81", x"84", x"86", x"83", x"89", x"92", x"8e", x"85", x"7d", x"7e", x"82", x"51", x"50", x"55", x"8a", 
        x"7c", x"7f", x"85", x"86", x"86", x"85", x"80", x"79", x"73", x"68", x"60", x"5e", x"5c", x"58", x"5c", 
        x"65", x"65", x"6d", x"63", x"4a", x"68", x"79", x"79", x"7b", x"7d", x"79", x"79", x"74", x"6f", x"73", 
        x"76", x"71", x"5e", x"4a", x"6f", x"95", x"a8", x"a4", x"9e", x"99", x"97", x"9b", x"a2", x"a6", x"81", 
        x"5e", x"65", x"6c", x"71", x"74", x"74", x"75", x"7a", x"93", x"a3", x"93", x"57", x"91", x"9c", x"9b", 
        x"9d", x"9e", x"99", x"82", x"76", x"74", x"73", x"72", x"63", x"3b", x"41", x"5f", x"65", x"64", x"56", 
        x"c8", x"d1", x"bf", x"95", x"72", x"5e", x"37", x"5e", x"70", x"74", x"56", x"4b", x"53", x"5f", x"78", 
        x"92", x"98", x"7e", x"70", x"74", x"7d", x"70", x"7b", x"88", x"81", x"65", x"79", x"8f", x"8e", x"90", 
        x"a7", x"9d", x"99", x"b2", x"89", x"8e", x"8d", x"77", x"a9", x"bc", x"9b", x"6b", x"a5", x"84", x"71", 
        x"60", x"70", x"8a", x"6d", x"66", x"7f", x"8d", x"7d", x"6d", x"67", x"60", x"5b", x"70", x"7f", x"57", 
        x"4c", x"73", x"86", x"88", x"9f", x"c2", x"ce", x"bf", x"dd", x"ed", x"f2", x"f1", x"f1", x"f0", x"e4", 
        x"d9", x"d5", x"c8", x"af", x"b1", x"cd", x"d1", x"cf", x"d6", x"de", x"e3", x"ea", x"ed", x"ef", x"ef", 
        x"ed", x"ec", x"ec", x"ee", x"ec", x"eb", x"eb", x"ec", x"ec", x"ec", x"eb", x"e9", x"ea", x"e5", x"e1", 
        x"da", x"d0", x"c6", x"8b", x"74", x"a1", x"a8", x"a5", x"a0", x"a4", x"ad", x"ad", x"b0", x"af", x"ad", 
        x"b0", x"ae", x"b0", x"b4", x"af", x"a6", x"90", x"59", x"3d", x"44", x"43", x"3e", x"36", x"31", x"28", 
        x"1c", x"15", x"0c", x"08", x"05", x"07", x"08", x"0a", x"0f", x"1e", x"35", x"4a", x"5f", x"78", x"7b", 
        x"7e", x"65", x"6b", x"d8", x"d9", x"d7", x"d7", x"d6", x"d7", x"d9", x"ce", x"d0", x"ce", x"d0", x"d3", 
        x"d1", x"d2", x"d1", x"d0", x"d2", x"d4", x"d3", x"d2", x"d3", x"d4", x"d3", x"d2", x"d3", x"d4", x"d4", 
        x"d2", x"d3", x"d5", x"d5", x"d5", x"d4", x"d3", x"d3", x"d3", x"d6", x"d4", x"d3", x"d3", x"d0", x"d1", 
        x"d0", x"d0", x"d2", x"d4", x"d5", x"d5", x"d2", x"d3", x"d6", x"d5", x"d7", x"d5", x"d0", x"d5", x"d4", 
        x"d6", x"d6", x"d3", x"e0", x"f4", x"f0", x"ef", x"ee", x"ef", x"ee", x"ef", x"ee", x"ee", x"ed", x"ee", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ef", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"ee", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"ed", 
        x"eb", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f1", x"f1", x"f2", 
        x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", 
        x"ef", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f1", x"f2", x"f3", x"f2", x"f3", x"f2", x"f4", x"f2", x"f2", x"f2", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f0", x"ed", x"ec", x"e9", x"e5", x"e1", x"dd", x"d8", x"d4", 
        x"d0", x"cd", x"cb", x"ca", x"ca", x"ca", x"cc", x"ce", x"d7", x"df", x"e3", x"e8", x"ec", x"ef", x"f2", 
        x"f2", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f1", x"f1", x"f1", x"f3", x"f2", x"f2", 
        x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f2", x"f1", x"f0", x"f1", x"f2", x"f2", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f2", x"f4", x"f6", x"f7", x"f4", x"f2", x"ef", x"ef", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f2", x"f0", x"f0", x"f2", x"f5", x"f7", x"f6", 
        x"f6", x"f6", x"f6", x"f0", x"9a", x"4e", x"4d", x"a7", x"db", x"d8", x"d3", x"d8", x"d6", x"ad", x"98", 
        x"9b", x"9b", x"99", x"99", x"99", x"96", x"96", x"96", x"95", x"93", x"95", x"93", x"92", x"92", x"91", 
        x"90", x"90", x"90", x"8e", x"8e", x"91", x"8d", x"8e", x"84", x"4e", x"45", x"62", x"89", x"8a", x"8a", 
        x"89", x"86", x"85", x"86", x"83", x"74", x"6f", x"6f", x"70", x"72", x"74", x"70", x"70", x"70", x"77", 
        x"81", x"88", x"86", x"87", x"8c", x"92", x"91", x"8a", x"82", x"82", x"83", x"59", x"4e", x"51", x"81", 
        x"7b", x"73", x"6d", x"66", x"60", x"5d", x"5d", x"5e", x"63", x"6c", x"6d", x"72", x"75", x"75", x"79", 
        x"7d", x"7f", x"85", x"7b", x"5e", x"74", x"83", x"7c", x"7e", x"7b", x"77", x"7c", x"7c", x"71", x"69", 
        x"69", x"60", x"50", x"36", x"5b", x"82", x"99", x"a5", x"b0", x"b8", x"c1", x"c5", x"cb", x"ce", x"9b", 
        x"58", x"5d", x"63", x"64", x"66", x"69", x"6c", x"6f", x"8a", x"a1", x"96", x"5f", x"8a", x"8f", x"89", 
        x"84", x"7c", x"79", x"67", x"5c", x"5a", x"5c", x"5e", x"54", x"35", x"35", x"52", x"5a", x"5b", x"57", 
        x"d1", x"e5", x"e3", x"e0", x"d4", x"c2", x"6a", x"9c", x"b8", x"aa", x"99", x"78", x"57", x"5f", x"75", 
        x"83", x"89", x"85", x"8a", x"94", x"91", x"83", x"85", x"8b", x"7b", x"72", x"85", x"89", x"79", x"75", 
        x"89", x"88", x"8f", x"98", x"83", x"81", x"90", x"86", x"97", x"98", x"78", x"5e", x"b7", x"a2", x"94", 
        x"63", x"6c", x"81", x"6f", x"5f", x"73", x"7d", x"86", x"9e", x"8c", x"6a", x"5f", x"78", x"7c", x"5b", 
        x"6b", x"7a", x"6d", x"4b", x"57", x"91", x"c5", x"93", x"8b", x"9e", x"b9", x"c8", x"d9", x"e8", x"ed", 
        x"ed", x"ee", x"e9", x"d3", x"dc", x"eb", x"e5", x"dd", x"d7", x"d0", x"cb", x"ca", x"ce", x"d4", x"da", 
        x"e1", x"e6", x"e9", x"ee", x"ef", x"ec", x"ec", x"ec", x"eb", x"eb", x"ec", x"eb", x"ed", x"ec", x"ed", 
        x"ee", x"ed", x"e4", x"9b", x"7a", x"b7", x"c7", x"bd", x"ad", x"a8", x"a9", x"a1", x"a4", x"ab", x"b4", 
        x"ba", x"b4", x"a0", x"88", x"69", x"50", x"4a", x"43", x"37", x"34", x"2c", x"20", x"15", x"11", x"0c", 
        x"03", x"02", x"04", x"0a", x"0e", x"15", x"2c", x"43", x"59", x"6b", x"78", x"80", x"7b", x"7e", x"7b", 
        x"7a", x"69", x"66", x"d6", x"db", x"d6", x"d7", x"d5", x"d7", x"d7", x"cc", x"d0", x"ce", x"d0", x"d3", 
        x"d2", x"d3", x"d2", x"d0", x"d1", x"d3", x"d2", x"d2", x"d3", x"d4", x"d3", x"d2", x"d2", x"d4", x"d5", 
        x"d4", x"d4", x"d3", x"d3", x"d5", x"d6", x"d6", x"d4", x"d4", x"d6", x"d4", x"d3", x"d3", x"d1", x"d1", 
        x"d1", x"d2", x"d3", x"d4", x"d5", x"d4", x"d4", x"d4", x"d6", x"d5", x"d9", x"d7", x"d1", x"d4", x"d3", 
        x"d6", x"d6", x"d3", x"e0", x"f4", x"ef", x"ed", x"ed", x"ee", x"ee", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", 
        x"ef", x"ee", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ed", 
        x"eb", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", 
        x"f0", x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f3", x"f4", x"f1", x"f0", x"f2", 
        x"f4", x"f4", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f0", 
        x"ef", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"ef", x"ef", x"f1", x"f2", x"f3", 
        x"f1", x"f1", x"f4", x"f3", x"f0", x"f0", x"f1", x"f4", x"f6", x"f3", x"f1", x"f2", x"f3", x"f3", x"f1", 
        x"f0", x"ec", x"ea", x"e9", x"e5", x"dd", x"d7", x"d2", x"d0", x"cf", x"cd", x"c9", x"c5", x"c6", x"ca", 
        x"d0", x"d6", x"dc", x"e3", x"e9", x"ee", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f2", x"f1", x"f0", x"ef", x"f1", x"f4", x"f4", x"f2", x"f1", 
        x"f1", x"f0", x"f1", x"f3", x"f5", x"f6", x"f7", x"f4", x"f2", x"ef", x"ef", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f4", x"f6", x"f6", 
        x"f6", x"f7", x"f7", x"f2", x"a0", x"4f", x"4a", x"a3", x"db", x"d8", x"d5", x"d9", x"d9", x"b3", x"99", 
        x"9b", x"9a", x"97", x"95", x"98", x"96", x"95", x"97", x"95", x"93", x"93", x"93", x"92", x"91", x"91", 
        x"91", x"90", x"8f", x"8d", x"8d", x"91", x"8d", x"8e", x"86", x"50", x"44", x"5e", x"86", x"8a", x"8a", 
        x"8a", x"87", x"86", x"89", x"87", x"77", x"6e", x"6f", x"6f", x"71", x"74", x"73", x"73", x"71", x"77", 
        x"7f", x"84", x"82", x"86", x"90", x"9a", x"96", x"88", x"7f", x"76", x"6f", x"4e", x"3d", x"38", x"5d", 
        x"62", x"65", x"6a", x"6c", x"6f", x"74", x"79", x"7a", x"7d", x"81", x"7f", x"80", x"81", x"7d", x"7e", 
        x"82", x"84", x"81", x"7c", x"64", x"71", x"7a", x"70", x"6d", x"63", x"58", x"58", x"5b", x"57", x"58", 
        x"67", x"6a", x"62", x"44", x"6f", x"a2", x"bd", x"c7", x"cd", x"d4", x"db", x"d9", x"da", x"db", x"b1", 
        x"6c", x"68", x"65", x"5c", x"58", x"58", x"5c", x"5d", x"6d", x"78", x"6b", x"41", x"65", x"70", x"6d", 
        x"6f", x"6f", x"6a", x"58", x"51", x"56", x"56", x"5c", x"62", x"45", x"40", x"71", x"7f", x"80", x"84", 
        x"d1", x"db", x"e3", x"e0", x"e1", x"de", x"7d", x"9c", x"d7", x"dd", x"e9", x"cf", x"ae", x"ce", x"ce", 
        x"bf", x"b2", x"a9", x"91", x"80", x"78", x"72", x"60", x"67", x"72", x"93", x"95", x"93", x"82", x"8c", 
        x"ad", x"a9", x"81", x"7f", x"9c", x"91", x"7b", x"75", x"80", x"8a", x"8a", x"6b", x"a5", x"b6", x"aa", 
        x"72", x"5d", x"72", x"79", x"6d", x"6f", x"7e", x"95", x"ad", x"8b", x"6d", x"70", x"8f", x"9d", x"7c", 
        x"90", x"94", x"7b", x"63", x"80", x"ae", x"e3", x"ac", x"87", x"8a", x"88", x"7f", x"87", x"86", x"97", 
        x"a9", x"bc", x"d3", x"db", x"e7", x"f2", x"f4", x"f4", x"f0", x"ed", x"ea", x"e4", x"df", x"da", x"d3", 
        x"cc", x"c8", x"c4", x"cc", x"d4", x"da", x"e6", x"ec", x"ec", x"ed", x"ee", x"ed", x"ef", x"ee", x"ee", 
        x"ed", x"ed", x"e8", x"9b", x"73", x"be", x"d8", x"da", x"d5", x"d4", x"db", x"d0", x"c8", x"b7", x"98", 
        x"79", x"58", x"47", x"45", x"45", x"3e", x"33", x"28", x"16", x"0f", x"0b", x"07", x"05", x"05", x"07", 
        x"0c", x"15", x"27", x"4a", x"67", x"6e", x"7e", x"80", x"7f", x"7a", x"7e", x"7a", x"7f", x"8b", x"8d", 
        x"93", x"80", x"6d", x"d6", x"dc", x"d5", x"d8", x"db", x"d8", x"d6", x"cc", x"d1", x"d0", x"d1", x"d4", 
        x"d2", x"d2", x"d3", x"d3", x"d2", x"d2", x"d0", x"d1", x"d2", x"d3", x"d3", x"d2", x"d2", x"d4", x"d5", 
        x"d4", x"d4", x"d4", x"d4", x"d4", x"d6", x"d6", x"d5", x"d4", x"d6", x"d4", x"d3", x"d4", x"d2", x"d2", 
        x"d3", x"d4", x"d5", x"d5", x"d4", x"d3", x"d3", x"d4", x"d6", x"d5", x"d8", x"d6", x"d1", x"d4", x"d2", 
        x"d6", x"d6", x"d4", x"e0", x"f4", x"ef", x"ed", x"ec", x"ee", x"ed", x"f0", x"f2", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"ec", 
        x"eb", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f2", x"f0", x"ef", x"f0", x"f1", x"f1", x"ef", x"ee", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f1", x"f3", x"f4", x"f2", x"f0", x"f1", 
        x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", 
        x"ef", x"f3", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f3", x"f4", x"f2", x"f1", x"f0", x"f3", 
        x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"ef", x"ef", x"f2", x"f2", x"f1", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f4", x"f8", x"f8", x"f3", x"f0", x"ee", x"ef", x"ef", x"ed", x"ea", x"e3", x"da", x"d1", 
        x"cc", x"c8", x"c5", x"c2", x"c1", x"c3", x"c6", x"cc", x"d6", x"db", x"e2", x"e6", x"ec", x"ed", x"f0", 
        x"f0", x"f1", x"f2", x"f2", x"f0", x"f0", x"f1", x"f3", x"f2", x"f1", x"f3", x"f5", x"f5", x"f1", x"f1", 
        x"f2", x"f0", x"f1", x"f3", x"f5", x"f5", x"f6", x"f4", x"f2", x"ef", x"ef", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f4", x"f6", x"f6", 
        x"f5", x"f7", x"f7", x"f5", x"a7", x"52", x"46", x"9c", x"da", x"d7", x"d4", x"d7", x"d7", x"b4", x"98", 
        x"9c", x"9b", x"99", x"97", x"98", x"98", x"96", x"99", x"96", x"95", x"93", x"94", x"93", x"91", x"91", 
        x"92", x"91", x"90", x"8e", x"8d", x"90", x"8e", x"8f", x"8a", x"55", x"45", x"5c", x"85", x"89", x"89", 
        x"8b", x"87", x"85", x"86", x"86", x"77", x"6e", x"72", x"72", x"73", x"71", x"6f", x"71", x"73", x"7e", 
        x"86", x"86", x"7d", x"73", x"6b", x"6a", x"62", x"57", x"5a", x"60", x"64", x"4b", x"45", x"44", x"75", 
        x"7e", x"7f", x"81", x"81", x"81", x"81", x"81", x"7e", x"7e", x"7f", x"81", x"84", x"85", x"80", x"7c", 
        x"77", x"6e", x"66", x"5d", x"3d", x"4d", x"61", x"60", x"68", x"6a", x"6e", x"75", x"79", x"74", x"72", 
        x"76", x"7c", x"74", x"45", x"6f", x"aa", x"c2", x"ca", x"cd", x"d2", x"d8", x"d5", x"d2", x"ce", x"ae", 
        x"6f", x"66", x"61", x"57", x"51", x"49", x"4b", x"4e", x"59", x"62", x"5b", x"34", x"55", x"69", x"62", 
        x"6d", x"82", x"89", x"80", x"7b", x"80", x"86", x"8b", x"89", x"59", x"45", x"7d", x"8b", x"8d", x"89", 
        x"b7", x"a7", x"b5", x"c9", x"d3", x"e5", x"9a", x"b3", x"e5", x"ec", x"e1", x"ca", x"d4", x"ee", x"e8", 
        x"e4", x"da", x"e2", x"cd", x"cb", x"b0", x"a4", x"99", x"81", x"79", x"7a", x"63", x"76", x"73", x"93", 
        x"b1", x"97", x"6d", x"7e", x"83", x"83", x"79", x"70", x"5b", x"65", x"77", x"8d", x"a5", x"86", x"84", 
        x"7c", x"62", x"5f", x"7d", x"6c", x"6d", x"81", x"71", x"6b", x"68", x"82", x"7c", x"77", x"7a", x"7c", 
        x"92", x"9b", x"9d", x"ad", x"ac", x"a4", x"d4", x"a9", x"8c", x"9b", x"99", x"94", x"90", x"8a", x"90", 
        x"8a", x"7f", x"7c", x"80", x"8b", x"a3", x"b9", x"ca", x"d6", x"e2", x"e9", x"f0", x"f1", x"f1", x"ef", 
        x"ee", x"eb", x"e6", x"de", x"d4", x"c9", x"c3", x"c4", x"c8", x"d1", x"db", x"e0", x"e3", x"e7", x"e9", 
        x"ec", x"f1", x"ea", x"9d", x"73", x"c3", x"da", x"db", x"d9", x"d1", x"bb", x"9a", x"78", x"52", x"3b", 
        x"3e", x"3f", x"36", x"28", x"18", x"0b", x"0e", x"15", x"1d", x"15", x"08", x"04", x"08", x"1f", x"42", 
        x"6c", x"8c", x"a7", x"b9", x"ae", x"83", x"78", x"76", x"77", x"70", x"70", x"6a", x"97", x"b2", x"9c", 
        x"8f", x"77", x"6a", x"d3", x"db", x"d5", x"d7", x"d5", x"d8", x"d7", x"cc", x"d1", x"d2", x"d2", x"d4", 
        x"d2", x"d3", x"d4", x"d5", x"d4", x"d2", x"cf", x"d0", x"d2", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", 
        x"d2", x"d4", x"d6", x"d6", x"d5", x"d4", x"d4", x"d6", x"d5", x"d6", x"d4", x"d3", x"d4", x"d3", x"d2", 
        x"d4", x"d6", x"d6", x"d4", x"d3", x"d3", x"d1", x"d4", x"d7", x"d4", x"d6", x"d4", x"d1", x"d4", x"d3", 
        x"d5", x"d6", x"d4", x"e0", x"f3", x"f1", x"ee", x"ed", x"ee", x"ec", x"ee", x"f0", x"ed", x"ed", x"ef", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", 
        x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"ec", 
        x"ea", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f2", x"f0", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"f1", x"f2", x"f1", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f1", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f4", x"f4", x"f2", x"f2", x"f3", x"f2", x"f0", x"f1", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", 
        x"ef", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", 
        x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f4", x"f2", x"f0", x"f0", x"f1", x"f2", 
        x"f3", x"f1", x"f3", x"f6", x"f5", x"f2", x"f1", x"f5", x"f8", x"f6", x"f3", x"f3", x"f4", x"f3", x"f0", 
        x"ee", x"ef", x"ef", x"ee", x"eb", x"e3", x"db", x"d4", x"c9", x"c7", x"c5", x"c0", x"c1", x"c2", x"c6", 
        x"ce", x"d3", x"da", x"e0", x"e5", x"e9", x"ec", x"ef", x"f1", x"f2", x"f5", x"f6", x"f4", x"f0", x"f2", 
        x"f3", x"f1", x"f2", x"f3", x"f5", x"f5", x"f6", x"f4", x"f2", x"ef", x"ef", x"f2", x"f1", x"f3", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f2", x"f1", x"f0", x"f0", x"f4", x"f7", x"f6", 
        x"f4", x"f6", x"f7", x"f6", x"ae", x"56", x"43", x"95", x"d9", x"d7", x"d2", x"d5", x"d9", x"b8", x"9b", 
        x"9f", x"9a", x"99", x"9b", x"98", x"98", x"97", x"9a", x"98", x"97", x"95", x"94", x"94", x"92", x"92", 
        x"93", x"92", x"91", x"90", x"8e", x"8f", x"8d", x"90", x"8d", x"59", x"46", x"59", x"83", x"89", x"8a", 
        x"8e", x"8b", x"89", x"89", x"89", x"7a", x"71", x"74", x"73", x"73", x"6e", x"67", x"5f", x"59", x"54", 
        x"56", x"59", x"60", x"65", x"6d", x"80", x"8a", x"85", x"87", x"88", x"8a", x"61", x"51", x"4c", x"83", 
        x"80", x"7c", x"7e", x"7f", x"80", x"81", x"7e", x"79", x"75", x"6c", x"62", x"5e", x"5c", x"5a", x"5b", 
        x"62", x"67", x"72", x"72", x"4d", x"64", x"81", x"80", x"7d", x"7c", x"7b", x"79", x"76", x"71", x"76", 
        x"75", x"79", x"75", x"47", x"6b", x"a4", x"b8", x"b9", x"ae", x"a6", x"a1", x"9b", x"96", x"92", x"84", 
        x"56", x"4a", x"4a", x"41", x"4b", x"4d", x"51", x"57", x"69", x"87", x"91", x"60", x"78", x"99", x"92", 
        x"83", x"7d", x"78", x"77", x"7e", x"89", x"8c", x"86", x"7e", x"50", x"33", x"54", x"5a", x"53", x"47", 
        x"e1", x"d5", x"bc", x"bb", x"cb", x"da", x"aa", x"c1", x"e5", x"e8", x"c3", x"cd", x"ea", x"ea", x"e9", 
        x"e5", x"e8", x"dd", x"b2", x"c9", x"b8", x"95", x"c5", x"aa", x"7f", x"94", x"a7", x"9b", x"8c", x"a3", 
        x"a2", x"85", x"9a", x"99", x"77", x"7b", x"61", x"6b", x"4f", x"5e", x"78", x"8d", x"96", x"a3", x"99", 
        x"85", x"71", x"77", x"8a", x"7c", x"72", x"71", x"63", x"6b", x"84", x"77", x"74", x"66", x"7d", x"8f", 
        x"83", x"8e", x"95", x"9b", x"9a", x"ab", x"d9", x"a8", x"88", x"94", x"91", x"8d", x"99", x"9f", x"9d", 
        x"9d", x"9c", x"9a", x"96", x"8f", x"8b", x"88", x"8b", x"92", x"95", x"9f", x"be", x"d3", x"dc", x"e2", 
        x"eb", x"ec", x"ed", x"f0", x"f4", x"ee", x"e8", x"e5", x"dc", x"d3", x"cc", x"c4", x"c2", x"c7", x"cd", 
        x"d4", x"e3", x"e0", x"9f", x"79", x"be", x"c2", x"a7", x"87", x"67", x"4a", x"3f", x"3d", x"3a", x"2f", 
        x"25", x"14", x"0d", x"15", x"1f", x"30", x"4b", x"74", x"8f", x"4f", x"17", x"07", x"20", x"7f", x"ab", 
        x"b0", x"b1", x"ae", x"b0", x"9b", x"85", x"96", x"a7", x"9a", x"6b", x"71", x"72", x"92", x"a0", x"98", 
        x"93", x"79", x"6b", x"ce", x"d9", x"d3", x"d5", x"d6", x"d8", x"d9", x"cb", x"d0", x"d0", x"d0", x"d1", 
        x"d3", x"d3", x"d2", x"d3", x"d4", x"d4", x"d3", x"d4", x"d5", x"d3", x"d2", x"d3", x"d4", x"d4", x"d4", 
        x"d4", x"d4", x"d5", x"d4", x"d5", x"d5", x"d6", x"d5", x"d4", x"d5", x"d4", x"d4", x"d4", x"d3", x"d3", 
        x"d3", x"d4", x"d4", x"d4", x"d3", x"d2", x"d1", x"d3", x"d4", x"d4", x"d8", x"d6", x"d0", x"d4", x"d3", 
        x"d4", x"d4", x"d4", x"df", x"f3", x"f0", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ed", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ed", x"ed", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f1", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"ef", x"ee", 
        x"e8", x"f1", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"ed", x"f1", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f5", x"f8", x"f6", x"f2", x"f1", x"f2", x"f6", x"f7", x"f5", x"f3", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f0", x"ee", x"f0", x"ef", x"eb", x"e6", x"df", x"d7", 
        x"d0", x"cb", x"c6", x"c3", x"c5", x"c7", x"c8", x"cc", x"d1", x"d9", x"df", x"e2", x"e5", x"e9", x"ec", 
        x"ed", x"ef", x"f4", x"f6", x"f5", x"f6", x"f6", x"f5", x"f3", x"f0", x"ee", x"f1", x"ef", x"f4", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f1", x"f2", x"f1", x"f2", 
        x"ed", x"f2", x"f1", x"f0", x"ef", x"ed", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f5", x"f6", x"f6", 
        x"f7", x"f7", x"f6", x"f6", x"b8", x"5d", x"43", x"8c", x"d9", x"d6", x"d3", x"d6", x"d9", x"bc", x"9c", 
        x"a1", x"9b", x"9b", x"99", x"9b", x"9b", x"99", x"97", x"95", x"94", x"94", x"92", x"95", x"95", x"92", 
        x"93", x"90", x"91", x"92", x"8c", x"8f", x"8f", x"91", x"8f", x"5f", x"47", x"59", x"81", x"8a", x"8c", 
        x"8c", x"8d", x"87", x"7e", x"78", x"6a", x"5f", x"5c", x"58", x"53", x"56", x"5c", x"61", x"69", x"4e", 
        x"59", x"82", x"87", x"88", x"89", x"8e", x"95", x"8b", x"83", x"82", x"86", x"5f", x"4d", x"4b", x"76", 
        x"7a", x"71", x"6e", x"66", x"62", x"63", x"60", x"5f", x"63", x"67", x"69", x"70", x"77", x"7a", x"7d", 
        x"82", x"7f", x"80", x"81", x"5a", x"64", x"7d", x"7e", x"7b", x"77", x"75", x"77", x"78", x"71", x"74", 
        x"73", x"70", x"65", x"3d", x"4d", x"73", x"84", x"8e", x"93", x"a2", x"af", x"bd", x"c3", x"c8", x"ab", 
        x"66", x"61", x"6c", x"48", x"68", x"81", x"83", x"86", x"8c", x"92", x"91", x"67", x"6e", x"89", x"83", 
        x"78", x"6c", x"5e", x"50", x"3e", x"3e", x"41", x"2e", x"37", x"34", x"27", x"40", x"51", x"5b", x"51", 
        x"ed", x"ed", x"e5", x"d5", x"b1", x"b7", x"9a", x"b5", x"d7", x"cd", x"a4", x"d9", x"ec", x"e8", x"ea", 
        x"e5", x"e8", x"b7", x"7d", x"7e", x"a9", x"9e", x"ba", x"a1", x"89", x"bf", x"d8", x"c6", x"a4", x"ab", 
        x"aa", x"97", x"bf", x"bf", x"94", x"99", x"87", x"84", x"7a", x"6e", x"66", x"69", x"61", x"7f", x"91", 
        x"80", x"5e", x"6b", x"81", x"86", x"86", x"66", x"6d", x"81", x"77", x"66", x"50", x"51", x"94", x"9c", 
        x"9f", x"9d", x"69", x"86", x"8f", x"a9", x"db", x"a4", x"86", x"89", x"86", x"96", x"9f", x"9e", x"9e", 
        x"a0", x"9c", x"9b", x"a0", x"a0", x"9a", x"99", x"9a", x"9b", x"95", x"8b", x"71", x"80", x"99", x"aa", 
        x"b7", x"bf", x"ca", x"da", x"e4", x"e7", x"eb", x"ef", x"ee", x"f0", x"f2", x"eb", x"e4", x"dc", x"d4", 
        x"ca", x"cb", x"cb", x"8e", x"5b", x"6e", x"5b", x"42", x"38", x"3b", x"35", x"2d", x"1e", x"10", x"08", 
        x"0b", x"22", x"3e", x"60", x"89", x"b6", x"d2", x"e4", x"cf", x"63", x"30", x"14", x"30", x"b8", x"d2", 
        x"ba", x"b1", x"a8", x"a8", x"a8", x"a8", x"b0", x"b3", x"9e", x"6e", x"6e", x"6a", x"86", x"98", x"93", 
        x"91", x"7a", x"6d", x"ce", x"d9", x"d7", x"d9", x"d5", x"d8", x"da", x"cc", x"d0", x"d1", x"d1", x"d3", 
        x"d3", x"d2", x"d2", x"d2", x"d3", x"d4", x"d3", x"d4", x"d3", x"d3", x"d4", x"d4", x"d4", x"d2", x"d3", 
        x"d4", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d4", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d2", 
        x"d2", x"d3", x"d4", x"d6", x"d5", x"d4", x"d2", x"d4", x"d3", x"d4", x"d8", x"d6", x"d0", x"d2", x"d1", 
        x"d3", x"d5", x"d5", x"df", x"f2", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"f0", x"ef", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"ed", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", 
        x"e8", x"f1", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f0", x"f1", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f2", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"ed", x"f1", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f3", x"f6", x"f9", x"f7", x"f3", x"f1", x"f2", x"f4", x"f5", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f2", x"ef", x"f1", x"f1", x"f1", x"f3", x"f2", x"ef", 
        x"f2", x"f1", x"f0", x"ef", x"eb", x"e5", x"de", x"d5", x"cd", x"c5", x"c1", x"c3", x"c6", x"c8", x"cb", 
        x"ce", x"d5", x"de", x"e3", x"e6", x"e8", x"eb", x"ee", x"ef", x"ef", x"f0", x"f2", x"ee", x"f3", x"f2", 
        x"f1", x"f2", x"f0", x"f0", x"ef", x"f0", x"ef", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"ed", x"ee", 
        x"eb", x"f1", x"f1", x"f1", x"f1", x"ee", x"f0", x"f0", x"ef", x"f0", x"f0", x"f2", x"f6", x"f5", x"f5", 
        x"f6", x"f6", x"f7", x"f8", x"be", x"5f", x"42", x"89", x"d6", x"d6", x"d4", x"d5", x"da", x"bd", x"99", 
        x"9e", x"9c", x"9d", x"9b", x"99", x"9a", x"99", x"96", x"92", x"92", x"94", x"95", x"8f", x"92", x"90", 
        x"91", x"93", x"92", x"93", x"94", x"94", x"92", x"94", x"90", x"63", x"48", x"52", x"75", x"79", x"77", 
        x"73", x"6c", x"66", x"64", x"65", x"60", x"5d", x"67", x"6f", x"73", x"75", x"78", x"79", x"7a", x"60", 
        x"65", x"82", x"84", x"85", x"85", x"82", x"8a", x"87", x"7b", x"74", x"74", x"55", x"42", x"36", x"5a", 
        x"63", x"5f", x"66", x"6b", x"70", x"76", x"79", x"7b", x"7f", x"81", x"7f", x"7e", x"7e", x"7c", x"7c", 
        x"82", x"82", x"7d", x"7e", x"60", x"68", x"7d", x"75", x"72", x"6e", x"67", x"63", x"60", x"58", x"57", 
        x"5b", x"58", x"51", x"39", x"50", x"74", x"9c", x"b4", x"bc", x"c7", x"cb", x"d4", x"d8", x"db", x"c9", 
        x"94", x"93", x"9c", x"6f", x"7e", x"8d", x"84", x"7e", x"72", x"68", x"63", x"45", x"44", x"4b", x"41", 
        x"39", x"35", x"36", x"36", x"38", x"49", x"51", x"4d", x"5b", x"4b", x"34", x"57", x"69", x"77", x"73", 
        x"e8", x"e6", x"e1", x"d6", x"bb", x"ba", x"93", x"a7", x"c8", x"b6", x"c7", x"e6", x"e5", x"ea", x"e7", 
        x"eb", x"c4", x"94", x"76", x"a2", x"ac", x"c8", x"bc", x"97", x"8f", x"9b", x"95", x"96", x"98", x"90", 
        x"8e", x"9b", x"94", x"ab", x"bc", x"a5", x"b8", x"ab", x"bf", x"b3", x"7d", x"6e", x"94", x"79", x"85", 
        x"76", x"74", x"75", x"77", x"87", x"69", x"6d", x"8f", x"6f", x"58", x"76", x"60", x"67", x"85", x"8c", 
        x"9d", x"83", x"6d", x"94", x"9a", x"ab", x"db", x"c9", x"99", x"9d", x"9d", x"a2", x"9c", x"9d", x"9b", 
        x"99", x"9b", x"9c", x"9e", x"9c", x"98", x"98", x"9b", x"a0", x"a1", x"9e", x"52", x"2c", x"66", x"56", 
        x"42", x"67", x"7f", x"80", x"87", x"b8", x"d7", x"a9", x"a8", x"bb", x"c9", x"d7", x"e5", x"f0", x"f5", 
        x"f5", x"f3", x"df", x"83", x"2c", x"31", x"2e", x"29", x"22", x"15", x"08", x"04", x"08", x"16", x"2c", 
        x"41", x"70", x"8e", x"9b", x"a8", x"b0", x"b0", x"b9", x"a9", x"58", x"46", x"2c", x"4a", x"c9", x"e2", 
        x"dd", x"de", x"dd", x"d5", x"cc", x"c4", x"b9", x"b7", x"a1", x"6c", x"6f", x"6d", x"89", x"9c", x"90", 
        x"91", x"7f", x"6c", x"cc", x"db", x"d6", x"d7", x"d3", x"d7", x"da", x"ce", x"d1", x"d1", x"d1", x"d5", 
        x"d4", x"d1", x"d0", x"d1", x"d2", x"d3", x"d2", x"d2", x"d2", x"d3", x"d4", x"d5", x"d4", x"d1", x"d1", 
        x"d3", x"d2", x"d2", x"d3", x"d4", x"d4", x"d5", x"d5", x"d2", x"d0", x"d2", x"d3", x"d3", x"d2", x"d2", 
        x"d2", x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", x"d4", x"d3", x"d4", x"d6", x"d6", x"d1", x"d3", x"d2", 
        x"d4", x"d5", x"d4", x"de", x"f1", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"ef", x"ee", x"ee", 
        x"ee", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ee", x"ee", x"ee", 
        x"ef", x"ef", x"f0", x"ef", x"ed", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", 
        x"e8", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f0", x"f0", x"f1", x"f3", x"f4", x"f3", x"f1", x"f2", x"f2", 
        x"ed", x"f1", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"f5", x"f8", x"f9", x"f8", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f3", x"f4", x"f2", 
        x"f1", x"f0", x"f0", x"f3", x"f6", x"f7", x"f5", x"f4", x"f4", x"f4", x"f3", x"ef", x"e8", x"df", x"d9", 
        x"d2", x"cd", x"ca", x"c8", x"c6", x"c9", x"cd", x"ce", x"cd", x"ce", x"d0", x"d7", x"d7", x"dd", x"e4", 
        x"e8", x"ed", x"f0", x"f4", x"f4", x"f5", x"f4", x"f5", x"f3", x"ef", x"ef", x"f1", x"f0", x"f2", x"f1", 
        x"ee", x"f2", x"f1", x"ef", x"f0", x"ef", x"f1", x"f1", x"f0", x"f1", x"ef", x"f1", x"f5", x"f6", x"f7", 
        x"f7", x"f6", x"f7", x"f8", x"c2", x"64", x"44", x"86", x"d4", x"d6", x"d5", x"d5", x"db", x"c1", x"98", 
        x"9d", x"9f", x"9d", x"9d", x"99", x"98", x"98", x"98", x"97", x"96", x"95", x"98", x"98", x"96", x"98", 
        x"99", x"94", x"90", x"88", x"85", x"7f", x"75", x"72", x"73", x"53", x"3e", x"47", x"66", x"6b", x"6e", 
        x"77", x"82", x"8b", x"8f", x"90", x"85", x"79", x"76", x"75", x"74", x"73", x"72", x"72", x"73", x"64", 
        x"62", x"75", x"71", x"6d", x"6d", x"6b", x"6e", x"6f", x"68", x"67", x"6f", x"57", x"46", x"4a", x"73", 
        x"89", x"85", x"83", x"83", x"82", x"80", x"80", x"7e", x"7b", x"7e", x"7e", x"7d", x"7b", x"75", x"71", 
        x"73", x"72", x"6d", x"6c", x"4d", x"52", x"66", x"61", x"5a", x"55", x"52", x"54", x"52", x"53", x"5e", 
        x"64", x"69", x"66", x"45", x"55", x"93", x"b8", x"ca", x"d5", x"d8", x"d3", x"d4", x"ce", x"c4", x"b0", 
        x"7c", x"69", x"61", x"3b", x"39", x"3e", x"36", x"32", x"2b", x"35", x"41", x"3a", x"39", x"62", x"70", 
        x"7a", x"86", x"91", x"86", x"79", x"7e", x"82", x"84", x"8a", x"66", x"3c", x"62", x"75", x"6f", x"5f", 
        x"e0", x"e4", x"d2", x"d7", x"cc", x"b4", x"92", x"8f", x"b8", x"a8", x"cf", x"e4", x"e6", x"e3", x"ce", 
        x"cf", x"bf", x"c0", x"97", x"a9", x"ba", x"be", x"b7", x"af", x"a4", x"84", x"94", x"97", x"90", x"92", 
        x"9b", x"9b", x"72", x"78", x"82", x"7e", x"94", x"a3", x"b6", x"ba", x"a1", x"6f", x"8e", x"70", x"7a", 
        x"96", x"89", x"7d", x"83", x"80", x"6c", x"60", x"6c", x"7f", x"5d", x"77", x"88", x"91", x"92", x"a3", 
        x"9f", x"71", x"8a", x"a8", x"c0", x"b7", x"d9", x"ad", x"81", x"98", x"a3", x"aa", x"ad", x"af", x"ae", 
        x"a6", x"9e", x"a3", x"9c", x"9b", x"94", x"95", x"9e", x"a2", x"9d", x"9d", x"8e", x"74", x"8b", x"62", 
        x"45", x"66", x"6a", x"3d", x"50", x"ab", x"db", x"90", x"88", x"8e", x"8a", x"8a", x"93", x"9f", x"a7", 
        x"bd", x"d5", x"d4", x"a9", x"7d", x"7c", x"6b", x"57", x"2f", x"0d", x"19", x"29", x"36", x"4e", x"63", 
        x"68", x"71", x"66", x"61", x"6c", x"69", x"5f", x"66", x"62", x"4e", x"4c", x"2f", x"42", x"79", x"8a", 
        x"93", x"97", x"a1", x"aa", x"af", x"b8", x"bb", x"ba", x"a6", x"6f", x"6d", x"6c", x"8b", x"a3", x"99", 
        x"94", x"77", x"6b", x"cd", x"dd", x"d6", x"d7", x"d7", x"d5", x"d9", x"ce", x"d1", x"d1", x"d0", x"d3", 
        x"d4", x"d1", x"cf", x"cf", x"d1", x"d2", x"d3", x"d2", x"d2", x"d3", x"d3", x"d4", x"d2", x"d0", x"d0", 
        x"d3", x"d2", x"d2", x"d2", x"d3", x"d4", x"d5", x"d6", x"d3", x"d1", x"d2", x"d4", x"d4", x"d3", x"d3", 
        x"d2", x"d1", x"d1", x"d0", x"cf", x"cf", x"d2", x"d4", x"d4", x"d3", x"d6", x"d6", x"d2", x"d4", x"d3", 
        x"d3", x"d3", x"d3", x"dd", x"f2", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"f0", x"ef", x"ee", 
        x"ee", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ee", x"ee", x"ee", 
        x"ee", x"ed", x"ee", x"ed", x"ed", x"ee", x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f0", x"ef", x"ef", x"f0", x"f2", 
        x"e8", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f1", x"f0", x"f0", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"ec", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f7", x"f9", x"f9", x"f8", x"f4", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f3", x"f3", x"f2", x"f0", x"f0", x"f2", x"f3", x"f2", x"f0", x"f0", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"ef", x"e9", x"e6", x"e2", x"db", x"d3", x"ce", x"c6", x"c7", x"c1", x"c1", x"c1", 
        x"c4", x"c9", x"cd", x"d1", x"d3", x"d7", x"de", x"e4", x"ec", x"f1", x"f3", x"f2", x"f2", x"f4", x"f2", 
        x"f0", x"f0", x"ef", x"ee", x"f0", x"ef", x"f1", x"f1", x"f0", x"f1", x"ef", x"ef", x"f4", x"f6", x"f7", 
        x"f8", x"f6", x"f7", x"fa", x"c6", x"67", x"47", x"7f", x"d3", x"d9", x"d6", x"d7", x"d9", x"c2", x"9a", 
        x"9e", x"a0", x"9c", x"9c", x"9e", x"9c", x"9c", x"9d", x"9e", x"9b", x"95", x"8e", x"89", x"80", x"7a", 
        x"78", x"71", x"74", x"73", x"74", x"77", x"77", x"75", x"79", x"5f", x"44", x"52", x"81", x"91", x"90", 
        x"8d", x"8e", x"91", x"8f", x"8c", x"7e", x"70", x"6e", x"6c", x"67", x"63", x"61", x"5f", x"62", x"55", 
        x"4d", x"6e", x"71", x"6c", x"70", x"79", x"80", x"87", x"89", x"89", x"92", x"6f", x"4b", x"51", x"70", 
        x"85", x"84", x"82", x"80", x"7d", x"79", x"77", x"71", x"69", x"6a", x"6a", x"69", x"6a", x"6a", x"6a", 
        x"67", x"65", x"5f", x"5c", x"39", x"3b", x"58", x"5e", x"68", x"69", x"6a", x"70", x"73", x"7d", x"8a", 
        x"8d", x"98", x"93", x"5d", x"50", x"92", x"a9", x"a8", x"a4", x"a0", x"99", x"9c", x"9a", x"96", x"88", 
        x"4d", x"33", x"35", x"28", x"2d", x"43", x"44", x"50", x"62", x"86", x"94", x"80", x"66", x"9b", x"9e", 
        x"9c", x"97", x"96", x"83", x"72", x"6e", x"69", x"60", x"60", x"4d", x"30", x"50", x"62", x"67", x"5c", 
        x"a4", x"d0", x"db", x"e9", x"e6", x"ac", x"79", x"5d", x"87", x"b8", x"d4", x"df", x"cf", x"c6", x"b6", 
        x"c3", x"da", x"c8", x"96", x"b6", x"ad", x"ac", x"d3", x"d0", x"ca", x"b7", x"d3", x"af", x"8c", x"90", 
        x"a1", x"8d", x"7a", x"78", x"6d", x"7b", x"80", x"a2", x"a8", x"9e", x"8f", x"62", x"8f", x"88", x"62", 
        x"78", x"76", x"6a", x"77", x"7f", x"8b", x"7f", x"65", x"83", x"62", x"55", x"5d", x"68", x"7d", x"95", 
        x"87", x"65", x"81", x"a8", x"c3", x"a7", x"c3", x"85", x"3c", x"5a", x"74", x"5a", x"6e", x"8b", x"93", 
        x"9c", x"a2", x"ab", x"b2", x"b2", x"9e", x"95", x"9c", x"9c", x"9a", x"96", x"aa", x"ad", x"a4", x"97", 
        x"9b", x"98", x"8e", x"7c", x"7f", x"b5", x"de", x"9d", x"9f", x"ab", x"a8", x"a1", x"94", x"85", x"7f", 
        x"85", x"93", x"9b", x"9f", x"ac", x"b9", x"bb", x"b5", x"63", x"2e", x"71", x"a0", x"9f", x"9c", x"90", 
        x"80", x"77", x"76", x"71", x"76", x"66", x"56", x"54", x"48", x"51", x"51", x"30", x"3b", x"48", x"4e", 
        x"57", x"56", x"57", x"5b", x"60", x"66", x"6d", x"70", x"74", x"6b", x"6c", x"6f", x"81", x"8b", x"7a", 
        x"6a", x"43", x"5b", x"ce", x"dd", x"d7", x"d8", x"d9", x"d4", x"d8", x"cd", x"d1", x"d1", x"d0", x"d1", 
        x"d3", x"d1", x"ce", x"ce", x"d0", x"d2", x"d3", x"d4", x"d2", x"d2", x"d2", x"d3", x"d2", x"d1", x"d1", 
        x"d2", x"d3", x"d3", x"d2", x"d2", x"d4", x"d5", x"d7", x"d4", x"d2", x"d3", x"d5", x"d4", x"d4", x"d4", 
        x"d3", x"d2", x"d1", x"d1", x"d1", x"d1", x"d2", x"d5", x"d4", x"d3", x"d5", x"d5", x"d2", x"d5", x"d3", 
        x"d2", x"d2", x"d2", x"de", x"f3", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"f1", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", 
        x"ed", x"ed", x"ec", x"ec", x"ee", x"ee", x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"e8", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f4", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", 
        x"ec", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", 
        x"f3", x"f8", x"fa", x"f9", x"f7", x"f4", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f0", x"ef", x"f1", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f0", x"f2", x"f4", x"f3", x"f1", x"f0", x"f0", x"f2", 
        x"f1", x"f2", x"f5", x"f6", x"f6", x"f8", x"f9", x"f4", x"f1", x"ef", x"e9", x"e9", x"e4", x"e1", x"d9", 
        x"d6", x"d2", x"cb", x"c7", x"c2", x"c1", x"c1", x"c1", x"c4", x"c8", x"ca", x"cd", x"d3", x"dd", x"e0", 
        x"ea", x"ef", x"f2", x"f1", x"f3", x"f2", x"f4", x"f2", x"f1", x"f2", x"ef", x"f0", x"f5", x"f7", x"f8", 
        x"f7", x"f5", x"f6", x"fa", x"c9", x"6a", x"49", x"7b", x"ce", x"d6", x"d4", x"d9", x"dc", x"c9", x"a5", 
        x"a6", x"a5", x"9e", x"99", x"92", x"8c", x"85", x"7e", x"78", x"75", x"72", x"6f", x"5e", x"73", x"75", 
        x"78", x"7c", x"85", x"8d", x"8f", x"93", x"98", x"95", x"95", x"73", x"4b", x"51", x"82", x"95", x"92", 
        x"87", x"7f", x"7b", x"77", x"74", x"66", x"5c", x"60", x"60", x"5c", x"5d", x"5f", x"62", x"6d", x"61", 
        x"53", x"80", x"86", x"82", x"84", x"87", x"86", x"88", x"86", x"8b", x"98", x"7a", x"4c", x"4b", x"62", 
        x"74", x"6c", x"69", x"69", x"69", x"68", x"6c", x"6d", x"6a", x"68", x"62", x"59", x"55", x"59", x"5d", 
        x"57", x"66", x"6c", x"73", x"58", x"56", x"7a", x"85", x"8c", x"90", x"94", x"9a", x"94", x"8d", x"85", 
        x"76", x"6e", x"60", x"3d", x"35", x"61", x"7b", x"87", x"8f", x"95", x"9b", x"a9", x"b4", x"be", x"b4", 
        x"6f", x"59", x"69", x"53", x"54", x"79", x"77", x"79", x"84", x"98", x"98", x"79", x"53", x"77", x"71", 
        x"6d", x"64", x"65", x"5d", x"53", x"4f", x"4c", x"4a", x"4d", x"44", x"29", x"43", x"59", x"68", x"68", 
        x"a3", x"ae", x"aa", x"b0", x"c1", x"af", x"7e", x"3c", x"8d", x"d6", x"be", x"dc", x"d7", x"d4", x"d6", 
        x"d6", x"b6", x"ca", x"d8", x"e0", x"9e", x"a3", x"ee", x"f0", x"c8", x"9a", x"af", x"9e", x"8f", x"87", 
        x"89", x"7c", x"7b", x"86", x"88", x"84", x"97", x"80", x"78", x"89", x"72", x"6c", x"91", x"70", x"67", 
        x"65", x"7f", x"75", x"75", x"74", x"72", x"7e", x"6d", x"7a", x"7a", x"68", x"63", x"6a", x"75", x"6d", 
        x"6d", x"6f", x"6d", x"7c", x"70", x"6d", x"a6", x"92", x"63", x"74", x"74", x"42", x"4d", x"7b", x"48", 
        x"41", x"73", x"68", x"61", x"76", x"92", x"92", x"9c", x"9e", x"9d", x"92", x"9c", x"b3", x"a1", x"a5", 
        x"bb", x"a5", x"a4", x"b7", x"98", x"b6", x"d9", x"69", x"47", x"79", x"6d", x"71", x"88", x"9a", x"a6", 
        x"a0", x"97", x"8e", x"90", x"96", x"96", x"90", x"93", x"46", x"30", x"91", x"ce", x"d2", x"d8", x"d6", 
        x"d3", x"d4", x"d2", x"cb", x"c2", x"b9", x"b6", x"b4", x"95", x"68", x"56", x"34", x"3c", x"6c", x"75", 
        x"76", x"6e", x"62", x"5f", x"59", x"4d", x"56", x"65", x"6c", x"6b", x"5a", x"47", x"35", x"2c", x"28", 
        x"26", x"16", x"53", x"d0", x"dc", x"d6", x"d6", x"d7", x"d6", x"d9", x"cc", x"d0", x"d1", x"d0", x"d2", 
        x"d3", x"d1", x"d0", x"d0", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d2", x"d3", x"d2", x"d1", x"d2", 
        x"d3", x"d3", x"d3", x"d3", x"d3", x"d4", x"d5", x"d5", x"d4", x"d3", x"d4", x"d4", x"d4", x"d4", x"d5", 
        x"d4", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d5", x"d4", x"d3", x"d4", x"d5", x"d2", x"d7", x"d6", 
        x"d4", x"d3", x"d2", x"dc", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"f0", x"ef", x"f1", x"f0", x"f0", 
        x"ef", x"f1", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ee", 
        x"ee", x"ee", x"ed", x"ed", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"e9", x"f1", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"f1", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", 
        x"ec", x"ef", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f1", x"f0", x"f1", x"f2", 
        x"f4", x"f9", x"f9", x"f8", x"f6", x"f4", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f0", x"f1", x"f4", 
        x"f4", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"ed", x"ee", 
        x"ef", x"f3", x"f7", x"f8", x"f5", x"f5", x"f5", x"f3", x"f1", x"f3", x"ed", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f2", x"ef", x"ed", x"e7", x"e6", x"e3", x"e0", x"dc", x"d6", x"cd", x"c5", x"c1", x"bb", x"b4", 
        x"b5", x"b4", x"ba", x"c4", x"d0", x"db", x"e3", x"e6", x"ea", x"ef", x"f1", x"f4", x"f4", x"f4", x"f7", 
        x"f7", x"f5", x"f6", x"f9", x"ce", x"6d", x"46", x"76", x"cc", x"db", x"db", x"d3", x"cb", x"b3", x"89", 
        x"80", x"7c", x"78", x"75", x"76", x"78", x"7b", x"7f", x"83", x"8a", x"90", x"84", x"5c", x"91", x"95", 
        x"95", x"97", x"96", x"97", x"97", x"95", x"95", x"94", x"91", x"6d", x"4c", x"4a", x"64", x"6f", x"6f", 
        x"6b", x"70", x"71", x"79", x"7d", x"74", x"6b", x"70", x"71", x"6e", x"72", x"73", x"73", x"78", x"6b", 
        x"5d", x"84", x"8b", x"89", x"88", x"87", x"7f", x"7a", x"75", x"71", x"74", x"5e", x"38", x"40", x"5a", 
        x"78", x"72", x"6f", x"6a", x"64", x"5f", x"5c", x"5c", x"5d", x"62", x"6c", x"76", x"7f", x"88", x"84", 
        x"70", x"93", x"9c", x"a0", x"7d", x"6b", x"81", x"80", x"70", x"61", x"56", x"58", x"4e", x"49", x"48", 
        x"40", x"3a", x"34", x"2d", x"38", x"65", x"96", x"b5", x"c1", x"c9", x"d0", x"d6", x"dc", x"e0", x"ce", 
        x"8c", x"73", x"7a", x"56", x"4b", x"64", x"57", x"5b", x"58", x"5c", x"5f", x"51", x"31", x"53", x"51", 
        x"53", x"56", x"62", x"63", x"5e", x"61", x"68", x"71", x"77", x"67", x"39", x"51", x"6a", x"7e", x"84", 
        x"b9", x"bd", x"c9", x"b6", x"b0", x"b4", x"84", x"4c", x"91", x"a3", x"ad", x"cc", x"d8", x"dc", x"e4", 
        x"d6", x"bd", x"e2", x"eb", x"ed", x"c6", x"ac", x"c2", x"d0", x"cb", x"9b", x"81", x"92", x"91", x"70", 
        x"7b", x"7a", x"82", x"7f", x"7a", x"86", x"b8", x"7f", x"64", x"70", x"6f", x"89", x"78", x"6e", x"7e", 
        x"5d", x"6c", x"6d", x"65", x"64", x"6d", x"73", x"70", x"75", x"93", x"a3", x"8e", x"71", x"8a", x"8c", 
        x"7f", x"72", x"79", x"85", x"8c", x"90", x"a9", x"b3", x"92", x"a2", x"8f", x"6f", x"69", x"7f", x"51", 
        x"56", x"8d", x"65", x"2e", x"38", x"8c", x"94", x"99", x"9d", x"98", x"94", x"a1", x"ad", x"a0", x"a3", 
        x"b7", x"a2", x"a5", x"c0", x"8f", x"ab", x"d9", x"62", x"38", x"83", x"42", x"2b", x"46", x"4e", x"57", 
        x"70", x"9a", x"a0", x"a0", x"9e", x"9d", x"94", x"90", x"3f", x"36", x"76", x"a2", x"a4", x"a4", x"a1", 
        x"ac", x"b5", x"c5", x"d2", x"cd", x"d6", x"e1", x"e4", x"c8", x"72", x"52", x"31", x"43", x"b5", x"cf", 
        x"c5", x"bb", x"b3", x"b4", x"ae", x"96", x"80", x"65", x"41", x"2f", x"26", x"23", x"1b", x"16", x"16", 
        x"17", x"1b", x"5c", x"d3", x"df", x"d8", x"d4", x"d6", x"d9", x"db", x"cc", x"d0", x"d1", x"d1", x"d2", 
        x"d2", x"d1", x"d1", x"d2", x"d3", x"d2", x"d1", x"d3", x"d3", x"d3", x"d2", x"d3", x"d3", x"d1", x"d2", 
        x"d3", x"d3", x"d2", x"d3", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d4", x"d2", x"d2", x"d3", x"d6", 
        x"d5", x"d3", x"d2", x"d1", x"d1", x"d2", x"d2", x"d4", x"d4", x"d2", x"d3", x"d4", x"d3", x"d7", x"d5", 
        x"d5", x"d4", x"d4", x"dd", x"f1", x"ef", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ed", x"ee", 
        x"ee", x"ee", x"ee", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", 
        x"f0", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f1", x"f2", x"f2", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", 
        x"e9", x"f2", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"f1", x"f0", x"ef", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", 
        x"ec", x"ef", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f3", x"f1", x"ef", x"f0", x"f2", 
        x"f4", x"fa", x"fa", x"f8", x"f6", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f2", x"ef", x"f0", x"f2", x"f2", x"ef", x"ef", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f3", 
        x"f4", x"f4", x"f6", x"f7", x"f5", x"f7", x"f6", x"f0", x"f0", x"f2", x"eb", x"f0", x"f1", x"f1", x"ee", 
        x"ef", x"f0", x"f0", x"f2", x"f0", x"f2", x"f3", x"f3", x"f1", x"ee", x"ec", x"eb", x"e8", x"e5", x"df", 
        x"dd", x"d4", x"ce", x"c7", x"c7", x"c2", x"c0", x"be", x"be", x"c5", x"cc", x"d3", x"db", x"e3", x"e9", 
        x"ed", x"ef", x"f0", x"f1", x"ca", x"6d", x"48", x"6a", x"a3", x"a3", x"a2", x"9d", x"a1", x"97", x"7f", 
        x"84", x"8f", x"96", x"97", x"98", x"98", x"98", x"99", x"99", x"99", x"9a", x"91", x"63", x"96", x"97", 
        x"95", x"8d", x"88", x"81", x"80", x"7a", x"6f", x"71", x"73", x"5b", x"44", x"44", x"68", x"81", x"8a", 
        x"88", x"8b", x"88", x"8b", x"8f", x"83", x"73", x"72", x"72", x"71", x"73", x"73", x"75", x"75", x"6a", 
        x"5b", x"72", x"72", x"6a", x"66", x"6a", x"69", x"6b", x"75", x"79", x"7a", x"60", x"38", x"43", x"4b", 
        x"68", x"67", x"69", x"6d", x"76", x"83", x"8a", x"8d", x"90", x"93", x"98", x"99", x"92", x"8c", x"79", 
        x"53", x"6e", x"65", x"5f", x"49", x"3f", x"55", x"4d", x"4e", x"48", x"42", x"44", x"41", x"4b", x"54", 
        x"5c", x"68", x"67", x"4d", x"45", x"84", x"b0", x"c6", x"c5", x"c2", x"bd", x"b5", x"b1", x"a7", x"92", 
        x"6b", x"5a", x"5b", x"44", x"39", x"4d", x"48", x"47", x"4b", x"60", x"70", x"6d", x"40", x"7a", x"86", 
        x"86", x"8c", x"93", x"8b", x"7e", x"7f", x"81", x"79", x"76", x"64", x"35", x"4a", x"58", x"5d", x"62", 
        x"9b", x"c7", x"e2", x"c7", x"d7", x"ce", x"88", x"5a", x"a0", x"a6", x"c1", x"be", x"b9", x"b6", x"b7", 
        x"a6", x"ba", x"cf", x"d2", x"de", x"c2", x"b0", x"ad", x"a2", x"a7", x"94", x"75", x"6f", x"79", x"82", 
        x"88", x"8e", x"7a", x"94", x"7e", x"96", x"a3", x"7f", x"68", x"63", x"7b", x"91", x"72", x"82", x"93", 
        x"7e", x"69", x"5a", x"4c", x"58", x"70", x"86", x"7f", x"71", x"71", x"9f", x"98", x"64", x"81", x"80", 
        x"86", x"7e", x"78", x"84", x"a3", x"9d", x"9b", x"9e", x"9f", x"cc", x"cb", x"c4", x"b9", x"a7", x"9f", 
        x"92", x"8a", x"87", x"51", x"40", x"85", x"91", x"9b", x"9e", x"98", x"95", x"a6", x"ac", x"a2", x"ac", 
        x"c5", x"a9", x"a5", x"c7", x"a1", x"b0", x"d8", x"69", x"59", x"90", x"4b", x"4d", x"68", x"6c", x"7f", 
        x"7c", x"9d", x"9e", x"9e", x"a1", x"a0", x"a3", x"a0", x"4e", x"5c", x"7d", x"9f", x"9e", x"9e", x"9c", 
        x"9a", x"93", x"a1", x"c8", x"a3", x"87", x"a3", x"ba", x"b4", x"6e", x"55", x"2e", x"47", x"c8", x"ea", 
        x"e0", x"d4", x"bb", x"99", x"70", x"4d", x"35", x"26", x"1d", x"18", x"12", x"14", x"1d", x"2f", x"45", 
        x"59", x"64", x"85", x"d4", x"dc", x"d8", x"d4", x"d4", x"d8", x"dc", x"ce", x"d2", x"d2", x"d0", x"d2", 
        x"d3", x"d4", x"d4", x"d3", x"d4", x"d1", x"d1", x"d3", x"d5", x"d3", x"d1", x"d2", x"d2", x"d1", x"d4", 
        x"d4", x"d3", x"d2", x"d2", x"d3", x"d4", x"d6", x"d5", x"d4", x"d6", x"d6", x"d2", x"d1", x"d5", x"d7", 
        x"d3", x"d3", x"d2", x"d0", x"d2", x"d3", x"d4", x"d4", x"d7", x"d0", x"d2", x"d5", x"d3", x"d7", x"d4", 
        x"d4", x"d3", x"d1", x"db", x"f2", x"ee", x"ed", x"ef", x"ef", x"ec", x"ec", x"ec", x"ed", x"ef", x"ee", 
        x"ed", x"ec", x"ee", x"f0", x"f1", x"ef", x"ee", x"ee", x"ec", x"ee", x"ef", x"ef", x"f1", x"ef", x"ee", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f2", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"ee", x"f0", x"ef", x"ee", x"ef", x"ee", x"ee", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f1", x"f2", x"f2", 
        x"f1", x"ef", x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", x"f1", x"f2", 
        x"e9", x"f2", x"f2", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f0", x"f1", x"f1", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", 
        x"ee", x"f0", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f3", x"f2", x"f3", x"f4", x"f3", x"f4", 
        x"f7", x"fa", x"f9", x"f6", x"f4", x"f2", x"f2", x"f2", x"f3", x"f3", x"f1", x"f1", x"f2", x"f2", x"f1", 
        x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", 
        x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f4", 
        x"f3", x"f3", x"f6", x"f7", x"f6", x"f5", x"f3", x"f0", x"f0", x"f1", x"eb", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"ef", x"ed", x"ee", x"ed", x"ed", x"eb", x"ea", x"e3", x"dd", x"d5", x"cc", x"c2", x"b4", x"b5", x"b1", 
        x"a7", x"ac", x"b2", x"b1", x"95", x"53", x"40", x"58", x"9e", x"c1", x"ca", x"d0", x"d7", x"cc", x"a3", 
        x"9d", x"a1", x"9f", x"9f", x"a2", x"9e", x"a0", x"9d", x"98", x"95", x"94", x"88", x"5d", x"74", x"75", 
        x"6d", x"6c", x"6c", x"6e", x"75", x"80", x"87", x"8a", x"93", x"7c", x"4b", x"4b", x"78", x"91", x"95", 
        x"8f", x"8b", x"8b", x"8c", x"92", x"88", x"76", x"71", x"69", x"67", x"60", x"5f", x"5c", x"58", x"59", 
        x"46", x"65", x"72", x"76", x"73", x"6f", x"6e", x"69", x"62", x"64", x"6a", x"69", x"3d", x"48", x"59", 
        x"95", x"9f", x"a1", x"a1", x"9e", x"98", x"8a", x"7a", x"6e", x"66", x"5d", x"54", x"4d", x"4f", x"4e", 
        x"34", x"4c", x"4e", x"4e", x"42", x"31", x"4d", x"51", x"56", x"58", x"64", x"69", x"6a", x"77", x"80", 
        x"81", x"7c", x"78", x"58", x"42", x"6b", x"82", x"8c", x"88", x"89", x"8e", x"95", x"9d", x"aa", x"a9", 
        x"6c", x"4c", x"54", x"45", x"33", x"5c", x"61", x"66", x"6f", x"8f", x"9f", x"9b", x"58", x"92", x"9b", 
        x"93", x"89", x"7f", x"72", x"62", x"57", x"5b", x"5c", x"5f", x"55", x"30", x"4f", x"71", x"77", x"6f", 
        x"a9", x"bb", x"c5", x"b3", x"cc", x"e0", x"9d", x"85", x"d3", x"d4", x"e5", x"df", x"dc", x"ce", x"d4", 
        x"dd", x"d1", x"c3", x"bc", x"a7", x"a2", x"ac", x"94", x"8b", x"77", x"7b", x"8a", x"87", x"75", x"87", 
        x"a6", x"99", x"80", x"8c", x"7c", x"73", x"8f", x"96", x"6e", x"7a", x"7a", x"7d", x"57", x"5b", x"60", 
        x"7e", x"54", x"53", x"68", x"74", x"77", x"72", x"7d", x"86", x"67", x"7b", x"7f", x"7c", x"86", x"8c", 
        x"8b", x"93", x"91", x"87", x"8b", x"b3", x"c3", x"b9", x"bf", x"d0", x"dc", x"da", x"d3", x"d1", x"dd", 
        x"e0", x"db", x"da", x"c0", x"a8", x"9f", x"8f", x"92", x"8e", x"8c", x"84", x"98", x"a0", x"9a", x"a5", 
        x"bd", x"a7", x"a5", x"c7", x"a4", x"ae", x"d6", x"75", x"98", x"a8", x"55", x"60", x"78", x"9a", x"a9", 
        x"7e", x"9a", x"9b", x"9b", x"9c", x"9d", x"a0", x"97", x"5a", x"66", x"82", x"a9", x"a7", x"a5", x"a4", 
        x"9e", x"9b", x"ad", x"de", x"a5", x"6d", x"7c", x"76", x"70", x"62", x"59", x"34", x"47", x"9f", x"a5", 
        x"7e", x"5b", x"40", x"31", x"1d", x"1c", x"1b", x"19", x"21", x"31", x"49", x"62", x"76", x"81", x"86", 
        x"89", x"80", x"89", x"d1", x"d9", x"d3", x"d2", x"d5", x"d7", x"dc", x"cd", x"d2", x"d1", x"d1", x"d2", 
        x"d1", x"d3", x"d3", x"d2", x"d3", x"d0", x"d2", x"d3", x"d4", x"d2", x"d1", x"d3", x"d1", x"d0", x"d2", 
        x"d1", x"d2", x"d3", x"d3", x"d3", x"d2", x"d3", x"d5", x"d4", x"d4", x"d6", x"d7", x"d5", x"d5", x"d8", 
        x"d5", x"d6", x"d6", x"d2", x"d4", x"d5", x"d7", x"d3", x"d6", x"d5", x"d9", x"da", x"d5", x"d5", x"d2", 
        x"d4", x"d6", x"d3", x"da", x"ee", x"eb", x"ed", x"ee", x"ee", x"ed", x"ee", x"ee", x"ec", x"ee", x"ee", 
        x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", x"ed", x"ed", x"ed", x"f1", x"ef", x"ee", 
        x"ef", x"f0", x"ef", x"ee", x"f1", x"f1", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"f1", x"f0", x"ee", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f0", x"ef", x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", x"f1", x"f2", 
        x"e9", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"ef", x"ef", x"f0", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f2", 
        x"ef", x"f0", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f4", x"f4", x"f3", x"f3", x"f4", x"f3", x"f4", 
        x"f8", x"f9", x"f6", x"f4", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f3", x"f2", x"f1", x"f1", x"f1", x"f4", 
        x"f2", x"f2", x"f5", x"f7", x"f5", x"f3", x"f1", x"ef", x"f0", x"f1", x"eb", x"f0", x"f0", x"ef", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"ef", x"f1", x"f2", x"ec", x"f0", x"eb", x"de", x"d9", x"ce", x"c6", x"b0", x"a0", x"aa", x"b4", x"b7", 
        x"b7", x"c4", x"ce", x"d0", x"af", x"64", x"4c", x"58", x"8c", x"ab", x"b6", x"be", x"cb", x"c1", x"9d", 
        x"9c", x"a0", x"97", x"96", x"90", x"89", x"87", x"7e", x"74", x"6f", x"70", x"72", x"50", x"7c", x"8b", 
        x"8c", x"95", x"98", x"96", x"94", x"93", x"92", x"8e", x"95", x"80", x"49", x"46", x"73", x"8e", x"95", 
        x"93", x"86", x"7f", x"7a", x"74", x"6d", x"59", x"57", x"5a", x"5a", x"5e", x"62", x"67", x"6a", x"6a", 
        x"48", x"5d", x"66", x"68", x"6c", x"70", x"7b", x"89", x"93", x"9b", x"aa", x"9c", x"4e", x"4d", x"5e", 
        x"85", x"74", x"6a", x"61", x"56", x"4f", x"52", x"56", x"54", x"50", x"54", x"51", x"50", x"58", x"54", 
        x"31", x"52", x"5b", x"5e", x"5f", x"4f", x"74", x"80", x"82", x"79", x"77", x"70", x"63", x"61", x"62", 
        x"5f", x"57", x"5a", x"46", x"32", x"5c", x"82", x"9a", x"a8", x"b3", x"c0", x"cd", x"ce", x"cf", x"cc", 
        x"91", x"70", x"79", x"65", x"4b", x"74", x"75", x"70", x"6a", x"7b", x"7d", x"7a", x"3b", x"61", x"69", 
        x"64", x"62", x"62", x"5f", x"58", x"55", x"58", x"54", x"56", x"54", x"33", x"3a", x"4c", x"4d", x"47", 
        x"49", x"59", x"57", x"63", x"7f", x"90", x"7b", x"6f", x"b3", x"c9", x"d7", x"d2", x"bb", x"c9", x"e8", 
        x"ed", x"f2", x"ec", x"c0", x"a8", x"c3", x"c9", x"bc", x"99", x"74", x"5f", x"88", x"99", x"64", x"62", 
        x"89", x"72", x"6a", x"69", x"75", x"7a", x"7e", x"84", x"88", x"7c", x"69", x"66", x"66", x"55", x"46", 
        x"84", x"7f", x"71", x"50", x"4c", x"5f", x"56", x"67", x"6a", x"7f", x"7a", x"6c", x"6d", x"86", x"81", 
        x"8d", x"89", x"95", x"8b", x"8c", x"b3", x"cb", x"a8", x"b2", x"c0", x"cc", x"b9", x"d4", x"d7", x"d9", 
        x"e3", x"ef", x"ee", x"ef", x"ee", x"e7", x"e1", x"d8", x"c4", x"b5", x"9f", x"8d", x"83", x"7e", x"8a", 
        x"9d", x"91", x"9b", x"b5", x"9e", x"af", x"d6", x"77", x"a5", x"a2", x"54", x"6e", x"9e", x"b0", x"a7", 
        x"83", x"9d", x"a0", x"a0", x"a2", x"9e", x"63", x"31", x"35", x"69", x"85", x"a7", x"a1", x"a7", x"b3", 
        x"ad", x"ae", x"ab", x"da", x"a4", x"76", x"8f", x"8a", x"83", x"6f", x"64", x"41", x"29", x"32", x"2b", 
        x"24", x"22", x"28", x"32", x"36", x"4c", x"57", x"63", x"79", x"84", x"8c", x"8e", x"8a", x"83", x"7b", 
        x"70", x"59", x"70", x"d1", x"dd", x"d4", x"d3", x"d5", x"d6", x"da", x"cd", x"d1", x"d1", x"d2", x"d2", 
        x"d0", x"d2", x"d2", x"d1", x"d2", x"d0", x"d1", x"d2", x"d3", x"d2", x"d3", x"d4", x"d0", x"d0", x"d2", 
        x"d1", x"d2", x"d3", x"d3", x"d3", x"d2", x"d3", x"d5", x"d7", x"d4", x"d3", x"d7", x"d7", x"d4", x"d7", 
        x"d3", x"d4", x"d4", x"d2", x"d3", x"d4", x"d5", x"d1", x"d4", x"d2", x"d4", x"d4", x"d2", x"d6", x"d5", 
        x"d6", x"d6", x"d0", x"d8", x"f0", x"ed", x"ee", x"ef", x"ec", x"ec", x"ee", x"ec", x"eb", x"ed", x"ed", 
        x"ee", x"ef", x"f0", x"f1", x"f1", x"ef", x"f1", x"f0", x"ef", x"ef", x"ee", x"ec", x"ef", x"ef", x"ee", 
        x"ee", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", x"f1", x"f2", 
        x"e9", x"f1", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f2", 
        x"ef", x"f0", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f1", 
        x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f1", x"f0", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f6", x"f3", x"f3", x"f4", x"f3", x"f4", 
        x"f8", x"f9", x"f5", x"f1", x"f0", x"f1", x"f3", x"f2", x"f3", x"f3", x"f1", x"f1", x"f2", x"f3", x"f4", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f5", 
        x"f3", x"f2", x"f4", x"f6", x"f3", x"f0", x"f0", x"f0", x"ef", x"f1", x"ec", x"ef", x"f0", x"f0", x"f0", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ee", 
        x"ef", x"f0", x"f0", x"e8", x"e9", x"b2", x"99", x"ac", x"b3", x"c9", x"be", x"a3", x"ce", x"f3", x"f5", 
        x"f5", x"f8", x"f9", x"f7", x"d9", x"7d", x"4a", x"61", x"a2", x"b2", x"9e", x"8b", x"8c", x"84", x"6c", 
        x"74", x"76", x"66", x"60", x"6b", x"72", x"81", x"89", x"92", x"99", x"9d", x"a3", x"69", x"8b", x"9d", 
        x"96", x"99", x"95", x"94", x"91", x"8e", x"90", x"8c", x"8e", x"7b", x"51", x"4b", x"64", x"73", x"6f", 
        x"6d", x"69", x"67", x"68", x"6c", x"72", x"6c", x"6c", x"6a", x"66", x"64", x"68", x"71", x"6a", x"72", 
        x"66", x"80", x"9a", x"9a", x"9b", x"93", x"86", x"7f", x"7b", x"75", x"72", x"61", x"2f", x"3a", x"3e", 
        x"5f", x"52", x"54", x"5f", x"65", x"66", x"65", x"62", x"5a", x"53", x"5b", x"5d", x"63", x"70", x"6d", 
        x"4a", x"73", x"7b", x"78", x"71", x"4f", x"63", x"62", x"5d", x"56", x"57", x"57", x"55", x"59", x"5c", 
        x"61", x"61", x"61", x"4f", x"3c", x"6e", x"95", x"aa", x"bd", x"c6", x"cb", x"d3", x"ce", x"c8", x"c1", 
        x"8d", x"6c", x"68", x"53", x"3c", x"58", x"53", x"54", x"55", x"65", x"61", x"5f", x"34", x"5e", x"65", 
        x"67", x"6a", x"6e", x"68", x"59", x"58", x"5c", x"63", x"68", x"65", x"50", x"5a", x"73", x"8e", x"97", 
        x"80", x"68", x"6f", x"60", x"49", x"48", x"44", x"32", x"51", x"73", x"80", x"7e", x"6c", x"9b", x"bd", 
        x"c8", x"d1", x"cb", x"b5", x"99", x"a1", x"9e", x"ab", x"a5", x"8b", x"a0", x"a7", x"97", x"7d", x"69", 
        x"6a", x"5b", x"67", x"63", x"53", x"5b", x"5b", x"6e", x"8c", x"74", x"66", x"5b", x"78", x"75", x"63", 
        x"73", x"84", x"81", x"5b", x"48", x"6d", x"5a", x"4e", x"5b", x"82", x"7d", x"83", x"7e", x"7d", x"89", 
        x"8b", x"7f", x"7d", x"6a", x"89", x"a0", x"b9", x"bb", x"cc", x"d0", x"d4", x"db", x"ea", x"ec", x"ea", 
        x"e8", x"ed", x"e9", x"e9", x"ea", x"ec", x"eb", x"eb", x"ee", x"ec", x"e7", x"e6", x"db", x"cc", x"c0", 
        x"b8", x"a5", x"a3", x"ac", x"97", x"ae", x"d3", x"7a", x"98", x"93", x"5d", x"87", x"ac", x"ad", x"a5", 
        x"84", x"9c", x"a1", x"a1", x"9e", x"a2", x"93", x"77", x"4b", x"65", x"82", x"91", x"7c", x"80", x"98", 
        x"90", x"8f", x"a3", x"d8", x"a8", x"83", x"95", x"8d", x"7b", x"68", x"5b", x"37", x"21", x"25", x"2f", 
        x"3a", x"50", x"72", x"9b", x"b7", x"ca", x"a5", x"8a", x"8b", x"86", x"7c", x"70", x"62", x"53", x"43", 
        x"37", x"29", x"59", x"ca", x"da", x"d4", x"d4", x"d6", x"d7", x"da", x"cc", x"d0", x"d0", x"d2", x"d1", 
        x"d0", x"d3", x"d3", x"d2", x"d2", x"d0", x"d1", x"d3", x"d4", x"d3", x"d4", x"d5", x"d1", x"d1", x"d3", 
        x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d4", x"d6", x"d8", x"d5", x"d1", x"d2", x"d4", x"d4", x"d6", 
        x"d2", x"d2", x"d3", x"d3", x"d4", x"d5", x"d3", x"d1", x"d4", x"d3", x"d5", x"d6", x"d4", x"d6", x"d7", 
        x"d9", x"dc", x"d7", x"db", x"ed", x"ec", x"ee", x"f1", x"f0", x"ef", x"ef", x"f0", x"ef", x"ee", x"ef", 
        x"f0", x"f1", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ed", x"ef", x"ef", x"ef", 
        x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"ef", x"ed", x"ef", x"ef", x"ee", x"ef", x"ef", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", x"f1", x"f2", 
        x"e9", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f2", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"ef", x"ee", x"ef", x"f1", x"f2", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"ee", x"f0", 
        x"f1", x"f2", x"f1", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", 
        x"ef", x"ee", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f6", x"f4", x"f3", x"f5", x"f5", x"f5", 
        x"f8", x"f9", x"f5", x"ef", x"ed", x"f0", x"f3", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f3", x"f4", 
        x"f3", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f2", x"f2", x"f2", x"f4", x"f7", 
        x"f5", x"f2", x"f4", x"f6", x"f3", x"f0", x"f0", x"f0", x"ef", x"f1", x"ec", x"ef", x"f0", x"f1", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"ef", x"f1", x"f4", x"ef", x"cf", x"7d", x"a2", x"e5", x"ef", x"f2", x"de", x"bb", x"d9", x"f5", x"f1", 
        x"ed", x"e6", x"e2", x"e1", x"c7", x"77", x"4c", x"56", x"94", x"ae", x"a8", x"a0", x"aa", x"ad", x"94", 
        x"92", x"90", x"84", x"81", x"79", x"79", x"7d", x"7c", x"80", x"85", x"85", x"87", x"62", x"7b", x"8f", 
        x"8d", x"8a", x"86", x"87", x"84", x"7c", x"76", x"6b", x"6c", x"5e", x"43", x"43", x"53", x"72", x"7c", 
        x"7d", x"7d", x"79", x"74", x"77", x"7c", x"82", x"8d", x"92", x"99", x"9c", x"97", x"96", x"77", x"72", 
        x"63", x"64", x"6b", x"64", x"5f", x"5a", x"54", x"51", x"55", x"5d", x"65", x"5f", x"37", x"46", x"49", 
        x"6e", x"67", x"65", x"68", x"69", x"6b", x"72", x"75", x"75", x"71", x"70", x"6f", x"70", x"72", x"69", 
        x"44", x"5d", x"60", x"58", x"51", x"39", x"54", x"5e", x"5c", x"5a", x"5c", x"5b", x"5a", x"5c", x"59", 
        x"60", x"67", x"6a", x"5b", x"43", x"72", x"9b", x"a7", x"ad", x"ad", x"a4", x"a4", x"9f", x"9e", x"9e", 
        x"72", x"58", x"5b", x"4a", x"36", x"55", x"5a", x"58", x"54", x"67", x"73", x"73", x"43", x"62", x"7b", 
        x"85", x"88", x"8f", x"90", x"88", x"8a", x"8e", x"9f", x"ad", x"b7", x"c0", x"ca", x"d2", x"da", x"d8", 
        x"8c", x"67", x"8d", x"81", x"6e", x"60", x"50", x"33", x"46", x"6b", x"6e", x"62", x"4d", x"54", x"6c", 
        x"89", x"76", x"82", x"8c", x"9e", x"9f", x"76", x"69", x"7d", x"72", x"80", x"7f", x"8f", x"90", x"7f", 
        x"61", x"61", x"72", x"62", x"53", x"47", x"51", x"79", x"6f", x"85", x"83", x"4f", x"61", x"83", x"6c", 
        x"5d", x"74", x"78", x"6a", x"44", x"45", x"44", x"5d", x"7e", x"8f", x"73", x"62", x"69", x"69", x"61", 
        x"7a", x"6d", x"7c", x"84", x"b8", x"ad", x"b5", x"d1", x"e0", x"c8", x"ad", x"d0", x"dc", x"e9", x"ed", 
        x"ec", x"ec", x"eb", x"eb", x"ec", x"ea", x"e9", x"ea", x"ed", x"e9", x"e8", x"e9", x"ee", x"f3", x"f3", 
        x"f5", x"f1", x"eb", x"e3", x"d1", x"d6", x"dd", x"b4", x"b0", x"97", x"7b", x"88", x"8c", x"97", x"91", 
        x"72", x"89", x"9b", x"9a", x"a0", x"a0", x"b7", x"c4", x"64", x"63", x"86", x"a2", x"97", x"95", x"9c", 
        x"8e", x"8d", x"a4", x"ca", x"a1", x"72", x"6e", x"5b", x"41", x"3d", x"47", x"47", x"55", x"72", x"96", 
        x"b6", x"cf", x"e0", x"e6", x"e0", x"d2", x"98", x"6e", x"61", x"51", x"43", x"35", x"29", x"2b", x"39", 
        x"49", x"4c", x"70", x"cd", x"dc", x"d6", x"d2", x"d7", x"d9", x"d9", x"cd", x"d1", x"d0", x"d1", x"cf", 
        x"d1", x"d5", x"d3", x"d2", x"d3", x"d0", x"d1", x"d3", x"d5", x"d4", x"d4", x"d6", x"d3", x"d2", x"d3", 
        x"d3", x"d4", x"d5", x"d5", x"d5", x"d5", x"d5", x"d5", x"d4", x"d2", x"d1", x"d1", x"d3", x"d5", x"d6", 
        x"d4", x"d3", x"d5", x"d6", x"d3", x"d3", x"d1", x"d3", x"d5", x"d2", x"d5", x"d9", x"d8", x"dc", x"dc", 
        x"d7", x"d1", x"c3", x"bc", x"ca", x"d6", x"db", x"e0", x"e2", x"de", x"de", x"e3", x"e6", x"e9", x"ea", 
        x"ee", x"f0", x"ee", x"ef", x"f2", x"f3", x"f1", x"f1", x"f1", x"ee", x"ed", x"ee", x"ef", x"ee", x"ef", 
        x"f0", x"ee", x"ec", x"ec", x"ee", x"ef", x"ef", x"ee", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"f2", 
        x"e9", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", x"f2", x"f1", x"ee", x"ef", x"f1", x"f2", x"f1", x"f1", x"f0", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"ee", x"ed", x"ef", 
        x"f0", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", 
        x"ef", x"ee", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f6", x"f4", x"f4", x"f6", x"f6", x"f5", 
        x"f6", x"f8", x"f4", x"ef", x"ee", x"f0", x"f3", x"f4", x"f2", x"f1", x"f2", x"f1", x"f1", x"f2", x"f3", 
        x"f3", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f2", x"f2", x"f4", x"f6", x"f8", 
        x"f6", x"f4", x"f6", x"f6", x"f2", x"f1", x"f1", x"f0", x"ee", x"f0", x"eb", x"ee", x"f0", x"f2", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"ed", x"ee", x"f1", x"ea", x"9f", x"4e", x"9c", x"e7", x"ea", x"e8", x"d0", x"ab", x"ba", x"d2", x"cc", 
        x"ca", x"c2", x"bf", x"c0", x"b1", x"70", x"49", x"52", x"a3", x"cd", x"d4", x"da", x"df", x"db", x"b0", 
        x"a5", x"a9", x"a9", x"a9", x"a5", x"9f", x"97", x"8e", x"85", x"7b", x"6a", x"5e", x"45", x"56", x"70", 
        x"6a", x"52", x"43", x"54", x"67", x"6d", x"69", x"65", x"70", x"68", x"44", x"3f", x"53", x"79", x"8c", 
        x"97", x"a1", x"a3", x"a0", x"9f", x"9d", x"96", x"8d", x"83", x"79", x"6e", x"65", x"5d", x"3c", x"3a", 
        x"33", x"37", x"4f", x"52", x"56", x"64", x"6c", x"69", x"6d", x"71", x"75", x"73", x"47", x"4f", x"4e", 
        x"7e", x"7e", x"78", x"77", x"74", x"72", x"6f", x"68", x"62", x"61", x"5d", x"5a", x"5c", x"61", x"5f", 
        x"40", x"57", x"61", x"5f", x"58", x"3f", x"50", x"58", x"56", x"55", x"5b", x"64", x"6a", x"70", x"73", 
        x"6f", x"6b", x"6a", x"5a", x"38", x"54", x"78", x"87", x"8e", x"96", x"9f", x"b1", x"bb", x"c4", x"ce", 
        x"8e", x"53", x"55", x"3f", x"27", x"46", x"51", x"55", x"63", x"86", x"95", x"92", x"79", x"8f", x"a7", 
        x"b6", x"b9", x"c2", x"cc", x"d1", x"d8", x"db", x"e3", x"e0", x"da", x"da", x"da", x"d7", x"d8", x"d4", 
        x"99", x"7c", x"8a", x"7c", x"76", x"61", x"67", x"50", x"72", x"78", x"81", x"aa", x"ac", x"95", x"8c", 
        x"8c", x"6c", x"64", x"59", x"7d", x"8c", x"6e", x"5c", x"6e", x"56", x"6b", x"84", x"88", x"84", x"51", 
        x"57", x"7a", x"60", x"46", x"55", x"7b", x"69", x"6d", x"8c", x"88", x"6a", x"5c", x"61", x"69", x"77", 
        x"62", x"63", x"81", x"6d", x"46", x"40", x"3e", x"4b", x"66", x"5e", x"5e", x"63", x"5e", x"58", x"6a", 
        x"78", x"76", x"7a", x"9f", x"bf", x"b1", x"c5", x"bf", x"c6", x"b5", x"c1", x"cf", x"e4", x"ef", x"ed", 
        x"eb", x"ec", x"ec", x"ed", x"ed", x"e7", x"ea", x"eb", x"ed", x"ef", x"ec", x"eb", x"ec", x"eb", x"ea", 
        x"ec", x"ec", x"ec", x"ee", x"e7", x"ec", x"ed", x"f1", x"e6", x"da", x"d6", x"c9", x"b7", x"b1", x"a2", 
        x"96", x"9d", x"92", x"8b", x"8c", x"88", x"9c", x"b2", x"5b", x"62", x"89", x"ad", x"b3", x"b2", x"aa", 
        x"96", x"89", x"6a", x"53", x"3d", x"2c", x"39", x"4e", x"64", x"85", x"a3", x"b7", x"cb", x"d8", x"e0", 
        x"df", x"d5", x"c1", x"a8", x"86", x"64", x"40", x"36", x"35", x"3a", x"41", x"4e", x"5c", x"65", x"6a", 
        x"70", x"73", x"7d", x"c7", x"dc", x"d8", x"d5", x"d8", x"da", x"d7", x"cc", x"d4", x"d0", x"d1", x"d0", 
        x"d0", x"d3", x"d2", x"d1", x"d2", x"d1", x"d2", x"d3", x"d5", x"d5", x"d1", x"d3", x"d4", x"d2", x"d2", 
        x"d2", x"d4", x"d7", x"d7", x"d6", x"d4", x"d4", x"d6", x"d1", x"cf", x"d1", x"d3", x"d4", x"d5", x"d4", 
        x"d2", x"d0", x"d4", x"d6", x"d1", x"d2", x"d3", x"d3", x"d5", x"da", x"e0", x"d9", x"c6", x"b3", x"a3", 
        x"94", x"8e", x"91", x"99", x"b7", x"d0", x"ca", x"c9", x"cc", x"c5", x"c7", x"cf", x"cc", x"c5", x"c4", 
        x"c7", x"c8", x"c7", x"ca", x"cf", x"d1", x"d1", x"da", x"e2", x"e3", x"e5", x"ea", x"ed", x"ec", x"f0", 
        x"f4", x"f3", x"f1", x"f3", x"f2", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"ef", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"ee", x"ef", x"f1", x"f0", x"f1", x"f1", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"f0", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f1", x"f0", x"f1", 
        x"e8", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ee", x"ef", x"f1", x"f1", x"f0", x"f0", x"f2", x"f2", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"f0", x"ef", x"ef", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ee", x"ef", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f4", 
        x"ef", x"ee", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f4", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f7", x"f5", x"f4", x"f6", x"f6", x"f5", 
        x"f6", x"f6", x"f3", x"f1", x"f1", x"f2", x"f3", x"f3", x"f1", x"f1", x"f3", x"f3", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f3", x"f3", x"f5", x"f7", x"f7", 
        x"f5", x"f5", x"f6", x"f5", x"f1", x"f1", x"f2", x"f0", x"ed", x"f0", x"eb", x"ed", x"f0", x"f2", x"f1", 
        x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ed", x"f0", 
        x"ef", x"ee", x"f0", x"ee", x"9f", x"53", x"7c", x"bc", x"c1", x"c4", x"b6", x"92", x"a5", x"d0", x"d4", 
        x"dd", x"e2", x"e6", x"ed", x"e2", x"8c", x"4a", x"55", x"b7", x"e4", x"e0", x"d9", x"d8", x"d0", x"a0", 
        x"91", x"8e", x"85", x"7d", x"7e", x"79", x"76", x"7e", x"7b", x"7a", x"73", x"71", x"52", x"51", x"72", 
        x"68", x"63", x"60", x"6e", x"81", x"85", x"7c", x"79", x"85", x"7d", x"53", x"4b", x"60", x"81", x"8b", 
        x"87", x"81", x"7c", x"70", x"68", x"64", x"59", x"54", x"55", x"4c", x"52", x"53", x"50", x"3d", x"43", 
        x"42", x"4d", x"6f", x"70", x"6d", x"75", x"79", x"74", x"74", x"70", x"75", x"74", x"3f", x"4a", x"4c", 
        x"6c", x"6a", x"6a", x"6c", x"6c", x"6c", x"69", x"61", x"5b", x"5b", x"5b", x"5a", x"5a", x"60", x"60", 
        x"42", x"59", x"66", x"68", x"67", x"4a", x"5a", x"68", x"6a", x"66", x"61", x"5e", x"5e", x"65", x"6d", 
        x"6d", x"6b", x"69", x"5a", x"3f", x"59", x"7e", x"a2", x"b3", x"b8", x"bf", x"c9", x"cb", x"cb", x"cf", 
        x"99", x"68", x"7c", x"80", x"7e", x"9c", x"ab", x"b3", x"b7", x"c7", x"cb", x"cd", x"d3", x"d9", x"d8", 
        x"de", x"db", x"d8", x"d7", x"d4", x"d3", x"d5", x"d7", x"d7", x"d7", x"d4", x"d7", x"d7", x"d9", x"d7", 
        x"8d", x"69", x"81", x"92", x"7b", x"61", x"5b", x"49", x"7d", x"6a", x"8e", x"c4", x"c0", x"97", x"86", 
        x"90", x"84", x"75", x"6c", x"6d", x"86", x"84", x"73", x"8c", x"7d", x"81", x"80", x"76", x"7b", x"5c", 
        x"6b", x"74", x"5b", x"64", x"5f", x"6f", x"85", x"83", x"86", x"7d", x"7a", x"73", x"79", x"83", x"6b", 
        x"59", x"71", x"7c", x"54", x"4c", x"42", x"40", x"4d", x"4a", x"3f", x"71", x"7a", x"68", x"74", x"76", 
        x"63", x"82", x"82", x"ac", x"ce", x"d2", x"d8", x"d3", x"d4", x"dc", x"e7", x"e2", x"e0", x"e6", x"ee", 
        x"eb", x"ea", x"ec", x"ed", x"ed", x"e9", x"ea", x"eb", x"ec", x"ec", x"ea", x"eb", x"ea", x"e7", x"e7", 
        x"ea", x"ec", x"eb", x"ec", x"e7", x"e9", x"eb", x"f1", x"ea", x"ec", x"ef", x"f0", x"ec", x"e9", x"e4", 
        x"df", x"d6", x"cb", x"c1", x"b6", x"a9", x"aa", x"a8", x"5e", x"67", x"89", x"95", x"86", x"6c", x"54", 
        x"43", x"38", x"39", x"43", x"5d", x"79", x"95", x"b6", x"c9", x"d6", x"dc", x"da", x"cf", x"bd", x"a7", 
        x"8c", x"73", x"56", x"45", x"3c", x"35", x"3a", x"4e", x"58", x"66", x"70", x"77", x"79", x"7b", x"7b", 
        x"7c", x"76", x"7d", x"c7", x"dd", x"d8", x"d8", x"d7", x"da", x"d5", x"cb", x"d5", x"d0", x"d1", x"d1", 
        x"ce", x"d0", x"d0", x"d0", x"d2", x"d1", x"d3", x"d2", x"d5", x"d4", x"cf", x"d1", x"d3", x"d2", x"d1", 
        x"d2", x"d4", x"d5", x"d6", x"d5", x"d4", x"d4", x"d7", x"d4", x"d2", x"d1", x"d2", x"d4", x"d6", x"d5", 
        x"d2", x"cf", x"d4", x"d8", x"d5", x"d7", x"d8", x"d5", x"ce", x"c5", x"b6", x"a9", x"9b", x"98", x"94", 
        x"93", x"8f", x"92", x"95", x"b4", x"d0", x"b9", x"b2", x"b6", x"b0", x"b3", x"bd", x"ba", x"b6", x"b9", 
        x"c2", x"c4", x"bf", x"be", x"c2", x"c0", x"bd", x"c5", x"cb", x"c5", x"c0", x"c4", x"c2", x"c1", x"c7", 
        x"d1", x"d1", x"d0", x"d6", x"de", x"e0", x"e1", x"e4", x"e8", x"eb", x"ed", x"ee", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", x"f2", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"ef", x"ee", x"ee", x"ed", x"ec", x"ef", x"f2", x"f2", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"f0", x"f1", x"f0", x"f1", 
        x"e8", x"f1", x"f2", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ee", x"ef", x"f2", x"f1", x"ef", x"f0", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f1", x"f1", x"f1", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", 
        x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f1", x"f2", x"f4", 
        x"ef", x"ed", x"f2", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f4", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f4", x"f3", x"f3", x"f8", x"f6", x"f4", x"f5", x"f5", x"f5", 
        x"f6", x"f6", x"f4", x"f2", x"f1", x"f1", x"f2", x"f3", x"f1", x"f1", x"f4", x"f5", x"f4", x"f2", x"f1", 
        x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f4", x"f3", x"f3", x"f3", x"f5", x"f8", x"f6", 
        x"f3", x"f5", x"f5", x"f3", x"ef", x"f0", x"f2", x"f0", x"ed", x"f0", x"ec", x"ed", x"f0", x"f2", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", 
        x"f0", x"ee", x"f0", x"ec", x"ac", x"80", x"79", x"c1", x"d6", x"de", x"da", x"a9", x"b8", x"f3", x"f5", 
        x"f9", x"f9", x"f6", x"f7", x"e7", x"8b", x"4b", x"51", x"9e", x"c0", x"ba", x"ad", x"af", x"a9", x"83", 
        x"7e", x"82", x"81", x"80", x"86", x"8a", x"89", x"8c", x"6f", x"6d", x"76", x"80", x"64", x"4d", x"82", 
        x"8d", x"93", x"99", x"98", x"98", x"93", x"8e", x"85", x"7f", x"70", x"4b", x"3f", x"43", x"55", x"52", 
        x"46", x"44", x"50", x"5b", x"5a", x"57", x"54", x"5a", x"61", x"5e", x"5f", x"67", x"6a", x"50", x"4e", 
        x"54", x"5b", x"76", x"6f", x"69", x"6a", x"69", x"67", x"68", x"66", x"6a", x"6f", x"3e", x"48", x"46", 
        x"66", x"67", x"67", x"69", x"69", x"67", x"66", x"63", x"60", x"5e", x"60", x"62", x"61", x"64", x"65", 
        x"4a", x"5f", x"69", x"68", x"6b", x"46", x"55", x"67", x"64", x"66", x"5e", x"50", x"4f", x"57", x"59", 
        x"54", x"4b", x"45", x"3d", x"30", x"4a", x"6c", x"98", x"ad", x"b8", x"c0", x"c8", x"ce", x"d0", x"d3", 
        x"c6", x"bb", x"c5", x"cf", x"d4", x"dc", x"dd", x"e0", x"de", x"dd", x"dd", x"dc", x"dd", x"d7", x"d3", 
        x"d7", x"d8", x"d6", x"d6", x"d6", x"d4", x"d6", x"d6", x"d6", x"d9", x"d4", x"d8", x"d7", x"d7", x"d6", 
        x"95", x"5d", x"7d", x"93", x"78", x"58", x"56", x"52", x"73", x"61", x"92", x"bd", x"b3", x"7f", x"74", 
        x"76", x"6f", x"79", x"6f", x"82", x"73", x"78", x"84", x"9d", x"a5", x"8d", x"7b", x"71", x"6e", x"6e", 
        x"76", x"7d", x"85", x"64", x"43", x"62", x"97", x"71", x"51", x"5f", x"72", x"74", x"57", x"68", x"69", 
        x"60", x"6d", x"72", x"68", x"54", x"34", x"55", x"70", x"53", x"61", x"82", x"7c", x"7f", x"8c", x"69", 
        x"65", x"83", x"7e", x"7d", x"7a", x"ab", x"c6", x"cc", x"cf", x"e2", x"e2", x"d5", x"d1", x"e2", x"f0", 
        x"ee", x"ec", x"ed", x"e9", x"e7", x"eb", x"ea", x"ea", x"eb", x"e9", x"ea", x"eb", x"eb", x"e6", x"e6", 
        x"e8", x"ec", x"eb", x"eb", x"ed", x"e4", x"e9", x"ec", x"eb", x"eb", x"eb", x"ea", x"e7", x"e8", x"ec", 
        x"e4", x"e5", x"eb", x"e5", x"eb", x"e3", x"e1", x"d5", x"78", x"5a", x"55", x"39", x"21", x"21", x"3f", 
        x"65", x"87", x"ad", x"c1", x"cf", x"d7", x"dd", x"e3", x"df", x"cb", x"ad", x"86", x"5d", x"3e", x"2f", 
        x"36", x"40", x"44", x"4a", x"51", x"5e", x"6d", x"78", x"78", x"7c", x"7f", x"7f", x"7e", x"7f", x"7f", 
        x"7f", x"77", x"7f", x"c8", x"dc", x"d6", x"d9", x"d7", x"d8", x"d8", x"cd", x"d2", x"d1", x"d0", x"d3", 
        x"ce", x"cf", x"d3", x"d5", x"d5", x"d3", x"d3", x"d0", x"d0", x"d2", x"d1", x"d3", x"d5", x"d3", x"d2", 
        x"d2", x"d2", x"d2", x"d5", x"d5", x"d3", x"d2", x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d4", x"d8", 
        x"d8", x"dc", x"e1", x"df", x"c9", x"b5", x"9c", x"8f", x"8c", x"90", x"a5", x"ca", x"c6", x"b0", x"a6", 
        x"a1", x"8f", x"7c", x"73", x"8b", x"9a", x"7a", x"78", x"88", x"84", x"8a", x"9e", x"a1", x"9b", x"9b", 
        x"ad", x"ae", x"a4", x"a7", x"ad", x"ab", x"a5", x"ab", x"b0", x"ae", x"ad", x"bd", x"bc", x"be", x"c0", 
        x"c7", x"ca", x"c5", x"c7", x"c7", x"c1", x"b8", x"b8", x"bd", x"b7", x"b1", x"ba", x"c2", x"c0", x"c2", 
        x"cc", x"d8", x"dc", x"dc", x"e2", x"e9", x"ec", x"ee", x"f5", x"f5", x"f4", x"f6", x"f6", x"f5", x"f3", 
        x"f2", x"f3", x"ef", x"ee", x"eb", x"ea", x"ef", x"f2", x"f3", x"f0", x"ee", x"f1", x"f3", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f0", x"ef", x"f1", x"f2", x"f0", x"f1", x"f4", x"f1", x"ed", x"ef", x"f3", x"f0", 
        x"e6", x"f0", x"f1", x"f1", x"f2", x"f0", x"ef", x"f0", x"f2", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", 
        x"f1", x"ed", x"ef", x"f1", x"f1", x"f1", x"f2", x"f0", x"ef", x"ee", x"ee", x"ee", x"ed", x"ee", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"ef", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f1", x"f0", x"f1", x"f3", x"f3", x"f2", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f3", 
        x"f0", x"ef", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f8", x"f6", x"f4", x"f4", x"f4", x"f5", 
        x"f5", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f4", x"f7", x"f7", x"f5", 
        x"f4", x"f5", x"f4", x"f2", x"f0", x"f0", x"f1", x"f1", x"ef", x"f0", x"ed", x"ef", x"f2", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f0", 
        x"ef", x"f0", x"ef", x"f1", x"b4", x"94", x"6f", x"dc", x"f8", x"f8", x"f4", x"c1", x"c1", x"f6", x"ef", 
        x"e9", x"dd", x"d3", x"c8", x"b7", x"6f", x"44", x"42", x"7e", x"a7", x"b6", x"b7", x"c8", x"c6", x"a0", 
        x"95", x"9f", x"ab", x"94", x"98", x"8e", x"80", x"8e", x"62", x"7f", x"9c", x"9d", x"7e", x"53", x"7c", 
        x"86", x"79", x"6d", x"67", x"61", x"59", x"58", x"57", x"5b", x"53", x"3c", x"39", x"40", x"51", x"4e", 
        x"58", x"6c", x"79", x"83", x"7a", x"70", x"5f", x"5f", x"66", x"64", x"64", x"64", x"63", x"4f", x"53", 
        x"55", x"50", x"6e", x"6d", x"70", x"75", x"72", x"71", x"74", x"64", x"61", x"65", x"42", x"53", x"51", 
        x"71", x"77", x"77", x"77", x"74", x"71", x"6d", x"67", x"61", x"5c", x"5b", x"5d", x"62", x"70", x"6f", 
        x"49", x"64", x"78", x"78", x"75", x"4b", x"45", x"56", x"46", x"39", x"2f", x"1f", x"20", x"31", x"39", 
        x"44", x"52", x"69", x"7f", x"8d", x"a2", x"ba", x"cd", x"d0", x"d4", x"d6", x"d7", x"d7", x"d7", x"d8", 
        x"d9", x"de", x"dd", x"dc", x"db", x"d8", x"d4", x"d5", x"d8", x"d8", x"d8", x"d8", x"da", x"d9", x"d5", 
        x"d8", x"da", x"d7", x"d6", x"d8", x"d3", x"d6", x"d4", x"d6", x"d7", x"d7", x"d8", x"d8", x"d7", x"d7", 
        x"a0", x"5a", x"7a", x"af", x"9a", x"63", x"86", x"74", x"56", x"6d", x"95", x"b3", x"b7", x"9d", x"82", 
        x"78", x"75", x"76", x"77", x"76", x"75", x"87", x"99", x"81", x"65", x"7e", x"7e", x"5c", x"71", x"71", 
        x"4e", x"3f", x"53", x"53", x"49", x"67", x"71", x"67", x"51", x"58", x"64", x"49", x"42", x"5e", x"5c", 
        x"3f", x"62", x"94", x"60", x"56", x"4a", x"32", x"40", x"59", x"53", x"5b", x"65", x"59", x"61", x"6a", 
        x"8f", x"8b", x"8f", x"88", x"82", x"a4", x"b4", x"b0", x"a3", x"aa", x"b6", x"bc", x"af", x"b8", x"cf", 
        x"d5", x"da", x"e0", x"e6", x"ea", x"eb", x"eb", x"ed", x"ee", x"ed", x"ec", x"ea", x"ea", x"e8", x"eb", 
        x"ea", x"ec", x"ea", x"ea", x"e9", x"da", x"e6", x"ea", x"eb", x"eb", x"ed", x"e7", x"e4", x"eb", x"ec", 
        x"e4", x"e3", x"e3", x"df", x"e9", x"ea", x"e3", x"c4", x"62", x"37", x"4e", x"69", x"87", x"a5", x"bf", 
        x"cf", x"d6", x"da", x"d9", x"d0", x"bd", x"a0", x"81", x"63", x"49", x"39", x"39", x"44", x"4b", x"4e", 
        x"54", x"5a", x"65", x"7d", x"92", x"95", x"83", x"7f", x"7f", x"7f", x"80", x"81", x"80", x"80", x"80", 
        x"80", x"77", x"7d", x"c5", x"da", x"d6", x"d8", x"d7", x"d8", x"da", x"ce", x"d1", x"d1", x"d2", x"d4", 
        x"d3", x"d1", x"d0", x"d0", x"d1", x"d3", x"d4", x"d1", x"d0", x"d4", x"d5", x"d4", x"d3", x"d4", x"d5", 
        x"d5", x"d6", x"d6", x"d5", x"d3", x"d2", x"d3", x"d2", x"d2", x"d3", x"d5", x"d5", x"d3", x"d1", x"cc", 
        x"bb", x"a6", x"98", x"95", x"98", x"9f", x"ad", x"b6", x"c1", x"c9", x"d2", x"d6", x"a2", x"7a", x"6b", 
        x"64", x"67", x"74", x"82", x"a6", x"b8", x"92", x"82", x"80", x"73", x"6d", x"72", x"6d", x"60", x"5f", 
        x"6b", x"6c", x"69", x"76", x"81", x"80", x"7b", x"88", x"93", x"8f", x"86", x"92", x"9b", x"98", x"93", 
        x"9a", x"a4", x"a0", x"a1", x"a7", x"aa", x"a7", x"ad", x"be", x"bd", x"b3", x"bc", x"c3", x"bf", x"b9", 
        x"bb", x"bd", x"b4", x"ae", x"b3", x"b4", x"b3", x"ae", x"b6", x"bd", x"bc", x"c2", x"cc", x"d5", x"d4", 
        x"d8", x"e1", x"e4", x"e2", x"e3", x"e5", x"eb", x"ee", x"ee", x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"f0", x"f3", x"f0", x"ef", x"f2", x"f2", x"f0", x"f3", x"f0", 
        x"e6", x"ee", x"f1", x"f0", x"f1", x"f0", x"ef", x"ef", x"f1", x"f3", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"f0", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ec", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"f1", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f3", 
        x"f0", x"ef", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", 
        x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f4", x"f5", x"f6", x"f7", x"f6", x"f4", x"f3", x"f4", x"f5", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f3", x"f1", x"f2", x"f2", x"f2", x"f5", x"f8", x"f7", x"f6", 
        x"f5", x"f4", x"f3", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"ed", x"ef", x"f3", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", 
        x"ee", x"f0", x"ef", x"f5", x"b4", x"73", x"65", x"cd", x"e4", x"d9", x"ce", x"9e", x"93", x"c2", x"bd", 
        x"bd", x"c3", x"cb", x"d2", x"d8", x"92", x"4f", x"40", x"95", x"d6", x"d5", x"d3", x"d9", x"db", x"af", 
        x"9c", x"aa", x"c1", x"a5", x"96", x"64", x"42", x"70", x"4b", x"55", x"66", x"5d", x"51", x"2f", x"4f", 
        x"5b", x"5d", x"5f", x"5f", x"5f", x"5f", x"60", x"63", x"6f", x"71", x"4f", x"42", x"5d", x"83", x"84", 
        x"87", x"8f", x"8a", x"83", x"74", x"66", x"50", x"4e", x"56", x"51", x"54", x"55", x"59", x"49", x"50", 
        x"57", x"46", x"67", x"5e", x"57", x"59", x"5c", x"62", x"6c", x"72", x"77", x"7c", x"58", x"54", x"4c", 
        x"69", x"6a", x"62", x"5e", x"5f", x"65", x"6f", x"71", x"70", x"71", x"73", x"73", x"6c", x"69", x"60", 
        x"39", x"42", x"51", x"49", x"42", x"37", x"42", x"60", x"6d", x"74", x"88", x"93", x"a1", x"b2", x"b7", 
        x"c1", x"c9", x"d2", x"d9", x"da", x"d8", x"da", x"dc", x"d8", x"d8", x"d8", x"d8", x"d8", x"d8", x"da", 
        x"d9", x"db", x"da", x"da", x"da", x"d9", x"d6", x"d7", x"d7", x"d7", x"d6", x"d7", x"da", x"db", x"d6", 
        x"d7", x"d9", x"d7", x"d6", x"d9", x"d6", x"d5", x"d3", x"d6", x"d4", x"d7", x"d8", x"d9", x"d9", x"da", 
        x"98", x"65", x"75", x"a1", x"94", x"6f", x"98", x"70", x"5a", x"73", x"8e", x"a0", x"8d", x"7e", x"7b", 
        x"90", x"87", x"72", x"76", x"5f", x"6e", x"71", x"6e", x"5f", x"4b", x"5f", x"46", x"37", x"6b", x"78", 
        x"56", x"3f", x"54", x"72", x"64", x"4e", x"4b", x"60", x"5e", x"5d", x"4f", x"4d", x"5f", x"4d", x"5f", 
        x"65", x"6e", x"73", x"4d", x"57", x"4a", x"2c", x"4e", x"63", x"45", x"67", x"7e", x"60", x"3c", x"55", 
        x"60", x"66", x"92", x"8b", x"a1", x"b2", x"c8", x"cf", x"b5", x"c5", x"ce", x"d3", x"bb", x"a6", x"bd", 
        x"b8", x"a3", x"9d", x"ae", x"b7", x"c0", x"cf", x"dc", x"df", x"e2", x"e8", x"ed", x"ee", x"eb", x"ec", 
        x"ea", x"ec", x"ed", x"ee", x"ea", x"d7", x"e3", x"ee", x"ee", x"eb", x"ea", x"e7", x"e6", x"e8", x"e8", 
        x"e8", x"e6", x"ec", x"e0", x"d2", x"c9", x"aa", x"92", x"91", x"ad", x"c2", x"d1", x"d9", x"db", x"d9", 
        x"d2", x"c4", x"a5", x"84", x"5e", x"3e", x"31", x"33", x"43", x"50", x"55", x"58", x"5e", x"65", x"75", 
        x"8d", x"a6", x"bc", x"cc", x"d6", x"bb", x"85", x"83", x"87", x"82", x"82", x"82", x"81", x"81", x"81", 
        x"82", x"77", x"7c", x"c3", x"db", x"d5", x"d7", x"d6", x"d8", x"db", x"ce", x"d1", x"d2", x"d3", x"d4", 
        x"d3", x"d2", x"d1", x"d3", x"d4", x"d3", x"d1", x"cf", x"ce", x"d0", x"d3", x"d4", x"d2", x"d3", x"d2", 
        x"d0", x"d3", x"d5", x"d6", x"d5", x"d5", x"d5", x"d7", x"d8", x"d5", x"c8", x"b5", x"9d", x"8d", x"87", 
        x"8f", x"a3", x"b4", x"c5", x"cd", x"d0", x"d5", x"d0", x"cd", x"cb", x"d2", x"e2", x"c1", x"95", x"8b", 
        x"8e", x"84", x"75", x"6e", x"90", x"a9", x"82", x"6e", x"72", x"7e", x"8a", x"94", x"92", x"8c", x"90", 
        x"94", x"90", x"87", x"85", x"84", x"77", x"6a", x"6d", x"6e", x"63", x"55", x"5c", x"66", x"64", x"65", 
        x"76", x"81", x"7c", x"7a", x"8a", x"92", x"89", x"84", x"94", x"98", x"8e", x"90", x"9a", x"9f", x"99", 
        x"97", x"9e", x"a2", x"b8", x"e0", x"d6", x"c8", x"ca", x"d1", x"d0", x"c7", x"c2", x"c6", x"c5", x"ba", 
        x"b5", x"b8", x"b6", x"af", x"ac", x"b2", x"b9", x"b9", x"bc", x"cb", x"d1", x"d1", x"db", x"e6", x"e6", 
        x"e2", x"e7", x"eb", x"eb", x"ea", x"ee", x"f1", x"f2", x"f0", x"f0", x"f1", x"f3", x"f3", x"f5", x"f0", 
        x"e9", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", 
        x"f1", x"ef", x"ee", x"f0", x"f2", x"f1", x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f3", 
        x"f0", x"ef", x"f2", x"f2", x"f2", x"f1", x"f0", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", 
        x"f3", x"f4", x"f5", x"f4", x"f2", x"f2", x"f5", x"f6", x"f6", x"f8", x"f6", x"f4", x"f3", x"f4", x"f5", 
        x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f4", x"f2", x"f2", x"f5", x"f4", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f2", x"f2", x"f6", x"f9", x"f8", x"f6", 
        x"f5", x"f4", x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"ed", x"ef", x"f3", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"ee", x"ee", 
        x"ef", x"f1", x"f1", x"f6", x"b4", x"74", x"5f", x"9b", x"ad", x"bf", x"ca", x"a4", x"9e", x"df", x"e6", 
        x"ea", x"ef", x"f0", x"f1", x"f3", x"a3", x"4f", x"3f", x"9d", x"e3", x"da", x"d6", x"d8", x"d1", x"a4", 
        x"8d", x"89", x"97", x"87", x"60", x"49", x"39", x"4f", x"3d", x"42", x"4e", x"50", x"4e", x"31", x"5b", 
        x"6b", x"6f", x"77", x"84", x"8a", x"8d", x"93", x"94", x"95", x"8c", x"62", x"4b", x"57", x"65", x"59", 
        x"5d", x"6b", x"6b", x"70", x"70", x"73", x"6b", x"66", x"69", x"5c", x"4d", x"45", x"49", x"39", x"30", 
        x"3e", x"40", x"5a", x"60", x"66", x"69", x"6a", x"6a", x"63", x"5d", x"5c", x"65", x"47", x"40", x"4f", 
        x"70", x"7e", x"82", x"82", x"7f", x"78", x"72", x"6a", x"5c", x"4f", x"4d", x"4b", x"46", x"4a", x"5a", 
        x"59", x"6d", x"85", x"8f", x"97", x"aa", x"c0", x"d1", x"d4", x"d9", x"e0", x"de", x"dd", x"da", x"d6", 
        x"d9", x"d7", x"d6", x"d9", x"dc", x"da", x"d9", x"d9", x"d5", x"d5", x"d5", x"d6", x"d8", x"d8", x"db", 
        x"da", x"dc", x"db", x"da", x"db", x"da", x"d8", x"d9", x"d8", x"d6", x"d5", x"d5", x"d8", x"da", x"d7", 
        x"d7", x"d9", x"d6", x"d4", x"d7", x"d6", x"d9", x"d7", x"d6", x"d4", x"d6", x"d8", x"da", x"d8", x"d9", 
        x"8c", x"6f", x"8d", x"87", x"7b", x"6c", x"77", x"60", x"6a", x"82", x"73", x"6f", x"56", x"65", x"7b", 
        x"94", x"91", x"7e", x"7d", x"7e", x"73", x"6f", x"79", x"83", x"5d", x"61", x"58", x"43", x"51", x"5d", 
        x"55", x"44", x"47", x"6b", x"80", x"6d", x"46", x"5a", x"50", x"5e", x"5f", x"69", x"79", x"56", x"5a", 
        x"69", x"6b", x"96", x"92", x"6a", x"48", x"3f", x"3f", x"2e", x"34", x"6b", x"66", x"53", x"4a", x"59", 
        x"57", x"74", x"90", x"78", x"7a", x"95", x"b5", x"b2", x"9a", x"ac", x"db", x"f0", x"d5", x"b5", x"d4", 
        x"e5", x"bf", x"c5", x"d7", x"cc", x"c0", x"b7", x"ba", x"b7", x"b3", x"b8", x"c2", x"cc", x"d4", x"df", 
        x"e3", x"e8", x"e9", x"dc", x"df", x"e4", x"eb", x"ec", x"e9", x"ee", x"ee", x"e8", x"e8", x"e5", x"e5", 
        x"eb", x"e1", x"e3", x"ce", x"ac", x"b5", x"c3", x"ce", x"d8", x"dd", x"d9", x"cf", x"be", x"a7", x"85", 
        x"63", x"4a", x"36", x"34", x"3d", x"4c", x"52", x"57", x"62", x"6d", x"79", x"8d", x"a5", x"ba", x"c9", 
        x"d2", x"d5", x"d6", x"d5", x"d6", x"ba", x"81", x"81", x"85", x"85", x"84", x"83", x"82", x"82", x"83", 
        x"84", x"7b", x"7e", x"c3", x"dd", x"d6", x"d6", x"d4", x"d7", x"da", x"cc", x"d0", x"d2", x"d4", x"d3", 
        x"d1", x"cf", x"cd", x"ce", x"d0", x"d1", x"d2", x"d2", x"d2", x"d3", x"d4", x"d4", x"d3", x"d6", x"d8", 
        x"d6", x"d3", x"d5", x"d7", x"d3", x"c7", x"b9", x"aa", x"9b", x"8c", x"8b", x"96", x"ab", x"bb", x"c5", 
        x"cc", x"d2", x"d1", x"d0", x"cf", x"d1", x"d0", x"d1", x"cf", x"cc", x"d2", x"db", x"aa", x"86", x"73", 
        x"67", x"6b", x"7a", x"7f", x"9b", x"b3", x"92", x"78", x"72", x"78", x"73", x"66", x"68", x"6e", x"6a", 
        x"61", x"62", x"68", x"6b", x"6f", x"73", x"7d", x"87", x"88", x"89", x"88", x"8d", x"8b", x"84", x"81", 
        x"84", x"7f", x"71", x"6d", x"74", x"74", x"68", x"5f", x"6b", x"70", x"66", x"68", x"72", x"77", x"76", 
        x"7a", x"83", x"82", x"98", x"d6", x"c4", x"9d", x"a6", x"b2", x"ad", x"a7", x"ae", x"b3", x"b6", x"b9", 
        x"c4", x"ca", x"c3", x"c6", x"c8", x"d0", x"cd", x"c3", x"c2", x"ca", x"c6", x"be", x"bd", x"bf", x"b8", 
        x"b0", x"b0", x"b7", x"b7", x"b8", x"c3", x"ce", x"d1", x"d0", x"d3", x"d9", x"de", x"e0", x"e3", x"e0", 
        x"e0", x"e6", x"ec", x"ed", x"ec", x"ed", x"ef", x"f0", x"f3", x"f2", x"f3", x"f3", x"f2", x"f1", x"f2", 
        x"f2", x"f2", x"f0", x"f0", x"f1", x"ef", x"ed", x"ee", x"ed", x"eb", x"ed", x"ef", x"ef", x"f0", x"ef", 
        x"f0", x"f1", x"f0", x"ef", x"ed", x"ee", x"f0", x"f1", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f1", x"f3", 
        x"f0", x"ef", x"f2", x"f3", x"f2", x"f0", x"f0", x"f3", x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", 
        x"f4", x"f4", x"f5", x"f4", x"f2", x"f2", x"f5", x"f7", x"f8", x"f8", x"f6", x"f4", x"f3", x"f4", x"f5", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f6", x"f3", x"f3", x"f5", x"f5", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f6", x"f9", x"f8", x"f6", 
        x"f5", x"f3", x"f1", x"f0", x"f1", x"f2", x"f3", x"f1", x"f1", x"f1", x"ed", x"ef", x"f3", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f0", x"f1", 
        x"f1", x"f0", x"f0", x"f4", x"b9", x"92", x"73", x"c0", x"d1", x"e9", x"f2", x"bf", x"aa", x"ec", x"f4", 
        x"f2", x"ee", x"ef", x"ed", x"e6", x"a1", x"59", x"45", x"81", x"ad", x"a6", x"99", x"90", x"8f", x"77", 
        x"70", x"77", x"a2", x"ba", x"86", x"63", x"66", x"74", x"49", x"47", x"69", x"76", x"73", x"4d", x"7b", 
        x"91", x"8f", x"8e", x"86", x"80", x"79", x"6e", x"64", x"62", x"61", x"44", x"38", x"4f", x"68", x"67", 
        x"69", x"74", x"72", x"6e", x"65", x"64", x"5a", x"58", x"60", x"67", x"71", x"6f", x"76", x"5c", x"4a", 
        x"5c", x"44", x"50", x"56", x"54", x"4e", x"55", x"5f", x"63", x"6f", x"77", x"7a", x"56", x"42", x"4e", 
        x"65", x"66", x"59", x"54", x"4d", x"46", x"54", x"65", x"70", x"83", x"96", x"aa", x"b7", x"bc", x"cb", 
        x"d1", x"d7", x"e0", x"df", x"da", x"dd", x"e0", x"da", x"d5", x"da", x"dc", x"db", x"db", x"d7", x"d6", 
        x"d7", x"d6", x"d7", x"d9", x"da", x"d9", x"da", x"dc", x"d8", x"d8", x"d7", x"d7", x"d7", x"d8", x"da", 
        x"d9", x"db", x"da", x"d8", x"d9", x"d9", x"d7", x"d8", x"d8", x"d7", x"d5", x"d5", x"d7", x"da", x"d9", 
        x"d8", x"da", x"d8", x"d4", x"d6", x"d6", x"d7", x"d6", x"d7", x"da", x"d9", x"d6", x"d7", x"da", x"dc", 
        x"8e", x"7e", x"9b", x"83", x"57", x"5b", x"7c", x"79", x"7a", x"76", x"78", x"63", x"5f", x"7d", x"82", 
        x"8f", x"8e", x"84", x"89", x"8f", x"65", x"75", x"71", x"67", x"79", x"79", x"6f", x"69", x"55", x"4f", 
        x"57", x"56", x"3d", x"32", x"3e", x"5f", x"59", x"58", x"5a", x"7f", x"87", x"62", x"63", x"5e", x"5d", 
        x"6d", x"72", x"91", x"70", x"66", x"7b", x"75", x"41", x"3f", x"4a", x"5a", x"79", x"57", x"4e", x"56", 
        x"53", x"5b", x"68", x"5f", x"5e", x"73", x"84", x"73", x"77", x"7c", x"98", x"be", x"b0", x"b6", x"c0", 
        x"d1", x"b9", x"d3", x"ba", x"a3", x"e0", x"f5", x"f1", x"ec", x"e3", x"d6", x"c9", x"c3", x"b8", x"b2", 
        x"ae", x"b6", x"bd", x"c2", x"c8", x"cd", x"d8", x"e6", x"e8", x"ee", x"ea", x"e2", x"ea", x"e8", x"d8", 
        x"db", x"d8", x"d5", x"d3", x"db", x"e2", x"dc", x"ca", x"b9", x"a0", x"80", x"5c", x"3c", x"29", x"2a", 
        x"39", x"4a", x"5c", x"62", x"68", x"70", x"7b", x"91", x"b0", x"ca", x"d9", x"e0", x"de", x"d5", x"cf", 
        x"d0", x"cf", x"d0", x"cf", x"d5", x"be", x"83", x"7e", x"81", x"86", x"85", x"84", x"83", x"83", x"83", 
        x"83", x"7b", x"7e", x"c0", x"dd", x"d7", x"d6", x"d4", x"d6", x"d9", x"ca", x"cd", x"d0", x"d2", x"d0", 
        x"ce", x"cf", x"d2", x"d3", x"d2", x"d1", x"d2", x"d3", x"d3", x"d2", x"d2", x"d6", x"d8", x"d2", x"cd", 
        x"c8", x"bc", x"ab", x"99", x"8b", x"83", x"84", x"98", x"af", x"cb", x"dc", x"e1", x"db", x"d4", x"d0", 
        x"cf", x"d1", x"d0", x"d1", x"d1", x"d2", x"cf", x"cf", x"cd", x"cc", x"d0", x"e0", x"be", x"96", x"87", 
        x"86", x"7e", x"72", x"6b", x"86", x"9d", x"7c", x"68", x"67", x"73", x"75", x"73", x"7b", x"81", x"82", 
        x"7f", x"87", x"8c", x"81", x"74", x"6c", x"76", x"6d", x"5b", x"5d", x"65", x"65", x"5a", x"5b", x"64", 
        x"6d", x"6e", x"71", x"7f", x"8d", x"8d", x"89", x"8c", x"95", x"95", x"89", x"82", x"85", x"85", x"77", 
        x"6f", x"73", x"73", x"94", x"df", x"b1", x"6d", x"70", x"85", x"87", x"81", x"84", x"8f", x"90", x"8b", 
        x"95", x"9b", x"90", x"93", x"a0", x"a6", x"99", x"99", x"a6", x"a9", x"a9", x"b4", x"c2", x"c1", x"c0", 
        x"cb", x"d0", x"cf", x"cc", x"c8", x"c9", x"ca", x"c5", x"bc", x"b8", x"b9", x"ba", x"b1", x"b0", x"b6", 
        x"bf", x"b6", x"c4", x"c7", x"c4", x"ca", x"d2", x"d3", x"d4", x"da", x"e0", x"e1", x"e1", x"e5", x"e9", 
        x"e9", x"e7", x"e9", x"ed", x"ef", x"ef", x"f0", x"f3", x"f3", x"f1", x"f3", x"f3", x"f2", x"f2", x"f2", 
        x"f0", x"ef", x"ef", x"f0", x"f1", x"f0", x"ed", x"ed", x"ee", x"ee", x"ef", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f3", 
        x"f0", x"ef", x"f2", x"f2", x"f2", x"f0", x"f0", x"f3", x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f4", 
        x"f4", x"f5", x"f5", x"f4", x"f2", x"f3", x"f5", x"f7", x"f9", x"f8", x"f6", x"f4", x"f3", x"f4", x"f5", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", 
        x"f1", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f6", x"f9", x"f6", x"f5", 
        x"f4", x"f2", x"f1", x"f0", x"f1", x"f2", x"f3", x"f1", x"f1", x"f1", x"ed", x"ef", x"f3", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", 
        x"f0", x"ee", x"ef", x"f5", x"c2", x"a2", x"79", x"d4", x"da", x"d7", x"e7", x"bc", x"a3", x"d7", x"da", 
        x"d4", x"c1", x"b8", x"b1", x"a6", x"77", x"47", x"33", x"62", x"9d", x"b4", x"c3", x"c9", x"d2", x"b6", 
        x"9f", x"9e", x"c3", x"db", x"a6", x"72", x"6f", x"76", x"5d", x"6a", x"81", x"75", x"75", x"46", x"59", 
        x"5e", x"56", x"58", x"5d", x"63", x"6c", x"71", x"72", x"6f", x"6b", x"52", x"43", x"47", x"5f", x"64", 
        x"66", x"7b", x"8b", x"92", x"8b", x"88", x"7b", x"73", x"6b", x"68", x"5d", x"5c", x"61", x"55", x"4f", 
        x"5a", x"3d", x"6f", x"7a", x"76", x"6f", x"66", x"57", x"49", x"44", x"43", x"46", x"3d", x"46", x"61", 
        x"70", x"83", x"95", x"ab", x"bf", x"c8", x"d9", x"e4", x"e5", x"e9", x"ea", x"e8", x"e4", x"dc", x"dd", 
        x"de", x"de", x"d9", x"d6", x"d8", x"d9", x"dd", x"da", x"d8", x"de", x"db", x"db", x"dc", x"da", x"db", 
        x"da", x"d8", x"d9", x"db", x"da", x"d8", x"d9", x"dd", x"da", x"d9", x"d9", x"d8", x"d9", x"d9", x"db", 
        x"da", x"dc", x"da", x"d8", x"d9", x"da", x"d8", x"d7", x"d8", x"d8", x"d7", x"d7", x"d8", x"db", x"de", 
        x"dd", x"dd", x"d9", x"d6", x"d6", x"d5", x"d7", x"d8", x"d6", x"d5", x"d5", x"d6", x"d8", x"d7", x"d9", 
        x"b6", x"81", x"65", x"5e", x"5a", x"63", x"5f", x"5d", x"5d", x"64", x"64", x"75", x"77", x"6a", x"6b", 
        x"86", x"8d", x"7c", x"7e", x"73", x"79", x"85", x"6e", x"6e", x"7c", x"74", x"7e", x"86", x"7d", x"5a", 
        x"42", x"36", x"5c", x"60", x"55", x"7d", x"7e", x"87", x"74", x"80", x"6e", x"6d", x"60", x"46", x"61", 
        x"5b", x"71", x"6d", x"66", x"78", x"82", x"6e", x"44", x"4f", x"4b", x"52", x"72", x"69", x"58", x"51", 
        x"54", x"5d", x"75", x"7b", x"7d", x"6a", x"8e", x"74", x"6e", x"77", x"6f", x"67", x"74", x"89", x"88", 
        x"93", x"a4", x"b0", x"8a", x"88", x"bf", x"d6", x"e1", x"eb", x"f1", x"f1", x"f0", x"f2", x"f1", x"ef", 
        x"e4", x"dc", x"d2", x"c6", x"b3", x"ab", x"b3", x"c7", x"c8", x"cd", x"ca", x"c9", x"da", x"dc", x"d0", 
        x"d3", x"d6", x"d1", x"c5", x"a9", x"89", x"70", x"5c", x"49", x"3c", x"3b", x"41", x"48", x"51", x"60", 
        x"70", x"7e", x"8e", x"99", x"ad", x"c6", x"d3", x"d6", x"d6", x"d5", x"d2", x"d0", x"d1", x"d3", x"d4", 
        x"d3", x"d2", x"d1", x"d0", x"d6", x"be", x"84", x"83", x"87", x"86", x"85", x"85", x"83", x"83", x"82", 
        x"82", x"78", x"7b", x"bb", x"dc", x"d7", x"d9", x"d7", x"d5", x"d9", x"cc", x"cc", x"ce", x"d2", x"d1", 
        x"d2", x"d2", x"d3", x"d3", x"d3", x"d7", x"da", x"da", x"d7", x"d0", x"c2", x"b2", x"a7", x"9f", x"98", 
        x"93", x"95", x"9c", x"ac", x"bc", x"ca", x"d3", x"d5", x"d4", x"d2", x"cf", x"ce", x"cf", x"d0", x"d0", 
        x"ce", x"d0", x"d1", x"d4", x"d1", x"ce", x"ce", x"d3", x"d1", x"ce", x"d1", x"dd", x"af", x"89", x"78", 
        x"77", x"72", x"72", x"7d", x"a0", x"b4", x"96", x"89", x"84", x"82", x"7f", x"7c", x"7f", x"80", x"79", 
        x"71", x"73", x"75", x"72", x"71", x"75", x"7e", x"79", x"70", x"77", x"80", x"7a", x"73", x"75", x"79", 
        x"76", x"6c", x"6a", x"73", x"75", x"6b", x"65", x"6c", x"72", x"6e", x"66", x"6c", x"77", x"79", x"73", 
        x"77", x"83", x"80", x"97", x"dc", x"bc", x"81", x"76", x"80", x"82", x"78", x"79", x"86", x"84", x"73", 
        x"78", x"84", x"83", x"7c", x"85", x"8f", x"88", x"84", x"8e", x"93", x"87", x"85", x"8f", x"8c", x"83", 
        x"8c", x"9e", x"9d", x"98", x"a1", x"ae", x"b1", x"ac", x"b1", x"b9", x"b9", x"bd", x"c3", x"cc", x"d6", 
        x"e4", x"c6", x"c7", x"ca", x"be", x"be", x"c3", x"bd", x"b6", x"b7", x"bd", x"bd", x"bb", x"bf", x"c3", 
        x"c2", x"c2", x"ca", x"ce", x"cd", x"cd", x"d1", x"d4", x"d5", x"d7", x"dc", x"df", x"e1", x"e6", x"ea", 
        x"ec", x"ed", x"ef", x"f1", x"f4", x"f3", x"f0", x"f1", x"f3", x"f3", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f3", 
        x"f0", x"ef", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f1", x"f2", x"f2", x"f2", x"f4", 
        x"f4", x"f4", x"f4", x"f3", x"f3", x"f4", x"f6", x"f8", x"f9", x"f8", x"f6", x"f4", x"f3", x"f4", x"f5", 
        x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f2", x"f1", x"f3", x"f3", x"f2", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f4", x"f4", x"f3", x"f5", x"f8", x"f6", x"f4", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f1", x"f1", x"f1", x"ed", x"ef", x"f3", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f0", x"ef", x"ef", x"f7", x"cb", x"a5", x"67", x"ad", x"c1", x"af", x"b4", x"96", x"81", x"b1", x"ba", 
        x"bf", x"c0", x"c6", x"d2", x"db", x"a7", x"5b", x"3c", x"85", x"d8", x"d6", x"d5", x"cf", x"c9", x"a2", 
        x"8a", x"8b", x"9f", x"ac", x"a0", x"72", x"55", x"5f", x"4c", x"4f", x"61", x"5c", x"5e", x"39", x"55", 
        x"70", x"6c", x"6f", x"74", x"77", x"7b", x"7b", x"7f", x"7f", x"7b", x"5b", x"49", x"55", x"72", x"7b", 
        x"74", x"78", x"79", x"78", x"72", x"70", x"6d", x"6b", x"6b", x"6c", x"66", x"63", x"60", x"46", x"35", 
        x"42", x"33", x"4c", x"5a", x"5f", x"63", x"72", x"81", x"8f", x"9b", x"a5", x"b0", x"b8", x"c4", x"d4", 
        x"d9", x"e0", x"e1", x"e0", x"de", x"db", x"df", x"e0", x"dd", x"dd", x"dd", x"dc", x"db", x"d9", x"d9", 
        x"d9", x"da", x"d7", x"d9", x"e0", x"dd", x"de", x"db", x"d5", x"db", x"db", x"dc", x"dc", x"da", x"d9", 
        x"d9", x"d6", x"d5", x"d9", x"dc", x"dc", x"db", x"dc", x"d8", x"d8", x"d9", x"d9", x"da", x"da", x"dc", 
        x"db", x"de", x"dc", x"d9", x"da", x"db", x"db", x"da", x"da", x"da", x"d8", x"d8", x"d8", x"da", x"d9", 
        x"d9", x"da", x"d9", x"d9", x"da", x"d7", x"dc", x"e0", x"dd", x"dd", x"d9", x"d9", x"d7", x"d1", x"ce", 
        x"c2", x"7d", x"51", x"4d", x"59", x"6a", x"5e", x"61", x"4c", x"59", x"58", x"74", x"7e", x"67", x"6b", 
        x"7a", x"86", x"6a", x"5f", x"4f", x"73", x"8e", x"7c", x"79", x"84", x"78", x"76", x"86", x"74", x"53", 
        x"42", x"2e", x"58", x"6a", x"60", x"75", x"6c", x"85", x"70", x"71", x"67", x"73", x"59", x"49", x"60", 
        x"36", x"4e", x"69", x"6e", x"70", x"6f", x"53", x"42", x"48", x"43", x"64", x"6b", x"65", x"53", x"45", 
        x"62", x"7b", x"7c", x"7c", x"7e", x"75", x"8d", x"6d", x"70", x"89", x"91", x"72", x"80", x"8a", x"84", 
        x"7e", x"84", x"7e", x"7d", x"8f", x"93", x"94", x"a4", x"b1", x"be", x"c3", x"d0", x"da", x"df", x"e9", 
        x"ef", x"f4", x"f4", x"f1", x"de", x"d5", x"c8", x"ca", x"be", x"bc", x"b5", x"b2", x"c4", x"cc", x"c1", 
        x"b1", x"99", x"77", x"5f", x"46", x"35", x"2f", x"35", x"3f", x"53", x"66", x"72", x"7c", x"89", x"9e", 
        x"b6", x"ca", x"d5", x"d7", x"d9", x"d8", x"d1", x"cc", x"d3", x"d4", x"d1", x"d0", x"d1", x"d3", x"d2", 
        x"d1", x"d1", x"d1", x"d0", x"d5", x"bf", x"88", x"83", x"86", x"85", x"85", x"85", x"84", x"82", x"81", 
        x"81", x"7a", x"7c", x"ba", x"dd", x"d9", x"da", x"d9", x"d5", x"da", x"cd", x"cd", x"cf", x"d3", x"d2", 
        x"d5", x"d7", x"d8", x"d6", x"d0", x"c6", x"bd", x"b2", x"a5", x"9b", x"90", x"8b", x"90", x"9b", x"ad", 
        x"c2", x"d0", x"db", x"dc", x"d7", x"d4", x"d2", x"d0", x"d1", x"d1", x"d0", x"ce", x"ce", x"cf", x"cf", 
        x"cf", x"d1", x"cf", x"cf", x"cd", x"cd", x"ce", x"d3", x"cf", x"cd", x"d1", x"e2", x"bc", x"92", x"7f", 
        x"82", x"77", x"6a", x"70", x"8e", x"9f", x"82", x"77", x"6c", x"66", x"70", x"7c", x"7c", x"7d", x"84", 
        x"87", x"87", x"83", x"83", x"87", x"85", x"83", x"81", x"7e", x"7d", x"7f", x"7b", x"74", x"71", x"70", 
        x"6e", x"6c", x"73", x"7f", x"82", x"77", x"73", x"7f", x"83", x"7c", x"73", x"76", x"7f", x"7c", x"6d", 
        x"6a", x"72", x"71", x"8e", x"db", x"b9", x"79", x"72", x"85", x"8b", x"83", x"87", x"92", x"91", x"84", 
        x"87", x"94", x"96", x"81", x"7d", x"85", x"7f", x"76", x"7c", x"8a", x"81", x"73", x"7b", x"86", x"80", 
        x"7d", x"89", x"8c", x"81", x"80", x"8f", x"94", x"89", x"84", x"8a", x"88", x"86", x"8e", x"9f", x"bc", 
        x"df", x"b2", x"aa", x"ba", x"b6", x"b9", x"c3", x"c4", x"c3", x"ca", x"cf", x"ca", x"c1", x"c0", x"c1", 
        x"bb", x"b3", x"b9", x"b8", x"ad", x"aa", x"b1", x"b3", x"af", x"b0", x"b6", x"b9", x"ba", x"c1", x"c8", 
        x"c8", x"ca", x"cf", x"d0", x"ce", x"d1", x"d9", x"dd", x"df", x"e3", x"e9", x"ed", x"f0", x"f2", x"f2", 
        x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f1", x"f0", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f2", x"f0", x"f1", x"f1", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", 
        x"f0", x"ef", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f4", x"f4", x"f4", x"f4", x"f3", 
        x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f4", 
        x"f5", x"f5", x"f3", x"f3", x"f3", x"f4", x"f7", x"f8", x"f8", x"f8", x"f6", x"f4", x"f3", x"f4", x"f5", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f0", x"ee", x"f2", x"f4", x"f2", x"f4", 
        x"f5", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f4", x"f5", x"f5", x"f4", x"f4", x"f3", x"f2", x"f5", x"f7", x"f5", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", x"f1", x"f1", x"f1", x"ee", x"ef", x"f3", x"f2", x"f1", 
        x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", x"ef", 
        x"f2", x"f0", x"ef", x"f6", x"d0", x"b8", x"65", x"97", x"b9", x"b3", x"b7", x"aa", x"96", x"d6", x"ed", 
        x"f3", x"f7", x"f4", x"f2", x"ef", x"af", x"62", x"43", x"79", x"b7", x"b1", x"b3", x"aa", x"a4", x"87", 
        x"73", x"78", x"89", x"98", x"ad", x"90", x"5a", x"6c", x"5b", x"4f", x"6a", x"67", x"6d", x"4b", x"5d", 
        x"7d", x"7a", x"7d", x"7e", x"80", x"84", x"80", x"7f", x"7d", x"74", x"57", x"4a", x"4b", x"61", x"6b", 
        x"6a", x"71", x"76", x"7e", x"72", x"6d", x"66", x"4d", x"4d", x"51", x"49", x"47", x"4f", x"54", x"53", 
        x"6d", x"86", x"98", x"af", x"c3", x"cd", x"da", x"e1", x"e4", x"e8", x"e4", x"e1", x"e2", x"e0", x"de", 
        x"dd", x"db", x"dc", x"da", x"d8", x"d8", x"dd", x"de", x"dd", x"dc", x"dd", x"dd", x"db", x"db", x"dd", 
        x"dd", x"dd", x"dc", x"dc", x"de", x"dc", x"de", x"de", x"d8", x"dc", x"da", x"da", x"da", x"db", x"da", 
        x"d9", x"d6", x"d5", x"da", x"dd", x"db", x"da", x"da", x"d8", x"d9", x"da", x"da", x"db", x"db", x"dc", 
        x"da", x"dd", x"da", x"d7", x"d8", x"da", x"da", x"d9", x"d9", x"d9", x"d9", x"da", x"dd", x"e0", x"df", 
        x"e0", x"e2", x"df", x"dc", x"d6", x"cb", x"ce", x"c7", x"bd", x"b7", x"a4", x"93", x"8d", x"7a", x"6f", 
        x"a0", x"79", x"60", x"65", x"72", x"9b", x"a0", x"78", x"4e", x"65", x"61", x"65", x"74", x"80", x"9e", 
        x"a4", x"a0", x"90", x"93", x"74", x"72", x"84", x"69", x"52", x"5d", x"5e", x"4c", x"68", x"55", x"38", 
        x"32", x"31", x"52", x"59", x"63", x"65", x"5d", x"67", x"58", x"4b", x"6f", x"80", x"5d", x"75", x"7f", 
        x"4a", x"59", x"68", x"46", x"30", x"4f", x"41", x"49", x"71", x"60", x"57", x"51", x"6e", x"6e", x"60", 
        x"77", x"97", x"6e", x"66", x"6e", x"68", x"64", x"5a", x"6b", x"82", x"88", x"81", x"8c", x"92", x"8f", 
        x"97", x"9e", x"8a", x"98", x"8b", x"74", x"86", x"89", x"85", x"83", x"7f", x"8c", x"91", x"95", x"9e", 
        x"a6", x"ae", x"b2", x"c7", x"d0", x"d4", x"cb", x"db", x"e9", x"e2", x"e8", x"db", x"cc", x"d2", x"c0", 
        x"ae", x"8a", x"41", x"3c", x"4f", x"5c", x"68", x"7a", x"87", x"9a", x"ae", x"bb", x"ca", x"d5", x"d9", 
        x"d8", x"d5", x"d1", x"cf", x"cf", x"d2", x"d1", x"d0", x"d2", x"d2", x"d1", x"d1", x"d1", x"d1", x"d0", 
        x"d0", x"d1", x"d1", x"d2", x"d6", x"bf", x"86", x"84", x"86", x"85", x"86", x"85", x"84", x"81", x"81", 
        x"81", x"7b", x"7d", x"bb", x"de", x"d6", x"d6", x"d5", x"d3", x"d9", x"cf", x"d5", x"d8", x"dd", x"d9", 
        x"ce", x"bc", x"a5", x"94", x"89", x"86", x"8f", x"99", x"a1", x"ad", x"bd", x"ce", x"d8", x"db", x"da", 
        x"d5", x"d1", x"ce", x"ce", x"d0", x"d1", x"cf", x"ce", x"cf", x"d0", x"d1", x"d0", x"ce", x"ce", x"d1", 
        x"cf", x"ce", x"ce", x"cf", x"cf", x"ce", x"cc", x"d0", x"d0", x"cf", x"d2", x"e0", x"b5", x"88", x"74", 
        x"6e", x"6a", x"69", x"70", x"91", x"b1", x"8f", x"75", x"6f", x"6d", x"6f", x"6d", x"69", x"70", x"77", 
        x"76", x"71", x"70", x"78", x"7f", x"7a", x"76", x"7e", x"84", x"7d", x"7b", x"80", x"87", x"80", x"76", 
        x"73", x"78", x"79", x"7a", x"75", x"74", x"7a", x"7e", x"7c", x"76", x"74", x"78", x"80", x"83", x"7f", 
        x"7f", x"85", x"83", x"97", x"d7", x"c0", x"87", x"82", x"8a", x"81", x"76", x"7b", x"83", x"7f", x"77", 
        x"7d", x"84", x"85", x"84", x"8a", x"97", x"93", x"89", x"8e", x"96", x"92", x"86", x"8d", x"94", x"85", 
        x"76", x"7a", x"83", x"7a", x"71", x"7c", x"8a", x"84", x"7b", x"85", x"95", x"8f", x"82", x"8b", x"b3", 
        x"dd", x"a5", x"88", x"96", x"94", x"88", x"84", x"88", x"86", x"8e", x"9b", x"9d", x"95", x"9c", x"ad", 
        x"ac", x"a2", x"a8", x"b3", x"ae", x"a6", x"ae", x"b9", x"b3", x"ad", x"b0", x"b7", x"b5", x"b2", x"b7", 
        x"b3", x"b2", x"b7", x"b4", x"ab", x"a7", x"ac", x"af", x"ac", x"ac", x"b6", x"b1", x"b1", x"b3", x"bb", 
        x"bf", x"be", x"c7", x"d0", x"d3", x"d6", x"de", x"e4", x"eb", x"ed", x"ed", x"f2", x"f5", x"f4", x"f5", 
        x"f5", x"f5", x"f5", x"f4", x"f2", x"f4", x"f5", x"f4", x"f0", x"ef", x"f2", x"f1", x"f1", x"f0", x"f1", 
        x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", x"f3", 
        x"f2", x"f0", x"f1", x"f1", x"f1", x"f3", x"f1", x"f0", x"f1", x"f1", x"f2", x"f2", x"f3", x"f1", x"f3", 
        x"f4", x"f1", x"f1", x"f1", x"f0", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f1", x"ef", x"f0", x"f2", 
        x"f3", x"f2", x"f3", x"f3", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f3", x"f3", x"f3", x"f2", x"f1", 
        x"ef", x"ed", x"f1", x"f0", x"f1", x"f2", x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f4", 
        x"f5", x"f5", x"f3", x"f3", x"f4", x"f6", x"f8", x"f8", x"f8", x"f7", x"f5", x"f4", x"f3", x"f4", x"f4", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"ef", x"ee", x"f1", x"f2", x"f1", x"f2", 
        x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f5", x"f6", x"f5", x"f5", x"f3", x"f2", x"f2", x"f6", x"f7", x"f5", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"ef", x"ed", x"f2", x"f3", x"f2", 
        x"f2", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f0", 
        x"f2", x"f0", x"ef", x"f3", x"d2", x"bf", x"76", x"c8", x"ea", x"eb", x"df", x"c8", x"a1", x"d0", x"dd", 
        x"d1", x"cd", x"c2", x"ba", x"ba", x"8e", x"57", x"3f", x"6a", x"ab", x"ae", x"b4", x"b9", x"bf", x"a4", 
        x"8e", x"95", x"b4", x"d2", x"d7", x"ce", x"94", x"77", x"69", x"60", x"73", x"6a", x"70", x"53", x"5a", 
        x"76", x"74", x"72", x"6f", x"71", x"74", x"6f", x"6e", x"71", x"6a", x"47", x"39", x"33", x"46", x"57", 
        x"4d", x"59", x"61", x"6e", x"75", x"78", x"7c", x"7b", x"8c", x"a2", x"ae", x"b6", x"c8", x"cc", x"d3", 
        x"e5", x"e9", x"e5", x"e6", x"e5", x"e1", x"e0", x"dd", x"dd", x"de", x"da", x"da", x"dd", x"dc", x"dd", 
        x"e1", x"df", x"de", x"de", x"dc", x"db", x"dc", x"da", x"da", x"dc", x"dd", x"dd", x"dc", x"dc", x"de", 
        x"de", x"dc", x"dc", x"dc", x"dc", x"dc", x"db", x"dc", x"da", x"dc", x"dd", x"dd", x"dd", x"dc", x"d9", 
        x"da", x"db", x"da", x"db", x"dd", x"dc", x"dc", x"da", x"d8", x"da", x"db", x"db", x"db", x"d9", x"d8", 
        x"d8", x"d9", x"da", x"d8", x"db", x"e1", x"e3", x"e4", x"e4", x"e1", x"df", x"d9", x"d0", x"ca", x"bd", 
        x"b3", x"a5", x"95", x"81", x"71", x"66", x"5c", x"4f", x"48", x"48", x"3e", x"33", x"36", x"35", x"34", 
        x"af", x"a4", x"8b", x"78", x"6e", x"9b", x"aa", x"6a", x"52", x"74", x"77", x"84", x"8a", x"8c", x"9a", 
        x"b0", x"b3", x"b1", x"c4", x"a1", x"98", x"af", x"92", x"64", x"52", x"52", x"52", x"5a", x"38", x"2c", 
        x"2e", x"43", x"56", x"64", x"47", x"3f", x"63", x"6b", x"64", x"50", x"6b", x"6a", x"62", x"7e", x"7d", 
        x"4d", x"59", x"59", x"55", x"41", x"47", x"3d", x"65", x"73", x"48", x"5b", x"6c", x"63", x"78", x"8a", 
        x"82", x"6c", x"67", x"61", x"73", x"80", x"a1", x"73", x"65", x"6e", x"69", x"72", x"71", x"86", x"8a", 
        x"91", x"97", x"8b", x"8f", x"7e", x"6c", x"86", x"8b", x"9b", x"9b", x"91", x"97", x"97", x"96", x"96", 
        x"95", x"91", x"8a", x"89", x"81", x"92", x"b8", x"a8", x"ad", x"b1", x"c2", x"bc", x"bb", x"dc", x"e2", 
        x"e6", x"ca", x"74", x"77", x"93", x"a4", x"b3", x"c3", x"cb", x"cf", x"d5", x"d6", x"d4", x"d2", x"cf", 
        x"cf", x"d0", x"d1", x"d1", x"d1", x"d0", x"d0", x"d0", x"d1", x"d1", x"d2", x"d2", x"d2", x"d1", x"d0", 
        x"cf", x"d1", x"d2", x"d2", x"d7", x"c1", x"86", x"86", x"88", x"87", x"87", x"86", x"84", x"7f", x"81", 
        x"80", x"7a", x"7c", x"bc", x"dc", x"d6", x"d9", x"d8", x"db", x"dc", x"c9", x"c3", x"b2", x"a2", x"91", 
        x"8b", x"8c", x"94", x"a0", x"aa", x"b6", x"c6", x"cf", x"d4", x"d6", x"d5", x"d2", x"d1", x"d0", x"d1", 
        x"d0", x"cf", x"cf", x"ce", x"cf", x"d2", x"d0", x"ce", x"cd", x"ce", x"cf", x"d0", x"ce", x"cd", x"d0", 
        x"d0", x"cf", x"d0", x"d0", x"d0", x"cf", x"d1", x"d1", x"d0", x"ce", x"cd", x"de", x"be", x"92", x"80", 
        x"7a", x"77", x"76", x"74", x"8d", x"aa", x"88", x"74", x"79", x"82", x"7e", x"76", x"78", x"7f", x"80", 
        x"7b", x"78", x"7b", x"7a", x"75", x"6f", x"72", x"76", x"73", x"6a", x"6c", x"75", x"79", x"73", x"6e", 
        x"76", x"81", x"7e", x"78", x"77", x"7f", x"84", x"7f", x"7b", x"7e", x"81", x"7f", x"7a", x"75", x"74", 
        x"77", x"77", x"72", x"91", x"da", x"be", x"86", x"83", x"89", x"86", x"86", x"91", x"95", x"8c", x"88", 
        x"91", x"93", x"8c", x"82", x"87", x"8c", x"80", x"78", x"80", x"87", x"86", x"7a", x"80", x"8a", x"87", 
        x"83", x"8d", x"96", x"90", x"87", x"8c", x"97", x"93", x"8a", x"8a", x"94", x"8d", x"79", x"7e", x"ae", 
        x"d8", x"a3", x"80", x"87", x"8b", x"86", x"89", x"98", x"99", x"91", x"93", x"93", x"8e", x"8e", x"93", 
        x"8e", x"85", x"7e", x"84", x"86", x"81", x"87", x"94", x"95", x"8f", x"98", x"aa", x"ad", x"a4", x"a6", 
        x"b2", x"b1", x"ad", x"b0", x"b4", x"b1", x"af", x"be", x"d0", x"bb", x"b2", x"ac", x"aa", x"ac", x"b2", 
        x"ad", x"a6", x"ac", x"b3", x"b3", x"b0", x"b2", x"bd", x"b9", x"b6", x"bb", x"c6", x"c9", x"c5", x"cc", 
        x"d1", x"d1", x"d4", x"e0", x"e5", x"e3", x"e6", x"ed", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f1", 
        x"f2", x"f4", x"f4", x"f2", x"f4", x"f1", x"f0", x"f2", x"f1", x"ef", x"f1", x"f1", x"f0", x"ef", x"f1", 
        x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"ef", x"f2", 
        x"f3", x"f0", x"f0", x"f2", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", x"f2", x"f1", x"f0", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f0", x"ed", x"f2", x"f2", x"f1", x"f2", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f4", 
        x"f5", x"f4", x"f4", x"f4", x"f5", x"f7", x"f9", x"fa", x"f9", x"f6", x"f5", x"f5", x"f5", x"f5", x"f5", 
        x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f3", x"f3", x"f3", x"f3", x"f6", x"f8", x"f6", x"f5", x"f3", x"f2", x"f3", x"f7", x"f8", x"f5", x"f3", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"eb", x"f1", x"f3", x"f2", 
        x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f0", 
        x"f1", x"f1", x"f1", x"f5", x"d6", x"bb", x"68", x"9e", x"be", x"b8", x"b6", x"95", x"75", x"b3", x"c7", 
        x"c6", x"ca", x"c9", x"cd", x"d6", x"a8", x"60", x"42", x"76", x"cf", x"d7", x"d4", x"d6", x"da", x"b5", 
        x"97", x"8f", x"9a", x"b5", x"aa", x"a7", x"88", x"65", x"58", x"5f", x"77", x"6a", x"6a", x"46", x"4b", 
        x"6b", x"67", x"65", x"62", x"5c", x"5f", x"60", x"5d", x"66", x"6d", x"58", x"58", x"5d", x"74", x"8e", 
        x"8f", x"a7", x"b3", x"c1", x"d0", x"d1", x"d2", x"d9", x"da", x"e1", x"e3", x"e2", x"e4", x"d3", x"d7", 
        x"e5", x"e1", x"de", x"df", x"df", x"de", x"de", x"de", x"df", x"df", x"dd", x"db", x"dd", x"de", x"de", 
        x"df", x"dd", x"dd", x"de", x"dc", x"dc", x"dd", x"db", x"db", x"dd", x"dd", x"dd", x"dc", x"dc", x"dc", 
        x"dd", x"de", x"dc", x"de", x"dd", x"dc", x"da", x"dd", x"d8", x"da", x"dc", x"dc", x"dc", x"dd", x"dd", 
        x"db", x"da", x"da", x"d8", x"d9", x"db", x"db", x"db", x"da", x"d9", x"d9", x"db", x"de", x"de", x"de", 
        x"dc", x"d9", x"d7", x"cd", x"c7", x"c3", x"b9", x"ac", x"a0", x"8d", x"81", x"74", x"65", x"5f", x"53", 
        x"4c", x"49", x"45", x"3e", x"3a", x"3b", x"3b", x"3a", x"3b", x"40", x"42", x"42", x"44", x"46", x"46", 
        x"b1", x"b4", x"9a", x"8f", x"7d", x"84", x"80", x"6c", x"6c", x"8d", x"77", x"71", x"7b", x"90", x"89", 
        x"8e", x"9f", x"92", x"94", x"90", x"98", x"af", x"a7", x"7a", x"40", x"42", x"6f", x"7e", x"41", x"35", 
        x"45", x"60", x"4e", x"5b", x"51", x"46", x"59", x"6f", x"6c", x"52", x"69", x"76", x"6a", x"80", x"7e", 
        x"7b", x"74", x"59", x"6b", x"54", x"50", x"69", x"7e", x"80", x"62", x"83", x"79", x"50", x"64", x"7b", 
        x"85", x"7e", x"66", x"63", x"83", x"86", x"ac", x"7c", x"5e", x"72", x"67", x"68", x"6e", x"6d", x"7f", 
        x"85", x"87", x"85", x"86", x"84", x"82", x"7b", x"82", x"93", x"9a", x"97", x"9e", x"a5", x"a4", x"a2", 
        x"a7", x"a5", x"9f", x"99", x"7c", x"82", x"ca", x"99", x"83", x"83", x"79", x"75", x"86", x"a0", x"a9", 
        x"aa", x"c1", x"b9", x"c9", x"d8", x"db", x"db", x"dc", x"d8", x"d2", x"cf", x"ce", x"ce", x"d0", x"d2", 
        x"d2", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", x"cf", x"d1", x"d2", x"d2", x"d2", x"d2", x"d1", 
        x"d1", x"d2", x"d3", x"d2", x"d7", x"c2", x"86", x"86", x"88", x"87", x"87", x"87", x"85", x"81", x"81", 
        x"7f", x"79", x"80", x"c4", x"e5", x"da", x"d1", x"c2", x"ac", x"9f", x"86", x"85", x"8a", x"9a", x"a9", 
        x"b8", x"c2", x"cd", x"d4", x"d6", x"d4", x"d4", x"d1", x"cf", x"d1", x"d0", x"d0", x"d2", x"d2", x"d2", 
        x"d0", x"ce", x"ce", x"ce", x"d0", x"d2", x"d0", x"d0", x"d0", x"cf", x"d0", x"d0", x"ce", x"ce", x"d1", 
        x"d1", x"d0", x"d2", x"d3", x"d3", x"d2", x"d2", x"d0", x"cf", x"ce", x"d2", x"de", x"b0", x"86", x"78", 
        x"71", x"66", x"64", x"6e", x"90", x"b2", x"8f", x"76", x"73", x"6c", x"64", x"66", x"6b", x"6b", x"63", 
        x"63", x"6a", x"75", x"76", x"74", x"7c", x"86", x"85", x"7e", x"7f", x"83", x"85", x"7d", x"76", x"74", 
        x"7d", x"7e", x"73", x"69", x"6b", x"6e", x"6b", x"63", x"65", x"6d", x"72", x"6e", x"6b", x"6f", x"7c", 
        x"84", x"81", x"79", x"8f", x"d3", x"c7", x"97", x"96", x"8e", x"80", x"7c", x"82", x"80", x"76", x"79", 
        x"87", x"87", x"7e", x"82", x"8b", x"92", x"8b", x"8a", x"95", x"97", x"8f", x"88", x"93", x"9a", x"8f", 
        x"81", x"82", x"83", x"7b", x"75", x"7b", x"89", x"87", x"7b", x"7c", x"88", x"87", x"85", x"8b", x"b3", 
        x"de", x"b0", x"90", x"98", x"9f", x"99", x"93", x"92", x"89", x"81", x"81", x"88", x"87", x"81", x"81", 
        x"86", x"85", x"86", x"92", x"a0", x"a0", x"96", x"95", x"9b", x"98", x"93", x"90", x"8f", x"88", x"7f", 
        x"84", x"84", x"7e", x"85", x"8d", x"8e", x"8d", x"b0", x"da", x"ab", x"86", x"8f", x"93", x"96", x"99", 
        x"97", x"98", x"9a", x"a1", x"ab", x"b0", x"b0", x"b1", x"ab", x"ae", x"b5", x"b9", x"b6", x"b4", x"b6", 
        x"ba", x"b4", x"b1", x"bb", x"bc", x"b2", x"b5", x"c0", x"c9", x"c7", x"c3", x"cb", x"d1", x"d0", x"d4", 
        x"dd", x"e6", x"e6", x"e7", x"ee", x"f0", x"f0", x"f4", x"f4", x"f3", x"f4", x"f4", x"f2", x"f0", x"f1", 
        x"f1", x"f1", x"f2", x"f3", x"f1", x"f2", x"f3", x"f2", x"f0", x"f1", x"f3", x"f3", x"f3", x"f2", x"f1", 
        x"f0", x"f3", x"f1", x"f1", x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", 
        x"ee", x"f1", x"f1", x"ef", x"f1", x"f2", x"f2", x"f0", x"f1", x"f2", x"f0", x"f2", x"f1", x"f2", x"f3", 
        x"f1", x"eb", x"f0", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", x"f4", x"f4", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f5", x"f4", x"f4", x"f4", x"f5", x"f7", x"f9", x"f9", x"f8", x"f6", x"f5", x"f4", x"f4", x"f5", x"f4", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f1", 
        x"f3", x"f4", x"f4", x"f3", x"f6", x"f8", x"f6", x"f4", x"f2", x"f2", x"f4", x"f7", x"f7", x"f4", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"eb", x"f1", x"f3", x"f2", 
        x"f2", x"f2", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f5", x"d9", x"bb", x"66", x"8a", x"be", x"bf", x"c8", x"9f", x"73", x"c6", x"ea", 
        x"ec", x"eb", x"f0", x"f5", x"f7", x"c1", x"69", x"4c", x"74", x"c1", x"c4", x"ac", x"a8", x"a5", x"87", 
        x"74", x"66", x"81", x"a4", x"a4", x"b0", x"ae", x"8e", x"67", x"56", x"63", x"50", x"52", x"34", x"3c", 
        x"5e", x"5d", x"66", x"72", x"75", x"80", x"93", x"9a", x"a7", x"b8", x"ba", x"c2", x"c9", x"d2", x"d9", 
        x"d9", x"dc", x"e0", x"e0", x"e2", x"de", x"dc", x"e0", x"dd", x"dc", x"df", x"df", x"e0", x"cf", x"d3", 
        x"e3", x"e0", x"df", x"df", x"df", x"dd", x"dc", x"dd", x"de", x"df", x"dd", x"dd", x"df", x"df", x"dd", 
        x"dc", x"db", x"dc", x"de", x"dc", x"dd", x"dc", x"db", x"db", x"dd", x"de", x"de", x"dd", x"dd", x"dd", 
        x"dd", x"db", x"dc", x"e0", x"df", x"de", x"dc", x"df", x"d9", x"dc", x"df", x"dd", x"db", x"db", x"d9", 
        x"db", x"da", x"da", x"dd", x"e1", x"e4", x"e4", x"e5", x"e2", x"dd", x"d8", x"d0", x"c4", x"b7", x"a9", 
        x"99", x"89", x"77", x"65", x"5b", x"56", x"4e", x"47", x"44", x"43", x"46", x"44", x"3e", x"3e", x"40", 
        x"3f", x"41", x"44", x"47", x"49", x"4d", x"50", x"4e", x"4b", x"48", x"47", x"46", x"42", x"3d", x"37", 
        x"97", x"b0", x"a4", x"89", x"91", x"96", x"84", x"69", x"62", x"8c", x"8a", x"89", x"93", x"9a", x"8b", 
        x"96", x"88", x"7c", x"7b", x"78", x"7e", x"61", x"60", x"73", x"78", x"8c", x"7b", x"79", x"72", x"65", 
        x"71", x"6e", x"48", x"55", x"60", x"6d", x"71", x"6c", x"77", x"41", x"51", x"6f", x"75", x"7d", x"83", 
        x"7c", x"4d", x"48", x"70", x"68", x"5d", x"60", x"65", x"7a", x"8c", x"74", x"72", x"6d", x"62", x"4e", 
        x"77", x"71", x"70", x"7b", x"6d", x"73", x"a9", x"98", x"60", x"68", x"73", x"6d", x"74", x"71", x"75", 
        x"8c", x"87", x"85", x"89", x"98", x"90", x"76", x"71", x"7f", x"92", x"92", x"9e", x"aa", x"ad", x"a7", 
        x"a3", x"a0", x"a8", x"af", x"99", x"8f", x"ce", x"a8", x"8c", x"8e", x"89", x"84", x"95", x"8e", x"84", 
        x"70", x"a7", x"d8", x"d8", x"da", x"d6", x"d3", x"d4", x"d3", x"d0", x"d1", x"d1", x"d2", x"d3", x"d3", 
        x"d2", x"d1", x"d0", x"d0", x"d1", x"d2", x"d2", x"d2", x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", 
        x"d3", x"d3", x"d3", x"d2", x"d8", x"c2", x"86", x"86", x"88", x"85", x"85", x"85", x"84", x"82", x"82", 
        x"83", x"7f", x"7b", x"9e", x"a6", x"97", x"90", x"9c", x"ad", x"ba", x"be", x"c9", x"cf", x"d3", x"d4", 
        x"d7", x"d7", x"d7", x"d6", x"d2", x"cf", x"cf", x"cf", x"ce", x"cf", x"ce", x"cf", x"d1", x"d0", x"d1", 
        x"cf", x"cd", x"cd", x"ce", x"d1", x"d3", x"d0", x"d0", x"d0", x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", 
        x"d2", x"d2", x"d2", x"d3", x"d3", x"d2", x"d1", x"ce", x"ce", x"ce", x"d0", x"e2", x"c1", x"96", x"83", 
        x"82", x"7c", x"7a", x"7d", x"8d", x"9e", x"84", x"7a", x"79", x"79", x"7d", x"89", x"8b", x"83", x"81", 
        x"8a", x"8d", x"81", x"74", x"72", x"76", x"72", x"65", x"5e", x"67", x"6d", x"68", x"63", x"64", x"69", 
        x"70", x"76", x"78", x"7d", x"86", x"8b", x"87", x"80", x"81", x"85", x"83", x"7a", x"75", x"7a", x"7d", 
        x"76", x"67", x"64", x"8a", x"d8", x"c3", x"85", x"7e", x"7e", x"82", x"91", x"9d", x"97", x"8e", x"92", 
        x"9b", x"98", x"8e", x"90", x"94", x"90", x"7f", x"7a", x"82", x"81", x"79", x"75", x"83", x"89", x"82", 
        x"7e", x"8b", x"95", x"90", x"8a", x"93", x"9b", x"94", x"8c", x"90", x"9a", x"95", x"86", x"80", x"aa", 
        x"db", x"a5", x"79", x"84", x"8b", x"83", x"7f", x"85", x"8b", x"8b", x"90", x"9f", x"a2", x"99", x"94", 
        x"9b", x"a0", x"98", x"8c", x"8a", x"85", x"7b", x"7f", x"8a", x"87", x"84", x"83", x"85", x"85", x"87", 
        x"95", x"a0", x"a2", x"9e", x"9a", x"99", x"99", x"b3", x"db", x"a6", x"72", x"7a", x"76", x"68", x"66", 
        x"70", x"74", x"6c", x"69", x"74", x"7c", x"7a", x"7a", x"83", x"8c", x"90", x"8d", x"8d", x"91", x"9c", 
        x"a2", x"a6", x"af", x"b6", x"b4", x"b4", x"b6", x"bb", x"c6", x"c3", x"bb", x"b8", x"bd", x"bd", x"b8", 
        x"bf", x"c2", x"b7", x"b1", x"bc", x"c2", x"c0", x"c2", x"c8", x"cf", x"d0", x"d5", x"dd", x"e1", x"df", 
        x"e2", x"eb", x"ee", x"ee", x"ef", x"f0", x"f2", x"f1", x"f1", x"f2", x"f0", x"f0", x"f2", x"f3", x"f3", 
        x"f1", x"f4", x"f0", x"f1", x"f2", x"f1", x"f3", x"f4", x"f1", x"ef", x"f1", x"f3", x"f3", x"f3", x"f3", 
        x"f2", x"f3", x"f3", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ee", x"f0", x"f3", 
        x"f1", x"e9", x"ef", x"f3", x"f2", x"f1", x"f0", x"f0", x"f0", x"f2", x"f4", x"f3", x"f3", x"f3", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f5", x"f4", x"f5", x"f5", x"f6", x"f8", x"f9", x"f9", x"f7", x"f5", x"f4", x"f3", x"f3", x"f4", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", 
        x"f3", x"f4", x"f4", x"f4", x"f7", x"f8", x"f5", x"f3", x"f2", x"f2", x"f5", x"f7", x"f5", x"f2", x"f1", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"eb", x"f1", x"f3", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"ef", 
        x"ee", x"f0", x"f0", x"f1", x"d9", x"c1", x"7a", x"af", x"db", x"df", x"e2", x"c6", x"8a", x"cc", x"f1", 
        x"ec", x"e1", x"d9", x"cd", x"c0", x"99", x"5d", x"4d", x"5c", x"98", x"ac", x"ac", x"b3", x"c1", x"b2", 
        x"91", x"74", x"a5", x"c9", x"ca", x"c7", x"bb", x"8d", x"63", x"57", x"67", x"6d", x"82", x"8e", x"a3", 
        x"b3", x"b9", x"c8", x"d2", x"d6", x"db", x"dd", x"da", x"dd", x"e1", x"e1", x"e3", x"e2", x"df", x"db", 
        x"df", x"dd", x"df", x"de", x"e0", x"df", x"db", x"dd", x"df", x"de", x"df", x"e0", x"e1", x"d1", x"d4", 
        x"e4", x"e2", x"df", x"df", x"df", x"de", x"dd", x"dd", x"df", x"df", x"dc", x"db", x"dd", x"dd", x"db", 
        x"db", x"db", x"de", x"e0", x"dd", x"de", x"de", x"dd", x"dd", x"db", x"dd", x"df", x"de", x"dc", x"da", 
        x"db", x"de", x"de", x"e0", x"df", x"df", x"dd", x"dd", x"d9", x"dc", x"df", x"df", x"df", x"dd", x"d9", 
        x"dc", x"d5", x"ca", x"c4", x"bb", x"aa", x"9b", x"89", x"77", x"69", x"5b", x"51", x"4b", x"49", x"47", 
        x"47", x"49", x"4b", x"49", x"48", x"48", x"47", x"45", x"45", x"49", x"4e", x"50", x"4f", x"51", x"4e", 
        x"4c", x"4a", x"49", x"46", x"42", x"3e", x"35", x"2c", x"27", x"21", x"19", x"14", x"12", x"12", x"10", 
        x"7b", x"8d", x"94", x"66", x"7b", x"9a", x"8d", x"70", x"75", x"91", x"96", x"8d", x"7f", x"8a", x"83", 
        x"85", x"74", x"7d", x"9c", x"82", x"87", x"8d", x"7b", x"6f", x"70", x"97", x"6e", x"7a", x"7e", x"64", 
        x"7f", x"64", x"5e", x"70", x"6a", x"62", x"7a", x"7d", x"84", x"72", x"50", x"3c", x"76", x"76", x"66", 
        x"82", x"66", x"85", x"89", x"6d", x"65", x"6e", x"48", x"48", x"73", x"6f", x"6f", x"5f", x"6c", x"51", 
        x"44", x"48", x"7c", x"8d", x"62", x"69", x"9b", x"6b", x"5b", x"77", x"5c", x"55", x"55", x"77", x"6c", 
        x"6c", x"6d", x"7d", x"75", x"8c", x"84", x"80", x"70", x"68", x"80", x"82", x"98", x"a6", x"ad", x"ac", 
        x"a3", x"98", x"a5", x"a1", x"89", x"93", x"d0", x"b4", x"9a", x"96", x"9a", x"99", x"9a", x"89", x"93", 
        x"81", x"a2", x"da", x"d4", x"d6", x"d7", x"d7", x"d8", x"d5", x"cd", x"cf", x"d2", x"d3", x"d2", x"cf", 
        x"cf", x"d0", x"d0", x"d0", x"d1", x"d2", x"d2", x"d2", x"d1", x"d3", x"d3", x"d2", x"d2", x"d3", x"d3", 
        x"d3", x"d3", x"d2", x"d3", x"d8", x"c3", x"86", x"86", x"88", x"87", x"86", x"84", x"82", x"81", x"7f", 
        x"81", x"7e", x"7a", x"a6", x"c2", x"c8", x"cc", x"d8", x"d8", x"e1", x"d9", x"d4", x"d5", x"d6", x"d5", 
        x"d4", x"d1", x"d0", x"d0", x"cf", x"ce", x"d2", x"d1", x"cf", x"cf", x"cf", x"d0", x"d2", x"cf", x"cf", 
        x"cf", x"cd", x"ce", x"cf", x"d2", x"d4", x"d1", x"d1", x"d2", x"d3", x"d3", x"d2", x"d2", x"d3", x"d4", 
        x"d3", x"d2", x"d2", x"d2", x"d1", x"d0", x"d2", x"d3", x"d2", x"ce", x"ce", x"de", x"b6", x"8c", x"74", 
        x"6c", x"63", x"68", x"79", x"96", x"b5", x"9c", x"87", x"75", x"6e", x"6e", x"70", x"6a", x"60", x"60", 
        x"69", x"6c", x"67", x"69", x"73", x"7b", x"7b", x"7c", x"81", x"8b", x"89", x"81", x"81", x"89", x"8b", 
        x"82", x"76", x"74", x"75", x"73", x"6d", x"64", x"5e", x"64", x"67", x"62", x"5e", x"63", x"70", x"7a", 
        x"79", x"70", x"71", x"89", x"cb", x"cd", x"9d", x"99", x"8c", x"86", x"88", x"83", x"7a", x"73", x"7a", 
        x"80", x"7a", x"72", x"77", x"81", x"83", x"7d", x"86", x"98", x"9c", x"92", x"8c", x"96", x"99", x"90", 
        x"89", x"8f", x"92", x"85", x"79", x"7c", x"80", x"7c", x"78", x"7e", x"84", x"80", x"7d", x"7d", x"a7", 
        x"dd", x"b5", x"90", x"97", x"9b", x"96", x"91", x"94", x"9d", x"99", x"89", x"84", x"88", x"82", x"7c", 
        x"82", x"83", x"7f", x"78", x"83", x"91", x"8d", x"8e", x"9a", x"a2", x"a0", x"98", x"9c", x"a1", x"9b", 
        x"8c", x"89", x"8a", x"86", x"83", x"85", x"87", x"a6", x"d8", x"a2", x"67", x"70", x"79", x"7a", x"7d", 
        x"85", x"87", x"7f", x"7b", x"84", x"88", x"80", x"76", x"78", x"77", x"6e", x"66", x"6a", x"75", x"70", 
        x"67", x"68", x"76", x"7a", x"75", x"7a", x"86", x"8f", x"92", x"8e", x"92", x"94", x"a4", x"d0", x"de", 
        x"c9", x"c6", x"c2", x"c0", x"c2", x"c3", x"c1", x"bd", x"be", x"be", x"bb", x"bb", x"bf", x"b9", x"b3", 
        x"b8", x"c1", x"bd", x"bb", x"c3", x"c9", x"cb", x"cf", x"d9", x"dd", x"db", x"e1", x"e8", x"e7", x"e9", 
        x"ea", x"ed", x"eb", x"f1", x"f1", x"f0", x"f1", x"f3", x"f3", x"f0", x"f1", x"f2", x"f0", x"f3", x"f5", 
        x"f4", x"f2", x"f3", x"f4", x"f2", x"f0", x"f0", x"f2", x"f2", x"f1", x"f2", x"f3", x"f1", x"f3", x"f5", 
        x"f3", x"eb", x"f1", x"f5", x"f4", x"f3", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f1", x"f2", x"f3", 
        x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f5", x"f4", x"f5", x"f5", x"f6", x"f8", x"f9", x"f8", x"f7", x"f5", x"f3", x"f3", x"f3", x"f4", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", 
        x"f4", x"f5", x"f5", x"f5", x"f8", x"f8", x"f5", x"f3", x"f2", x"f2", x"f4", x"f6", x"f4", x"f1", x"f1", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"eb", x"f1", x"f3", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"ee", x"ef", 
        x"ec", x"f0", x"f1", x"f2", x"df", x"bf", x"7d", x"a6", x"d4", x"cb", x"c4", x"b1", x"77", x"9d", x"bd", 
        x"b9", x"ba", x"c0", x"c4", x"ce", x"af", x"62", x"43", x"6b", x"c5", x"d9", x"d5", x"d6", x"d5", x"b3", 
        x"77", x"73", x"a6", x"cc", x"cf", x"ca", x"cc", x"c0", x"be", x"c3", x"ce", x"da", x"de", x"e0", x"e6", 
        x"df", x"e0", x"e3", x"e1", x"e2", x"e3", x"e1", x"de", x"e0", x"df", x"dc", x"de", x"e0", x"e2", x"db", 
        x"dc", x"dc", x"dd", x"dd", x"e0", x"e3", x"dd", x"dd", x"e1", x"df", x"dc", x"dc", x"e0", x"d3", x"d4", 
        x"e4", x"e3", x"de", x"de", x"df", x"df", x"df", x"df", x"df", x"df", x"dc", x"db", x"dd", x"df", x"de", 
        x"df", x"df", x"e1", x"e1", x"dd", x"dd", x"de", x"dd", x"df", x"e0", x"de", x"de", x"de", x"e0", x"e0", 
        x"e1", x"e2", x"e1", x"e1", x"e1", x"e2", x"dd", x"d8", x"d0", x"c9", x"bd", x"b1", x"a4", x"94", x"84", 
        x"77", x"66", x"55", x"4b", x"46", x"45", x"45", x"44", x"46", x"49", x"4c", x"4b", x"4b", x"4c", x"4c", 
        x"4d", x"4f", x"4f", x"50", x"50", x"52", x"53", x"4e", x"4b", x"4c", x"49", x"42", x"3b", x"35", x"2f", 
        x"27", x"1e", x"18", x"14", x"12", x"12", x"11", x"10", x"11", x"0e", x"06", x"04", x"0b", x"1a", x"20", 
        x"ac", x"9b", x"7d", x"67", x"83", x"77", x"63", x"62", x"74", x"78", x"76", x"85", x"7c", x"79", x"79", 
        x"97", x"90", x"91", x"a2", x"82", x"83", x"8e", x"7d", x"6b", x"64", x"75", x"69", x"69", x"60", x"61", 
        x"81", x"6b", x"70", x"70", x"4f", x"41", x"65", x"96", x"87", x"6f", x"58", x"61", x"6b", x"71", x"48", 
        x"6e", x"5e", x"6c", x"63", x"5c", x"64", x"5a", x"30", x"52", x"56", x"57", x"65", x"68", x"76", x"81", 
        x"63", x"4e", x"60", x"58", x"47", x"63", x"87", x"5c", x"54", x"6c", x"5d", x"51", x"59", x"75", x"60", 
        x"59", x"64", x"68", x"6f", x"7c", x"67", x"83", x"7f", x"8c", x"96", x"94", x"a2", x"a8", x"ad", x"af", 
        x"b2", x"a5", x"9c", x"a5", x"8e", x"99", x"cc", x"a6", x"a5", x"a1", x"95", x"96", x"a2", x"a6", x"98", 
        x"7d", x"9f", x"d7", x"d7", x"d6", x"d6", x"d6", x"d8", x"d6", x"ce", x"d0", x"d4", x"d5", x"d2", x"ce", 
        x"cf", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d0", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", 
        x"d2", x"d2", x"d1", x"d3", x"d9", x"c3", x"87", x"86", x"88", x"85", x"85", x"84", x"83", x"84", x"81", 
        x"81", x"78", x"80", x"c8", x"e1", x"db", x"da", x"d8", x"d7", x"e3", x"d6", x"d0", x"d1", x"d1", x"d0", 
        x"d6", x"d5", x"d4", x"d3", x"d1", x"ce", x"cf", x"cf", x"ce", x"cf", x"cf", x"d0", x"d1", x"cf", x"cf", 
        x"cf", x"ce", x"d0", x"d1", x"d3", x"d4", x"d3", x"d4", x"d5", x"d5", x"d3", x"d1", x"d1", x"d2", x"d5", 
        x"d3", x"d2", x"d2", x"d1", x"d0", x"cf", x"d4", x"d2", x"d1", x"ce", x"ce", x"e1", x"c1", x"95", x"7e", 
        x"7f", x"7a", x"77", x"76", x"88", x"a4", x"83", x"71", x"78", x"80", x"85", x"87", x"82", x"81", x"82", 
        x"81", x"80", x"81", x"83", x"84", x"80", x"75", x"70", x"72", x"71", x"69", x"62", x"68", x"6f", x"70", 
        x"69", x"69", x"75", x"7e", x"7f", x"7a", x"75", x"79", x"82", x"82", x"77", x"79", x"83", x"87", x"84", 
        x"7b", x"72", x"6f", x"8a", x"d1", x"c9", x"8b", x"7c", x"76", x"7e", x"89", x"8b", x"85", x"87", x"96", 
        x"99", x"90", x"8b", x"95", x"99", x"93", x"86", x"85", x"87", x"7e", x"74", x"73", x"80", x"80", x"77", 
        x"74", x"7f", x"85", x"80", x"83", x"92", x"9d", x"9b", x"8d", x"87", x"95", x"98", x"8f", x"88", x"ac", 
        x"df", x"b0", x"7d", x"82", x"88", x"86", x"81", x"7f", x"87", x"86", x"86", x"8e", x"9a", x"9c", x"90", 
        x"8c", x"90", x"92", x"8d", x"92", x"9b", x"92", x"8b", x"89", x"89", x"89", x"8a", x"89", x"89", x"8a", 
        x"88", x"89", x"8f", x"98", x"99", x"95", x"94", x"aa", x"d6", x"ae", x"7c", x"83", x"8a", x"87", x"7f", 
        x"76", x"79", x"76", x"71", x"70", x"74", x"74", x"6f", x"71", x"76", x"7a", x"78", x"7b", x"82", x"85", 
        x"7f", x"7d", x"86", x"89", x"7d", x"74", x"70", x"73", x"71", x"66", x"6d", x"70", x"84", x"c5", x"dd", 
        x"c0", x"c2", x"c6", x"c7", x"c6", x"c6", x"c7", x"c6", x"c5", x"c5", x"c7", x"c8", x"c6", x"c2", x"c4", 
        x"c6", x"c5", x"c2", x"c3", x"c9", x"c4", x"bf", x"bb", x"c0", x"bf", x"b6", x"ba", x"c2", x"bb", x"b6", 
        x"bc", x"cb", x"c6", x"c7", x"d0", x"d5", x"d6", x"db", x"e4", x"e8", x"e6", x"e6", x"ea", x"ed", x"ed", 
        x"ed", x"ee", x"ef", x"f1", x"f1", x"f1", x"f3", x"f4", x"f5", x"f5", x"f3", x"f1", x"f0", x"f2", x"f3", 
        x"f0", x"eb", x"f2", x"f4", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f4", x"f3", x"f1", x"f2", x"f3", 
        x"f3", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f5", x"f4", x"f5", x"f5", x"f7", x"f8", x"fa", x"f8", x"f6", x"f5", x"f3", x"f3", x"f3", x"f4", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f5", x"f6", x"f6", x"f8", x"f8", x"f4", x"f2", x"f2", x"f2", x"f3", x"f4", x"f3", x"f1", x"f1", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"eb", x"f1", x"f3", x"f1", 
        x"f1", x"f1", x"f0", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f2", 
        x"ef", x"f3", x"f5", x"f5", x"e4", x"c3", x"78", x"7b", x"b5", x"b8", x"b9", x"b6", x"75", x"9c", x"dc", 
        x"e8", x"e9", x"ef", x"f1", x"f2", x"c8", x"6d", x"40", x"6c", x"c2", x"d8", x"d9", x"d9", x"db", x"cf", 
        x"bd", x"c8", x"d4", x"df", x"e0", x"db", x"e1", x"e3", x"e4", x"e1", x"e1", x"e3", x"e3", x"e3", x"e2", 
        x"de", x"df", x"e2", x"e2", x"e0", x"df", x"e1", x"e1", x"e0", x"df", x"e0", x"e3", x"df", x"e2", x"dd", 
        x"dc", x"e0", x"e0", x"df", x"df", x"e2", x"dd", x"dd", x"dd", x"dc", x"de", x"dd", x"e2", x"d7", x"d3", 
        x"e2", x"e4", x"de", x"de", x"e0", x"e0", x"df", x"df", x"df", x"e0", x"de", x"dd", x"de", x"df", x"de", 
        x"de", x"df", x"e0", x"e0", x"df", x"de", x"e0", x"df", x"de", x"e1", x"de", x"de", x"dd", x"d9", x"d3", 
        x"cc", x"c3", x"bb", x"b1", x"a2", x"96", x"86", x"77", x"6a", x"5f", x"50", x"4a", x"4c", x"4d", x"4b", 
        x"4b", x"4c", x"4e", x"50", x"51", x"53", x"55", x"55", x"55", x"58", x"59", x"57", x"54", x"54", x"53", 
        x"4f", x"4c", x"45", x"42", x"3c", x"34", x"2d", x"22", x"1e", x"1a", x"16", x"15", x"16", x"14", x"14", 
        x"13", x"14", x"18", x"1c", x"1f", x"21", x"20", x"22", x"22", x"1e", x"0e", x"04", x"0c", x"23", x"27", 
        x"b5", x"ae", x"78", x"68", x"82", x"72", x"78", x"80", x"7c", x"7e", x"77", x"78", x"79", x"75", x"70", 
        x"8b", x"8a", x"6c", x"7c", x"77", x"74", x"80", x"7d", x"83", x"6b", x"69", x"68", x"64", x"55", x"59", 
        x"76", x"71", x"70", x"7a", x"58", x"58", x"5b", x"64", x"7b", x"70", x"74", x"6b", x"7f", x"6a", x"3f", 
        x"6d", x"61", x"5e", x"50", x"68", x"5e", x"4e", x"48", x"60", x"59", x"5e", x"3e", x"45", x"70", x"70", 
        x"47", x"6c", x"73", x"54", x"60", x"71", x"75", x"62", x"5a", x"68", x"55", x"36", x"4f", x"68", x"67", 
        x"70", x"6f", x"78", x"8a", x"7c", x"66", x"8b", x"8f", x"88", x"87", x"84", x"92", x"a1", x"b1", x"b6", 
        x"bd", x"b2", x"a2", x"a3", x"9c", x"a7", x"d6", x"aa", x"b4", x"ac", x"8e", x"88", x"9b", x"a8", x"94", 
        x"85", x"a6", x"da", x"d4", x"d2", x"d4", x"d5", x"d7", x"d7", x"d1", x"d3", x"d4", x"d3", x"d2", x"d1", 
        x"d2", x"d3", x"d3", x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d3", x"d3", x"d2", x"d1", 
        x"d0", x"d1", x"d1", x"d2", x"d9", x"c4", x"87", x"86", x"87", x"83", x"85", x"87", x"87", x"88", x"82", 
        x"82", x"76", x"7b", x"ca", x"e3", x"dc", x"de", x"d8", x"d7", x"e3", x"d4", x"d2", x"d2", x"d3", x"d2", 
        x"d3", x"d3", x"d2", x"d0", x"d0", x"d1", x"d1", x"cf", x"ce", x"ce", x"cc", x"cd", x"ce", x"ce", x"ce", 
        x"cf", x"d0", x"d3", x"d2", x"d4", x"d5", x"d3", x"d4", x"d6", x"d6", x"d3", x"d1", x"d0", x"d2", x"d5", 
        x"d4", x"d2", x"d3", x"d2", x"d2", x"d1", x"d4", x"d3", x"d0", x"cc", x"cf", x"dd", x"b3", x"86", x"6d", 
        x"69", x"69", x"6f", x"75", x"93", x"b9", x"9a", x"85", x"80", x"7e", x"74", x"6d", x"70", x"72", x"6c", 
        x"61", x"5e", x"66", x"6c", x"6b", x"6c", x"6f", x"7a", x"84", x"85", x"81", x"80", x"8a", x"88", x"85", 
        x"82", x"84", x"89", x"87", x"78", x"70", x"6f", x"72", x"73", x"6b", x"61", x"63", x"6b", x"6d", x"67", 
        x"65", x"6b", x"6f", x"84", x"c8", x"d0", x"9d", x"93", x"93", x"9c", x"9e", x"91", x"85", x"81", x"85", 
        x"7c", x"71", x"74", x"7b", x"79", x"72", x"74", x"83", x"8d", x"87", x"82", x"88", x"9a", x"9a", x"8e", 
        x"8c", x"99", x"a1", x"92", x"82", x"7f", x"80", x"7f", x"76", x"76", x"81", x"80", x"79", x"74", x"96", 
        x"d7", x"ba", x"86", x"93", x"a1", x"a2", x"99", x"8f", x"96", x"9b", x"98", x"90", x"90", x"91", x"86", 
        x"7d", x"80", x"89", x"85", x"80", x"83", x"84", x"83", x"88", x"97", x"a2", x"9e", x"93", x"91", x"96", 
        x"96", x"94", x"98", x"9c", x"96", x"89", x"82", x"9d", x"d7", x"b3", x"7c", x"7a", x"79", x"79", x"79", 
        x"78", x"7a", x"83", x"87", x"83", x"83", x"88", x"88", x"83", x"81", x"82", x"81", x"79", x"6e", x"75", 
        x"7c", x"78", x"74", x"78", x"79", x"74", x"69", x"6b", x"78", x"7d", x"7d", x"75", x"80", x"c1", x"d9", 
        x"c1", x"c1", x"bc", x"b6", x"b6", x"b9", x"ba", x"b8", x"b7", x"ba", x"c2", x"c6", x"c6", x"c6", x"c6", 
        x"c6", x"c7", x"ca", x"cd", x"d0", x"ca", x"c8", x"c6", x"ce", x"d1", x"c8", x"c9", x"d0", x"cb", x"bb", 
        x"bf", x"d1", x"b7", x"ad", x"b1", x"b2", x"af", x"b0", x"b5", x"b8", x"b2", x"b2", x"c0", x"c2", x"c0", 
        x"c6", x"d0", x"d3", x"d4", x"e2", x"e5", x"e2", x"df", x"e4", x"eb", x"e9", x"ea", x"ed", x"ef", x"ee", 
        x"ed", x"ea", x"f3", x"f4", x"f4", x"f4", x"f5", x"f5", x"f5", x"f6", x"f7", x"f5", x"f2", x"f3", x"f5", 
        x"f5", x"f3", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f3", x"f3", x"f3", x"f3", x"f4", 
        x"f5", x"f4", x"f5", x"f5", x"f7", x"f9", x"fa", x"f7", x"f5", x"f5", x"f4", x"f3", x"f3", x"f4", x"f3", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f5", x"f6", x"f6", x"f8", x"f7", x"f4", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"eb", x"f1", x"f2", x"f1", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f3", 
        x"ef", x"f3", x"f5", x"f4", x"e6", x"c4", x"84", x"8c", x"da", x"ec", x"e7", x"dc", x"83", x"a3", x"e8", 
        x"f3", x"ee", x"f0", x"f0", x"ec", x"db", x"b7", x"b4", x"cc", x"e3", x"de", x"e0", x"e3", x"e5", x"e3", 
        x"e7", x"e5", x"e1", x"e2", x"df", x"df", x"e0", x"e3", x"e0", x"de", x"dd", x"e0", x"e3", x"e4", x"e1", 
        x"df", x"e1", x"e1", x"e1", x"e0", x"df", x"e1", x"e1", x"de", x"e1", x"e4", x"e4", x"de", x"df", x"dc", 
        x"dd", x"df", x"df", x"e0", x"de", x"e0", x"de", x"df", x"de", x"de", x"e1", x"de", x"e1", x"d7", x"cf", 
        x"de", x"e2", x"e0", x"e0", x"e0", x"e0", x"df", x"df", x"e0", x"e1", x"e0", x"e0", x"e3", x"e3", x"e2", 
        x"e0", x"e0", x"dc", x"dc", x"da", x"d3", x"d0", x"cb", x"c0", x"b9", x"ae", x"a1", x"94", x"83", x"71", 
        x"62", x"57", x"50", x"47", x"3e", x"42", x"48", x"4f", x"54", x"57", x"57", x"59", x"5c", x"5d", x"5a", 
        x"5a", x"5b", x"5a", x"58", x"58", x"5a", x"59", x"54", x"4b", x"45", x"40", x"3a", x"32", x"2c", x"23", 
        x"1d", x"18", x"11", x"11", x"10", x"0e", x"0f", x"11", x"17", x"1d", x"1e", x"23", x"25", x"21", x"28", 
        x"26", x"27", x"29", x"28", x"28", x"2c", x"27", x"2e", x"39", x"3b", x"1e", x"06", x"1d", x"4a", x"4d", 
        x"72", x"83", x"79", x"73", x"8b", x"91", x"82", x"76", x"62", x"60", x"7a", x"7f", x"96", x"83", x"82", 
        x"79", x"71", x"60", x"59", x"71", x"77", x"76", x"58", x"62", x"63", x"53", x"55", x"62", x"62", x"5e", 
        x"60", x"53", x"42", x"52", x"59", x"77", x"7e", x"5c", x"4f", x"5f", x"85", x"66", x"4c", x"33", x"32", 
        x"4d", x"62", x"69", x"70", x"62", x"61", x"5b", x"56", x"65", x"5e", x"71", x"68", x"69", x"77", x"66", 
        x"4c", x"7a", x"65", x"53", x"4c", x"59", x"74", x"66", x"73", x"89", x"73", x"51", x"5d", x"6e", x"6a", 
        x"6f", x"6d", x"76", x"99", x"9a", x"62", x"7d", x"7f", x"74", x"85", x"83", x"4a", x"36", x"67", x"67", 
        x"72", x"94", x"91", x"8b", x"8f", x"9f", x"d4", x"a4", x"97", x"9b", x"8f", x"87", x"a4", x"b0", x"96", 
        x"7c", x"a0", x"d8", x"d8", x"d5", x"d7", x"d7", x"d8", x"d7", x"d0", x"d2", x"d1", x"d1", x"d2", x"d3", 
        x"d4", x"d4", x"d3", x"d3", x"d2", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", x"d1", 
        x"cf", x"cf", x"d0", x"d2", x"d6", x"c3", x"8a", x"83", x"86", x"86", x"89", x"89", x"87", x"86", x"83", 
        x"83", x"7a", x"7d", x"c5", x"e0", x"d9", x"d9", x"d7", x"d6", x"e1", x"d2", x"cf", x"cf", x"cf", x"cf", 
        x"d0", x"d2", x"d2", x"d1", x"d2", x"d3", x"d1", x"d0", x"d2", x"d1", x"cf", x"cf", x"d0", x"d0", x"d0", 
        x"d0", x"d1", x"d3", x"d4", x"d5", x"d6", x"d4", x"d3", x"d4", x"d4", x"d3", x"d2", x"d2", x"d3", x"d3", 
        x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d1", x"d3", x"d3", x"ce", x"cf", x"e3", x"c3", x"94", x"7f", 
        x"82", x"7f", x"7a", x"76", x"86", x"a4", x"87", x"77", x"79", x"77", x"78", x"80", x"87", x"86", x"7e", 
        x"7e", x"81", x"84", x"80", x"78", x"71", x"76", x"78", x"74", x"6e", x"70", x"77", x"79", x"6e", x"66", 
        x"67", x"74", x"7c", x"78", x"72", x"76", x"81", x"86", x"80", x"78", x"79", x"80", x"85", x"80", x"78", 
        x"77", x"7b", x"77", x"89", x"ce", x"cb", x"8c", x"78", x"7b", x"86", x"86", x"7e", x"82", x"8d", x"98", 
        x"90", x"87", x"90", x"96", x"90", x"86", x"88", x"93", x"92", x"83", x"79", x"7d", x"87", x"82", x"78", 
        x"77", x"80", x"82", x"78", x"76", x"83", x"8f", x"8f", x"88", x"88", x"94", x"94", x"8d", x"84", x"a4", 
        x"dd", x"c0", x"91", x"87", x"86", x"87", x"86", x"84", x"8b", x"8e", x"89", x"81", x"89", x"92", x"93", 
        x"8f", x"95", x"99", x"94", x"8d", x"8e", x"95", x"98", x"90", x"8a", x"8c", x"8d", x"84", x"7d", x"82", 
        x"90", x"92", x"8d", x"8b", x"90", x"94", x"90", x"9e", x"d3", x"b7", x"85", x"85", x"80", x"82", x"8a", 
        x"88", x"80", x"81", x"86", x"81", x"77", x"73", x"7f", x"82", x"7b", x"72", x"75", x"7d", x"7d", x"7a", 
        x"86", x"8c", x"89", x"85", x"82", x"81", x"7f", x"7b", x"79", x"77", x"76", x"70", x"7e", x"bf", x"d6", 
        x"b6", x"b5", x"b7", x"b9", x"b9", x"bb", x"bf", x"b9", x"b6", x"b6", x"bb", x"be", x"c0", x"bc", x"b7", 
        x"b6", x"b8", x"b6", x"b7", x"b9", x"b8", x"b9", x"b9", x"bf", x"c4", x"bf", x"bc", x"c1", x"c7", x"bf", 
        x"c2", x"d5", x"a8", x"96", x"99", x"96", x"97", x"9d", x"a2", x"a1", x"9f", x"a2", x"a7", x"a7", x"a6", 
        x"aa", x"af", x"af", x"ac", x"b7", x"bc", x"b7", x"b2", x"b8", x"bf", x"bc", x"b9", x"c3", x"c9", x"c8", 
        x"cd", x"d4", x"d8", x"d7", x"d8", x"de", x"e2", x"e0", x"e1", x"e7", x"eb", x"ea", x"eb", x"f0", x"f5", 
        x"f6", x"f5", x"f5", x"f5", x"f5", x"f5", x"f5", x"f3", x"f2", x"f4", x"f4", x"f2", x"f3", x"f2", x"f3", 
        x"f3", x"f5", x"f3", x"f5", x"f6", x"f7", x"f7", x"f4", x"f4", x"f3", x"f2", x"f2", x"f3", x"f4", x"f4", 
        x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f3", 
        x"f2", x"f3", x"f2", x"f3", x"f3", x"f2", x"f3", x"f4", x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f5", 
        x"f3", x"f4", x"f6", x"f5", x"f7", x"f7", x"f4", x"f4", x"f3", x"f2", x"f1", x"f0", x"f1", x"f0", x"f1", 
        x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"ef", x"f0", x"f1", x"f0", x"ec", x"f2", x"f3", x"f0", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f0", x"f0", 
        x"ef", x"f2", x"f4", x"f4", x"e9", x"bf", x"8e", x"9b", x"d8", x"e9", x"e7", x"d7", x"ac", x"c7", x"e4", 
        x"e8", x"e4", x"e0", x"df", x"df", x"e5", x"e9", x"e8", x"e5", x"e5", x"e3", x"e2", x"e4", x"e3", x"e2", 
        x"e2", x"e3", x"e3", x"e2", x"e4", x"e3", x"e0", x"e1", x"e1", x"e2", x"e3", x"e1", x"e1", x"e4", x"e2", 
        x"df", x"e0", x"e1", x"e0", x"e1", x"e2", x"e3", x"e1", x"df", x"e1", x"e1", x"e0", x"df", x"de", x"dd", 
        x"df", x"e1", x"e4", x"e2", x"e0", x"e0", x"de", x"df", x"e0", x"e0", x"e1", x"dd", x"e0", x"d8", x"cf", 
        x"df", x"e4", x"e2", x"e4", x"e6", x"e7", x"e5", x"e5", x"e2", x"de", x"da", x"d1", x"cb", x"c6", x"bc", 
        x"b4", x"a8", x"98", x"8c", x"81", x"74", x"6a", x"62", x"59", x"55", x"4e", x"48", x"48", x"4d", x"52", 
        x"54", x"59", x"5e", x"63", x"62", x"63", x"60", x"60", x"5e", x"60", x"5f", x"5d", x"56", x"4d", x"48", 
        x"44", x"3f", x"3a", x"35", x"30", x"25", x"1c", x"16", x"0f", x"0e", x"14", x"17", x"17", x"15", x"16", 
        x"1b", x"1a", x"18", x"18", x"18", x"17", x"1d", x"21", x"24", x"25", x"23", x"2e", x"34", x"30", x"32", 
        x"36", x"40", x"49", x"4f", x"5a", x"5d", x"5e", x"63", x"69", x"64", x"30", x"08", x"23", x"5d", x"60", 
        x"74", x"72", x"6d", x"7b", x"79", x"7c", x"77", x"71", x"7b", x"86", x"6d", x"76", x"7c", x"63", x"76", 
        x"86", x"77", x"7a", x"79", x"7b", x"71", x"70", x"5c", x"58", x"5b", x"55", x"61", x"70", x"5b", x"49", 
        x"50", x"4c", x"4d", x"3b", x"25", x"55", x"7f", x"67", x"62", x"6c", x"6d", x"5d", x"4d", x"57", x"45", 
        x"4b", x"60", x"62", x"5c", x"58", x"73", x"55", x"61", x"7a", x"5e", x"6b", x"78", x"70", x"6f", x"6d", 
        x"5e", x"5b", x"55", x"77", x"7f", x"5e", x"58", x"76", x"82", x"7b", x"5d", x"71", x"6c", x"78", x"80", 
        x"7d", x"7f", x"7d", x"a3", x"ac", x"79", x"7d", x"6b", x"72", x"87", x"93", x"6f", x"4e", x"71", x"5a", 
        x"6c", x"97", x"81", x"86", x"82", x"84", x"d8", x"b0", x"79", x"6b", x"52", x"53", x"6b", x"79", x"76", 
        x"74", x"9f", x"d9", x"d6", x"d5", x"d7", x"d5", x"d7", x"d7", x"d2", x"d1", x"d2", x"d2", x"d4", x"d4", 
        x"d4", x"d4", x"d2", x"d2", x"d2", x"d3", x"d2", x"d2", x"d1", x"d4", x"d3", x"d1", x"d1", x"d2", x"d1", 
        x"d0", x"ce", x"d1", x"d2", x"d4", x"c3", x"8f", x"83", x"87", x"87", x"87", x"84", x"81", x"84", x"85", 
        x"83", x"7c", x"81", x"c5", x"e2", x"dc", x"db", x"d9", x"d7", x"e1", x"d5", x"cd", x"d0", x"d0", x"d0", 
        x"d2", x"d2", x"d3", x"d3", x"d2", x"d0", x"cf", x"cf", x"cf", x"cf", x"d0", x"d0", x"d1", x"d1", x"d2", 
        x"d2", x"d0", x"d1", x"d4", x"d6", x"d7", x"d6", x"d4", x"d3", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", 
        x"d3", x"d4", x"d4", x"d4", x"d4", x"d3", x"d4", x"d4", x"d2", x"ce", x"cf", x"e0", x"be", x"8c", x"79", 
        x"76", x"74", x"75", x"7d", x"92", x"ad", x"95", x"83", x"77", x"6e", x"74", x"77", x"74", x"6d", x"68", 
        x"6f", x"74", x"72", x"6d", x"70", x"79", x"7b", x"77", x"74", x"79", x"80", x"84", x"7f", x"79", x"76", 
        x"7a", x"84", x"83", x"77", x"70", x"74", x"79", x"74", x"6a", x"67", x"70", x"78", x"76", x"6e", x"6d", 
        x"74", x"79", x"72", x"82", x"c8", x"cd", x"93", x"81", x"8d", x"95", x"90", x"84", x"83", x"86", x"88", 
        x"80", x"77", x"84", x"8d", x"87", x"7b", x"7b", x"86", x"88", x"81", x"80", x"8a", x"96", x"91", x"87", 
        x"86", x"90", x"94", x"8b", x"81", x"88", x"91", x"8e", x"80", x"79", x"88", x"8d", x"86", x"7c", x"9b", 
        x"d9", x"ba", x"84", x"84", x"91", x"97", x"96", x"96", x"96", x"99", x"98", x"91", x"94", x"9a", x"9a", 
        x"8d", x"81", x"7f", x"83", x"83", x"7f", x"85", x"8c", x"8e", x"86", x"87", x"92", x"98", x"93", x"91", 
        x"97", x"9a", x"96", x"91", x"96", x"9c", x"96", x"a3", x"d3", x"b4", x"7b", x"7a", x"76", x"74", x"7a", 
        x"7d", x"79", x"76", x"77", x"7c", x"7f", x"7f", x"83", x"86", x"82", x"79", x"7a", x"83", x"87", x"85", 
        x"83", x"80", x"81", x"7c", x"73", x"70", x"78", x"7c", x"70", x"67", x"6a", x"6d", x"7e", x"bd", x"d8", 
        x"ba", x"b9", x"b6", x"b9", x"c0", x"c1", x"bb", x"b6", x"b6", x"b8", x"bb", x"bb", x"bb", x"b2", x"b5", 
        x"b7", x"ba", x"b8", x"b9", x"b7", x"b6", x"b9", x"be", x"c0", x"bc", x"b6", x"b5", x"b5", x"b8", x"b7", 
        x"ba", x"d1", x"9a", x"7d", x"7a", x"75", x"7c", x"89", x"88", x"81", x"86", x"8e", x"8b", x"8b", x"92", 
        x"95", x"91", x"91", x"98", x"9e", x"9f", x"9f", x"a3", x"a8", x"ac", x"ac", x"ac", x"b6", x"b6", x"b2", 
        x"c4", x"cd", x"bb", x"b1", x"af", x"b6", x"bc", x"b8", x"b5", x"be", x"c2", x"c0", x"c5", x"cf", x"d3", 
        x"d1", x"d4", x"dc", x"df", x"df", x"e2", x"e5", x"e7", x"e8", x"eb", x"ef", x"f1", x"f3", x"f4", x"f6", 
        x"f4", x"f4", x"f2", x"f8", x"f8", x"f8", x"f7", x"f3", x"f4", x"f4", x"f3", x"f3", x"f3", x"f5", x"f4", 
        x"f2", x"f2", x"f4", x"f4", x"f3", x"f3", x"f3", x"f1", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f3", 
        x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f1", x"f2", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f4", x"f7", x"f4", x"f7", x"f8", x"f7", x"f4", x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", 
        x"f1", x"f1", x"f2", x"f2", x"ef", x"ef", x"f0", x"ee", x"ef", x"f1", x"ef", x"ed", x"f1", x"f3", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"f2", x"f3", x"f2", x"f4", x"ea", x"d2", x"c0", x"ce", x"e2", x"e5", x"e6", x"e6", x"e7", x"e9", x"e6", 
        x"e3", x"e3", x"e3", x"e2", x"e2", x"e4", x"e4", x"e3", x"e2", x"e2", x"e2", x"e3", x"e2", x"e1", x"e4", 
        x"e2", x"e1", x"e3", x"e2", x"e3", x"e0", x"e0", x"e3", x"e2", x"e0", x"df", x"df", x"df", x"e0", x"e1", 
        x"df", x"dd", x"de", x"e1", x"e3", x"e4", x"e4", x"e2", x"e1", x"e2", x"e2", x"e1", x"e0", x"e0", x"e2", 
        x"e1", x"e0", x"e3", x"e3", x"de", x"df", x"de", x"df", x"e1", x"e0", x"e5", x"e2", x"e5", x"dc", x"d0", 
        x"df", x"e1", x"d7", x"d2", x"cb", x"c3", x"b6", x"ae", x"a5", x"96", x"8f", x"7f", x"72", x"6f", x"67", 
        x"60", x"5a", x"53", x"4e", x"4f", x"52", x"55", x"58", x"5c", x"63", x"65", x"64", x"63", x"64", x"65", 
        x"65", x"63", x"5f", x"5e", x"58", x"52", x"46", x"42", x"3c", x"38", x"32", x"2f", x"29", x"20", x"1f", 
        x"1d", x"1c", x"1d", x"1d", x"1e", x"19", x"1e", x"1f", x"18", x"1c", x"25", x"28", x"29", x"28", x"27", 
        x"24", x"22", x"25", x"25", x"2e", x"33", x"3a", x"40", x"4a", x"52", x"53", x"61", x"60", x"5d", x"64", 
        x"67", x"6b", x"6c", x"6c", x"75", x"69", x"5c", x"5b", x"5b", x"57", x"2e", x"09", x"18", x"4a", x"4c", 
        x"7b", x"6e", x"76", x"77", x"64", x"60", x"59", x"5f", x"8a", x"8e", x"55", x"70", x"77", x"61", x"75", 
        x"96", x"6b", x"51", x"63", x"91", x"82", x"56", x"42", x"5f", x"6a", x"61", x"8c", x"76", x"4b", x"4a", 
        x"54", x"4d", x"5c", x"6d", x"50", x"5e", x"76", x"5b", x"5e", x"6c", x"6a", x"52", x"5a", x"73", x"4e", 
        x"39", x"4d", x"5e", x"3e", x"4c", x"69", x"58", x"5c", x"7e", x"82", x"70", x"63", x"38", x"4b", x"56", 
        x"4b", x"55", x"46", x"6f", x"8c", x"66", x"4c", x"65", x"6d", x"73", x"68", x"94", x"7b", x"88", x"6e", 
        x"58", x"73", x"7e", x"ad", x"97", x"8a", x"8b", x"8b", x"ac", x"c1", x"be", x"b7", x"ae", x"a2", x"96", 
        x"b0", x"a9", x"9d", x"a9", x"a0", x"8b", x"d5", x"b3", x"8d", x"71", x"2f", x"27", x"38", x"1e", x"16", 
        x"4d", x"96", x"d9", x"d6", x"d5", x"d7", x"d5", x"d7", x"d7", x"d2", x"d0", x"d1", x"d2", x"d4", x"d5", 
        x"d5", x"d5", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d1", x"d2", x"d3", x"d4", x"d4", x"d3", x"d2", 
        x"d2", x"d1", x"d3", x"d3", x"d5", x"c2", x"8a", x"83", x"87", x"84", x"85", x"83", x"84", x"8d", x"8e", 
        x"89", x"80", x"88", x"cc", x"e4", x"de", x"db", x"db", x"d7", x"e1", x"d6", x"ce", x"d2", x"d3", x"d4", 
        x"d2", x"d1", x"d1", x"d1", x"d1", x"d0", x"cf", x"ce", x"ce", x"cf", x"d0", x"d1", x"d2", x"d2", x"d2", 
        x"d1", x"d0", x"d1", x"d3", x"d5", x"d6", x"d5", x"d5", x"d3", x"d2", x"d1", x"d1", x"d3", x"d3", x"d3", 
        x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d0", x"d1", x"d0", x"cc", x"cf", x"e4", x"c8", x"96", x"7f", 
        x"79", x"7d", x"7a", x"77", x"89", x"ae", x"94", x"7f", x"7b", x"7e", x"88", x"89", x"82", x"7d", x"81", 
        x"86", x"81", x"78", x"77", x"7c", x"7c", x"77", x"6c", x"65", x"6d", x"76", x"77", x"6c", x"66", x"69", 
        x"72", x"78", x"74", x"6d", x"76", x"7f", x"83", x"81", x"7c", x"7d", x"84", x"86", x"7f", x"77", x"79", 
        x"80", x"7f", x"73", x"85", x"ce", x"c8", x"84", x"70", x"7f", x"87", x"83", x"7c", x"81", x"8c", x"94", 
        x"8e", x"85", x"8e", x"98", x"95", x"8b", x"8a", x"92", x"92", x"86", x"79", x"7c", x"83", x"80", x"77", 
        x"78", x"87", x"8e", x"86", x"79", x"7e", x"8a", x"8f", x"88", x"85", x"91", x"9b", x"9a", x"8c", x"a1", 
        x"dc", x"c1", x"90", x"8c", x"8e", x"91", x"8d", x"83", x"7e", x"88", x"8f", x"88", x"82", x"82", x"8b", 
        x"8c", x"85", x"88", x"96", x"9a", x"94", x"92", x"96", x"9d", x"9a", x"96", x"99", x"99", x"92", x"89", 
        x"87", x"8a", x"8b", x"89", x"88", x"8b", x"8c", x"9d", x"cd", x"b7", x"7a", x"7d", x"86", x"8b", x"8a", 
        x"89", x"87", x"85", x"85", x"87", x"88", x"87", x"7d", x"78", x"75", x"6f", x"70", x"77", x"79", x"7e", 
        x"7a", x"76", x"7b", x"81", x"82", x"7e", x"7d", x"83", x"83", x"7b", x"70", x"6d", x"80", x"c0", x"d9", 
        x"b2", x"b3", x"b7", x"ba", x"bb", x"bd", x"bf", x"b7", x"b9", x"bf", x"c2", x"bc", x"b9", x"b8", x"b8", 
        x"b8", x"be", x"bf", x"bc", x"b3", x"b3", x"b7", x"bd", x"bf", x"bc", x"ba", x"ba", x"bb", x"bd", x"bc", 
        x"be", x"d5", x"a4", x"89", x"85", x"84", x"8e", x"8d", x"80", x"78", x"81", x"86", x"7a", x"78", x"7f", 
        x"80", x"78", x"7c", x"89", x"8a", x"81", x"82", x"8b", x"8d", x"8a", x"8c", x"91", x"93", x"91", x"98", 
        x"c5", x"cd", x"9c", x"96", x"95", x"98", x"a2", x"a7", x"a4", x"a6", x"a9", x"aa", x"b0", x"b8", x"b7", 
        x"b2", x"b6", x"be", x"bd", x"ba", x"ba", x"c0", x"c4", x"c4", x"c5", x"cf", x"d3", x"d1", x"d5", x"d9", 
        x"df", x"dc", x"dc", x"e4", x"e7", x"ec", x"f1", x"f0", x"ef", x"f3", x"f6", x"f6", x"f5", x"f6", x"f6", 
        x"f5", x"f3", x"f5", x"f5", x"f1", x"f3", x"f5", x"f3", x"f3", x"f1", x"f0", x"f0", x"f1", x"f2", x"f1", 
        x"f2", x"f4", x"f4", x"f2", x"ef", x"f2", x"f3", x"ef", x"f2", x"f0", x"f1", x"f3", x"f4", x"f4", x"f5", 
        x"f5", x"f6", x"f7", x"f2", x"f4", x"f6", x"f7", x"f4", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f2", 
        x"f0", x"f1", x"f3", x"f3", x"f1", x"f1", x"f2", x"ef", x"ef", x"ef", x"ef", x"ee", x"f0", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"ef", x"f1", 
        x"f3", x"f4", x"f4", x"f4", x"e7", x"e1", x"e1", x"e8", x"e8", x"e4", x"e7", x"e8", x"e9", x"e7", x"e5", 
        x"e5", x"e6", x"e6", x"e4", x"e4", x"e6", x"e6", x"e5", x"e4", x"e4", x"e3", x"e2", x"e1", x"e1", x"e4", 
        x"e3", x"e2", x"e3", x"e0", x"e0", x"e0", x"e1", x"e1", x"df", x"de", x"e1", x"e3", x"e1", x"e1", x"e1", 
        x"df", x"df", x"e1", x"e0", x"e2", x"e4", x"e4", x"e1", x"e0", x"e2", x"e3", x"e1", x"df", x"e0", x"e0", 
        x"df", x"e0", x"e3", x"e8", x"e8", x"e9", x"ea", x"e7", x"e2", x"de", x"d9", x"ce", x"c6", x"b0", x"97", 
        x"99", x"8e", x"7b", x"71", x"6b", x"6a", x"61", x"5d", x"5b", x"54", x"55", x"55", x"53", x"56", x"5c", 
        x"63", x"66", x"65", x"67", x"6c", x"70", x"6e", x"6a", x"69", x"68", x"61", x"5a", x"51", x"48", x"3e", 
        x"38", x"33", x"2d", x"29", x"23", x"20", x"1c", x"1f", x"1e", x"1e", x"1f", x"24", x"27", x"26", x"27", 
        x"28", x"29", x"28", x"28", x"26", x"24", x"39", x"45", x"3f", x"3d", x"3e", x"44", x"48", x"4b", x"4f", 
        x"4f", x"55", x"62", x"5c", x"63", x"69", x"69", x"69", x"67", x"61", x"68", x"7d", x"7c", x"79", x"7e", 
        x"7f", x"84", x"85", x"83", x"84", x"6a", x"56", x"55", x"55", x"54", x"30", x"09", x"12", x"44", x"4c", 
        x"72", x"67", x"8b", x"6e", x"7b", x"84", x"56", x"67", x"83", x"7c", x"57", x"6b", x"74", x"53", x"51", 
        x"78", x"87", x"69", x"4c", x"6c", x"63", x"4e", x"36", x"41", x"3d", x"33", x"64", x"53", x"6b", x"5a", 
        x"5f", x"5d", x"67", x"81", x"77", x"6d", x"59", x"54", x"68", x"58", x"55", x"75", x"76", x"45", x"46", 
        x"32", x"4c", x"61", x"41", x"53", x"62", x"66", x"7c", x"6f", x"5f", x"4a", x"60", x"61", x"5a", x"5f", 
        x"3a", x"55", x"5a", x"58", x"4c", x"5d", x"62", x"54", x"70", x"91", x"a4", x"af", x"94", x"70", x"5f", 
        x"6b", x"75", x"76", x"84", x"89", x"6e", x"6a", x"9d", x"c5", x"dd", x"cb", x"d0", x"d8", x"e2", x"d2", 
        x"c5", x"d2", x"d4", x"cc", x"c9", x"c9", x"ce", x"a1", x"8c", x"72", x"65", x"60", x"57", x"38", x"29", 
        x"4f", x"98", x"dd", x"d6", x"d5", x"d7", x"d5", x"d7", x"d7", x"d2", x"d2", x"d2", x"d2", x"d3", x"d3", 
        x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", x"d3", x"d3", x"d3", x"d2", x"d0", x"d0", x"d2", x"d5", x"d5", 
        x"d0", x"cf", x"d2", x"ce", x"d3", x"c2", x"8b", x"85", x"89", x"8d", x"90", x"8c", x"86", x"7d", x"6b", 
        x"56", x"39", x"5a", x"c4", x"e2", x"db", x"de", x"da", x"d5", x"df", x"d4", x"cc", x"d0", x"d2", x"d4", 
        x"d1", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", x"d1", 
        x"d0", x"d0", x"d1", x"d3", x"d4", x"d4", x"d4", x"d5", x"d4", x"d2", x"d1", x"d1", x"d3", x"d4", x"d3", 
        x"d2", x"d2", x"d3", x"d4", x"d4", x"d3", x"d4", x"d2", x"d0", x"ce", x"cf", x"e1", x"c6", x"93", x"82", 
        x"7b", x"72", x"67", x"67", x"86", x"b7", x"97", x"76", x"73", x"73", x"75", x"74", x"77", x"79", x"7c", 
        x"7f", x"7f", x"7d", x"7e", x"82", x"88", x"88", x"87", x"89", x"8d", x"8d", x"88", x"85", x"82", x"83", 
        x"82", x"7a", x"71", x"6d", x"71", x"73", x"6d", x"64", x"63", x"6a", x"75", x"74", x"6c", x"69", x"71", 
        x"7b", x"7b", x"73", x"81", x"c6", x"d0", x"94", x"86", x"93", x"97", x"8e", x"7d", x"82", x"87", x"85", 
        x"7a", x"72", x"79", x"83", x"81", x"79", x"7b", x"86", x"8b", x"83", x"82", x"8b", x"9a", x"9d", x"92", 
        x"89", x"8f", x"95", x"91", x"87", x"89", x"8f", x"8e", x"84", x"7a", x"7b", x"80", x"86", x"80", x"95", 
        x"d4", x"c0", x"8e", x"89", x"86", x"91", x"98", x"93", x"91", x"96", x"9a", x"97", x"91", x"8f", x"92", 
        x"92", x"8b", x"86", x"87", x"87", x"80", x"7c", x"81", x"8c", x"92", x"8f", x"89", x"88", x"8e", x"91", 
        x"92", x"97", x"9d", x"a1", x"9c", x"94", x"92", x"a0", x"d0", x"c3", x"80", x"78", x"77", x"7b", x"74", 
        x"6d", x"6d", x"73", x"79", x"79", x"77", x"77", x"7d", x"7b", x"7c", x"7d", x"84", x"8c", x"8a", x"86", 
        x"85", x"87", x"87", x"86", x"86", x"82", x"76", x"6e", x"6a", x"6e", x"6c", x"6e", x"78", x"b6", x"dd", 
        x"c0", x"c2", x"c7", x"c8", x"c5", x"bd", x"be", x"c2", x"be", x"b5", x"b5", x"b3", x"b2", x"ac", x"b4", 
        x"ba", x"bc", x"b9", x"ba", x"bb", x"be", x"c1", x"c4", x"c4", x"c0", x"ba", x"ba", x"bd", x"be", x"ba", 
        x"ba", x"d2", x"a2", x"7f", x"80", x"85", x"87", x"81", x"80", x"89", x"8e", x"8a", x"88", x"8e", x"8c", 
        x"86", x"85", x"8b", x"8d", x"81", x"79", x"7e", x"84", x"80", x"7a", x"7f", x"85", x"7f", x"7a", x"85", 
        x"bb", x"c3", x"7f", x"76", x"76", x"76", x"7c", x"7e", x"79", x"75", x"7d", x"85", x"89", x"89", x"88", 
        x"8a", x"8d", x"95", x"9f", x"a3", x"a5", x"a7", x"aa", x"ae", x"b4", x"c0", x"be", x"c2", x"d1", x"c8", 
        x"c7", x"c0", x"b5", x"c3", x"c8", x"c3", x"c1", x"c7", x"cd", x"d1", x"d3", x"d8", x"db", x"dc", x"dd", 
        x"e0", x"e1", x"e7", x"ec", x"e9", x"e9", x"ed", x"f3", x"f4", x"f4", x"f4", x"f3", x"f4", x"f4", x"f0", 
        x"f7", x"f4", x"f1", x"f4", x"f2", x"f3", x"f6", x"f3", x"f3", x"f1", x"f1", x"f3", x"f2", x"f0", x"f3", 
        x"f5", x"f7", x"f7", x"f5", x"f7", x"f6", x"f5", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f3", x"f3", x"f1", x"f0", x"f1", x"ef", x"f0", x"f3", x"f2", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"ee", x"f1", 
        x"f4", x"f4", x"f5", x"f5", x"e5", x"db", x"e2", x"e8", x"e6", x"e8", x"ea", x"e8", x"e7", x"e7", x"e6", 
        x"e6", x"e7", x"e7", x"e4", x"e4", x"e7", x"e7", x"e6", x"e4", x"e3", x"e1", x"e1", x"e2", x"e0", x"e2", 
        x"e2", x"e1", x"e1", x"de", x"dc", x"df", x"e2", x"e2", x"e0", x"df", x"e2", x"e3", x"e2", x"e2", x"e4", 
        x"e3", x"e0", x"e0", x"e3", x"e4", x"e5", x"e5", x"e3", x"e2", x"e2", x"e6", x"e6", x"e5", x"e5", x"df", 
        x"d8", x"d3", x"cc", x"c2", x"ba", x"ab", x"9f", x"91", x"83", x"7d", x"77", x"6d", x"6b", x"69", x"64", 
        x"67", x"61", x"5a", x"5a", x"5f", x"64", x"65", x"68", x"65", x"65", x"68", x"6c", x"70", x"6f", x"70", 
        x"6d", x"68", x"5e", x"55", x"4d", x"45", x"39", x"31", x"2d", x"29", x"24", x"24", x"26", x"27", x"27", 
        x"28", x"28", x"27", x"2a", x"29", x"2a", x"28", x"2d", x"2d", x"29", x"25", x"26", x"29", x"2a", x"2d", 
        x"33", x"3c", x"3e", x"49", x"4a", x"48", x"68", x"77", x"77", x"72", x"6d", x"71", x"70", x"6c", x"6b", 
        x"66", x"66", x"69", x"58", x"54", x"54", x"4a", x"46", x"44", x"3c", x"57", x"84", x"8c", x"86", x"8a", 
        x"87", x"88", x"86", x"85", x"89", x"6b", x"54", x"54", x"56", x"57", x"38", x"10", x"12", x"42", x"4e", 
        x"7a", x"5c", x"79", x"80", x"71", x"6d", x"5b", x"59", x"67", x"69", x"71", x"63", x"55", x"4c", x"35", 
        x"3e", x"61", x"73", x"5b", x"5c", x"62", x"44", x"4a", x"4c", x"4c", x"51", x"43", x"51", x"74", x"53", 
        x"70", x"7f", x"6e", x"6f", x"7c", x"61", x"3a", x"51", x"7d", x"5d", x"58", x"71", x"71", x"75", x"83", 
        x"67", x"77", x"69", x"50", x"58", x"59", x"70", x"89", x"6b", x"4e", x"5d", x"69", x"5b", x"50", x"72", 
        x"5c", x"3c", x"40", x"57", x"51", x"55", x"72", x"61", x"72", x"79", x"90", x"a8", x"8b", x"78", x"7f", 
        x"6b", x"76", x"a9", x"a9", x"ad", x"74", x"87", x"ae", x"d2", x"d1", x"bd", x"dd", x"e4", x"eb", x"c7", 
        x"a7", x"d6", x"e5", x"e9", x"ea", x"e9", x"e5", x"cd", x"b7", x"a3", x"b4", x"b8", x"8b", x"96", x"95", 
        x"7b", x"9d", x"da", x"d6", x"d5", x"d7", x"d5", x"d7", x"d7", x"d3", x"d4", x"d3", x"d2", x"d1", x"d2", 
        x"d2", x"d3", x"d3", x"d3", x"d4", x"d4", x"d2", x"d1", x"cf", x"d3", x"d3", x"d1", x"d0", x"d0", x"d1", 
        x"d0", x"d2", x"d4", x"d3", x"d9", x"c8", x"91", x"85", x"7f", x"70", x"5f", x"4b", x"37", x"2b", x"22", 
        x"1d", x"19", x"46", x"c1", x"e3", x"db", x"e0", x"da", x"d7", x"e0", x"d4", x"cb", x"ce", x"d0", x"d1", 
        x"d1", x"cf", x"cf", x"cf", x"d0", x"d0", x"d1", x"d2", x"d2", x"d1", x"d1", x"d1", x"d0", x"cf", x"d0", 
        x"d0", x"d0", x"d1", x"d2", x"d3", x"d3", x"d3", x"d5", x"d4", x"d2", x"d1", x"d1", x"d2", x"d3", x"d4", 
        x"d2", x"d1", x"d2", x"d4", x"d4", x"d4", x"d5", x"d0", x"cf", x"d0", x"d0", x"e2", x"cb", x"98", x"7f", 
        x"79", x"7b", x"74", x"7b", x"8b", x"a4", x"8b", x"80", x"89", x"87", x"83", x"7e", x"83", x"87", x"82", 
        x"7f", x"80", x"84", x"87", x"83", x"77", x"72", x"75", x"7a", x"79", x"74", x"73", x"7a", x"7f", x"81", 
        x"7e", x"7a", x"7b", x"80", x"83", x"83", x"81", x"7f", x"82", x"86", x"86", x"7f", x"7a", x"7d", x"84", 
        x"87", x"80", x"78", x"86", x"c7", x"c9", x"86", x"78", x"86", x"87", x"7e", x"76", x"81", x"8a", x"89", 
        x"83", x"87", x"93", x"9a", x"93", x"88", x"88", x"91", x"97", x"8f", x"83", x"84", x"8d", x"8a", x"7d", 
        x"75", x"7d", x"86", x"84", x"7b", x"7d", x"86", x"8b", x"86", x"82", x"8e", x"9a", x"a5", x"9b", x"a0", 
        x"d7", x"c6", x"93", x"91", x"8b", x"92", x"96", x"8f", x"89", x"82", x"87", x"88", x"83", x"81", x"88", 
        x"8f", x"8c", x"87", x"89", x"90", x"93", x"90", x"91", x"95", x"9b", x"98", x"91", x"90", x"96", x"98", 
        x"93", x"8f", x"8c", x"8c", x"88", x"82", x"81", x"94", x"ca", x"bd", x"7a", x"72", x"72", x"7f", x"83", 
        x"81", x"82", x"89", x"8f", x"8c", x"84", x"80", x"88", x"8a", x"86", x"7d", x"7a", x"7c", x"76", x"74", 
        x"75", x"79", x"7b", x"80", x"81", x"7a", x"72", x"6e", x"70", x"79", x"77", x"78", x"82", x"b9", x"dc", 
        x"c1", x"bf", x"bd", x"b6", x"b7", x"b3", x"ae", x"b7", x"bb", x"b7", x"b3", x"b4", x"bb", x"bd", x"c0", 
        x"c4", x"c3", x"bd", x"ba", x"be", x"c1", x"bc", x"b8", x"b8", x"b5", x"b1", x"b1", x"b8", x"bd", x"ba", 
        x"ba", x"d3", x"a8", x"82", x"8e", x"96", x"90", x"8a", x"8d", x"92", x"8d", x"87", x"8c", x"8f", x"88", 
        x"81", x"85", x"8c", x"8a", x"82", x"85", x"8b", x"8a", x"84", x"85", x"8c", x"8b", x"85", x"84", x"90", 
        x"bd", x"cb", x"87", x"72", x"73", x"74", x"76", x"76", x"73", x"6f", x"6f", x"73", x"75", x"72", x"73", 
        x"78", x"76", x"72", x"76", x"7c", x"7c", x"7a", x"7e", x"86", x"8c", x"8c", x"8b", x"aa", x"d1", x"b1", 
        x"94", x"8d", x"95", x"a9", x"ae", x"a5", x"a0", x"ad", x"b9", x"b3", x"b2", x"bb", x"c3", x"c0", x"bb", 
        x"bf", x"c8", x"c6", x"c1", x"c3", x"ca", x"d0", x"d4", x"d4", x"d5", x"d6", x"de", x"df", x"e6", x"e6", 
        x"e8", x"e8", x"e9", x"f0", x"f0", x"f0", x"f4", x"f5", x"f4", x"f1", x"ef", x"f3", x"f3", x"f0", x"f3", 
        x"f5", x"f7", x"f5", x"f6", x"f9", x"f7", x"f4", x"f2", x"f1", x"f3", x"f3", x"f3", x"f3", x"f1", x"f1", 
        x"f2", x"f2", x"f1", x"f0", x"f0", x"ef", x"f1", x"f3", x"f1", x"ef", x"f2", x"f0", x"ef", x"f2", x"f0", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f0", x"f0", x"f2", 
        x"f3", x"f3", x"f4", x"f6", x"e5", x"d8", x"e2", x"e7", x"e5", x"e9", x"ea", x"e9", x"e9", x"e7", x"e6", 
        x"e6", x"e7", x"e7", x"e5", x"e4", x"e5", x"e4", x"e4", x"e2", x"e2", x"e1", x"e2", x"e4", x"e2", x"e4", 
        x"e3", x"e4", x"e5", x"e2", x"e0", x"e0", x"e1", x"e3", x"e4", x"e4", x"e3", x"e2", x"e2", x"e2", x"e5", 
        x"e5", x"e3", x"e3", x"e5", x"e4", x"e0", x"dc", x"d7", x"d0", x"c5", x"bd", x"b2", x"a9", x"9f", x"90", 
        x"84", x"7d", x"76", x"71", x"6e", x"69", x"69", x"6a", x"68", x"6a", x"69", x"6a", x"6c", x"70", x"72", 
        x"75", x"77", x"79", x"7a", x"7b", x"78", x"73", x"70", x"67", x"5c", x"52", x"4d", x"49", x"3b", x"33", 
        x"31", x"30", x"29", x"28", x"2a", x"2c", x"2a", x"2a", x"2c", x"2d", x"2c", x"2d", x"2f", x"2e", x"2e", 
        x"30", x"2b", x"28", x"2a", x"2c", x"32", x"39", x"44", x"48", x"48", x"49", x"4f", x"57", x"5f", x"63", 
        x"60", x"66", x"65", x"6c", x"64", x"55", x"72", x"84", x"87", x"7b", x"6d", x"6f", x"6c", x"69", x"67", 
        x"63", x"5b", x"52", x"48", x"49", x"4a", x"44", x"3f", x"43", x"3e", x"56", x"7f", x"85", x"85", x"85", 
        x"82", x"86", x"83", x"81", x"87", x"6b", x"53", x"54", x"54", x"56", x"3a", x"11", x"0d", x"3d", x"4e", 
        x"7f", x"7c", x"70", x"66", x"71", x"81", x"8a", x"6f", x"68", x"5f", x"68", x"63", x"54", x"5f", x"58", 
        x"4f", x"46", x"5f", x"5a", x"60", x"71", x"4d", x"56", x"4e", x"44", x"4f", x"57", x"54", x"72", x"46", 
        x"46", x"51", x"41", x"68", x"68", x"62", x"73", x"75", x"7b", x"5a", x"52", x"69", x"7a", x"7e", x"69", 
        x"79", x"85", x"71", x"6a", x"62", x"61", x"57", x"53", x"5f", x"68", x"6f", x"59", x"42", x"3b", x"58", 
        x"5a", x"38", x"4b", x"86", x"66", x"4e", x"5d", x"4a", x"6f", x"7d", x"81", x"92", x"73", x"7e", x"94", 
        x"73", x"8a", x"a1", x"95", x"a5", x"94", x"97", x"ab", x"cc", x"c2", x"d1", x"e4", x"e7", x"e4", x"cb", 
        x"b0", x"c7", x"c2", x"d9", x"e4", x"da", x"d1", x"d1", x"bd", x"a5", x"be", x"d2", x"ac", x"ce", x"c9", 
        x"b5", x"c5", x"da", x"d5", x"d5", x"d7", x"d5", x"d7", x"d7", x"d2", x"d2", x"d2", x"d1", x"d1", x"d2", 
        x"d3", x"d4", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"ce", x"d1", x"d3", x"d2", x"d1", x"d0", x"d3", 
        x"d9", x"de", x"db", x"cc", x"bd", x"99", x"56", x"35", x"25", x"1e", x"1d", x"1b", x"17", x"18", x"21", 
        x"31", x"40", x"5e", x"c5", x"e5", x"db", x"d9", x"d9", x"d9", x"e2", x"d6", x"cd", x"cf", x"d0", x"d1", 
        x"d0", x"cf", x"cf", x"cf", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", x"d1", x"d2", x"d1", 
        x"d0", x"d1", x"d2", x"d2", x"d3", x"d3", x"d3", x"d5", x"d4", x"d3", x"d2", x"d2", x"d1", x"d2", x"d4", 
        x"d3", x"d1", x"d2", x"d4", x"d5", x"d4", x"d2", x"d2", x"d4", x"d2", x"d1", x"e0", x"c0", x"8c", x"78", 
        x"70", x"68", x"58", x"69", x"90", x"bd", x"9a", x"79", x"6d", x"60", x"5c", x"5f", x"66", x"62", x"5d", 
        x"60", x"6c", x"78", x"7b", x"78", x"78", x"7d", x"8c", x"97", x"90", x"87", x"86", x"8c", x"8e", x"87", 
        x"7d", x"7d", x"84", x"89", x"7d", x"71", x"68", x"67", x"6f", x"72", x"6d", x"63", x"62", x"6e", x"78", 
        x"79", x"73", x"6f", x"79", x"b7", x"d1", x"9b", x"92", x"9a", x"93", x"8c", x"8f", x"97", x"99", x"8a", 
        x"77", x"75", x"7a", x"79", x"6f", x"6a", x"71", x"7c", x"83", x"7c", x"73", x"79", x"88", x"8d", x"89", 
        x"8b", x"9a", x"a0", x"9d", x"91", x"90", x"96", x"9c", x"97", x"89", x"80", x"85", x"91", x"88", x"92", 
        x"d4", x"c1", x"81", x"82", x"7c", x"82", x"89", x"89", x"8b", x"8c", x"98", x"a5", x"a2", x"9a", x"94", 
        x"96", x"97", x"92", x"8d", x"90", x"92", x"89", x"82", x"7f", x"82", x"82", x"80", x"83", x"8b", x"8e", 
        x"8c", x"89", x"89", x"93", x"9e", x"9e", x"93", x"9a", x"ce", x"c5", x"84", x"7c", x"79", x"80", x"81", 
        x"7c", x"77", x"75", x"75", x"72", x"6c", x"6a", x"73", x"7b", x"7b", x"74", x"74", x"7e", x"84", x"8c", 
        x"8a", x"8a", x"93", x"a3", x"a1", x"8d", x"7c", x"7f", x"8a", x"89", x"75", x"6b", x"7b", x"b8", x"d8", 
        x"b1", x"a9", x"ad", x"ad", x"ae", x"ad", x"b7", x"bc", x"c1", x"c0", x"be", x"bb", x"bf", x"c2", x"bc", 
        x"b6", x"b3", x"b5", x"b1", x"ad", x"ad", x"b3", x"b5", x"b1", x"b3", x"ba", x"bf", x"c1", x"c4", x"c3", 
        x"c0", x"d9", x"b6", x"92", x"91", x"87", x"83", x"84", x"81", x"7b", x"7c", x"81", x"87", x"87", x"83", 
        x"87", x"90", x"92", x"8b", x"88", x"90", x"91", x"87", x"81", x"84", x"87", x"7d", x"79", x"7f", x"8b", 
        x"b2", x"cc", x"90", x"7b", x"7e", x"7e", x"7f", x"82", x"82", x"7f", x"80", x"7f", x"79", x"75", x"75", 
        x"77", x"74", x"73", x"75", x"76", x"73", x"6f", x"6f", x"72", x"74", x"74", x"70", x"9d", x"d7", x"ab", 
        x"7b", x"76", x"74", x"77", x"76", x"70", x"70", x"76", x"78", x"77", x"75", x"7c", x"87", x"8a", x"8f", 
        x"9c", x"a6", x"9d", x"98", x"a8", x"bb", x"bc", x"b2", x"b8", x"cd", x"c2", x"bb", x"bd", x"c1", x"bb", 
        x"b8", x"bc", x"c5", x"ca", x"cd", x"d0", x"d3", x"d5", x"dd", x"e2", x"e1", x"e5", x"e8", x"e9", x"f0", 
        x"f4", x"f6", x"f1", x"f4", x"f9", x"f8", x"f6", x"f3", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f0", 
        x"f1", x"f3", x"f2", x"f2", x"f3", x"f3", x"f1", x"f1", x"f0", x"ee", x"f1", x"ef", x"ed", x"f2", x"ef", 
        x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", 
        x"f3", x"f2", x"f3", x"f6", x"e8", x"d5", x"e3", x"eb", x"e9", x"e8", x"e6", x"e8", x"e8", x"e7", x"e4", 
        x"e5", x"e7", x"e8", x"e6", x"e6", x"e6", x"e6", x"e4", x"e2", x"e1", x"e0", x"e1", x"e5", x"e2", x"e3", 
        x"e4", x"e3", x"e4", x"e1", x"e2", x"e1", x"e0", x"e2", x"e7", x"e7", x"e2", x"e4", x"e2", x"de", x"db", 
        x"d1", x"c5", x"bc", x"b0", x"a3", x"94", x"86", x"7f", x"78", x"70", x"6d", x"6c", x"6c", x"6f", x"71", 
        x"72", x"75", x"75", x"75", x"74", x"73", x"78", x"7d", x"7e", x"81", x"83", x"83", x"7d", x"77", x"71", 
        x"69", x"61", x"5a", x"4f", x"47", x"3c", x"33", x"2e", x"2a", x"2a", x"2a", x"33", x"30", x"16", x"0b", 
        x"21", x"3c", x"40", x"3e", x"3d", x"3b", x"36", x"34", x"30", x"2a", x"2a", x"2d", x"33", x"3a", x"43", 
        x"4b", x"4d", x"52", x"5c", x"63", x"68", x"69", x"6e", x"70", x"6f", x"6c", x"66", x"61", x"60", x"5b", 
        x"51", x"55", x"52", x"51", x"48", x"3f", x"68", x"7e", x"82", x"7b", x"70", x"72", x"6f", x"6b", x"69", 
        x"66", x"5d", x"4c", x"4b", x"4e", x"4c", x"49", x"44", x"47", x"41", x"58", x"82", x"84", x"82", x"83", 
        x"83", x"88", x"85", x"82", x"89", x"72", x"55", x"56", x"55", x"56", x"3d", x"14", x"0c", x"36", x"4c", 
        x"72", x"9d", x"7c", x"5b", x"7b", x"86", x"83", x"7a", x"68", x"54", x"57", x"4a", x"49", x"7a", x"7c", 
        x"7a", x"59", x"4f", x"4f", x"4e", x"60", x"62", x"59", x"5d", x"3d", x"32", x"48", x"44", x"4e", x"78", 
        x"73", x"4c", x"3c", x"5c", x"70", x"74", x"6f", x"6e", x"4c", x"2e", x"32", x"62", x"73", x"65", x"3f", 
        x"5b", x"77", x"6e", x"47", x"54", x"62", x"86", x"6b", x"73", x"57", x"71", x"6c", x"46", x"5a", x"64", 
        x"58", x"6d", x"78", x"6c", x"48", x"70", x"8d", x"8e", x"87", x"77", x"84", x"9d", x"82", x"94", x"92", 
        x"7f", x"7b", x"6e", x"96", x"8f", x"a0", x"ac", x"b9", x"b8", x"bb", x"ce", x"df", x"e4", x"e7", x"e5", 
        x"dd", x"e5", x"ce", x"ae", x"a0", x"8a", x"ac", x"bf", x"c4", x"a9", x"90", x"c2", x"b0", x"a1", x"bb", 
        x"ce", x"a1", x"d3", x"d5", x"d5", x"d7", x"d5", x"d7", x"d7", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", 
        x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d3", x"d5", x"d7", x"d6", x"d4", x"d4", x"d2", x"c9", x"b5", 
        x"9c", x"80", x"5e", x"3a", x"21", x"17", x"12", x"17", x"1a", x"22", x"2e", x"40", x"54", x"64", x"6e", 
        x"75", x"6e", x"71", x"be", x"df", x"da", x"db", x"dc", x"d9", x"e2", x"d6", x"cd", x"cf", x"cf", x"cf", 
        x"d0", x"d0", x"d1", x"d1", x"d0", x"cf", x"ce", x"ce", x"cf", x"d0", x"d1", x"d2", x"d3", x"d3", x"d2", 
        x"d0", x"d2", x"d4", x"d3", x"d3", x"d3", x"d3", x"d5", x"d5", x"d4", x"d3", x"d2", x"d1", x"d1", x"d6", 
        x"d4", x"d2", x"d3", x"d5", x"d6", x"d5", x"d3", x"d1", x"d3", x"d3", x"d1", x"e3", x"ce", x"9e", x"84", 
        x"7e", x"8a", x"87", x"84", x"83", x"9f", x"8e", x"7d", x"7c", x"7c", x"86", x"8c", x"8d", x"89", x"86", 
        x"87", x"89", x"89", x"81", x"7b", x"78", x"77", x"72", x"6a", x"5f", x"60", x"66", x"6b", x"69", x"61", 
        x"5e", x"6b", x"76", x"74", x"72", x"72", x"77", x"83", x"8d", x"8e", x"89", x"7f", x"7f", x"88", x"88", 
        x"81", x"78", x"73", x"84", x"c7", x"d1", x"8a", x"79", x"7f", x"77", x"74", x"7f", x"86", x"8b", x"85", 
        x"83", x"92", x"9b", x"99", x"8d", x"8b", x"94", x"97", x"92", x"85", x"89", x"92", x"99", x"90", x"7e", 
        x"74", x"7a", x"7c", x"78", x"6e", x"6d", x"78", x"84", x"82", x"78", x"7a", x"87", x"9c", x"a3", x"a3", 
        x"d3", x"cb", x"a1", x"a2", x"9c", x"9c", x"a0", x"9f", x"9d", x"92", x"8d", x"8b", x"84", x"80", x"7e", 
        x"82", x"83", x"84", x"82", x"85", x"8d", x"8b", x"88", x"8c", x"98", x"a5", x"a5", x"9b", x"93", x"91", 
        x"95", x"97", x"94", x"8f", x"8e", x"8d", x"83", x"8c", x"c6", x"c7", x"7f", x"73", x"77", x"76", x"75", 
        x"7a", x"7a", x"79", x"7a", x"7f", x"84", x"86", x"82", x"7e", x"7d", x"79", x"75", x"77", x"79", x"7c", 
        x"82", x"88", x"8e", x"98", x"8c", x"7a", x"66", x"66", x"6f", x"78", x"71", x"69", x"73", x"b2", x"df", 
        x"c4", x"b8", x"b8", x"bd", x"c2", x"bb", x"ba", x"bf", x"bd", x"b2", x"ac", x"af", x"b8", x"b3", x"ac", 
        x"ae", x"b1", x"b1", x"af", x"b5", x"bc", x"be", x"bc", x"ba", x"ba", x"bd", x"c0", x"c2", x"bf", x"b6", 
        x"b4", x"d0", x"ae", x"7f", x"7f", x"81", x"87", x"87", x"82", x"84", x"90", x"97", x"92", x"8c", x"8f", 
        x"93", x"8d", x"86", x"84", x"87", x"86", x"7f", x"7d", x"85", x"8b", x"85", x"7f", x"83", x"92", x"94", 
        x"b9", x"da", x"9a", x"7f", x"82", x"81", x"7e", x"7f", x"80", x"7d", x"7e", x"7f", x"7d", x"7c", x"7e", 
        x"81", x"81", x"81", x"80", x"7e", x"80", x"82", x"81", x"7e", x"7d", x"7f", x"7a", x"9b", x"d8", x"ae", 
        x"74", x"71", x"6f", x"72", x"76", x"72", x"6d", x"70", x"71", x"75", x"75", x"77", x"79", x"74", x"6e", 
        x"70", x"6b", x"66", x"66", x"6c", x"71", x"6f", x"6a", x"83", x"c1", x"ab", x"87", x"91", x"94", x"8c", 
        x"92", x"9c", x"9e", x"9e", x"a7", x"b0", x"b1", x"b4", x"b7", x"bc", x"b7", x"b9", x"be", x"bd", x"c0", 
        x"c8", x"d0", x"cd", x"d2", x"d7", x"da", x"dd", x"e0", x"e1", x"e3", x"e5", x"e7", x"ea", x"ed", x"ec", 
        x"ed", x"ef", x"ed", x"ee", x"f1", x"f0", x"ee", x"f1", x"f2", x"f1", x"f5", x"f0", x"ef", x"f4", x"f1", 
        x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f3", x"f3", 
        x"f3", x"f3", x"f2", x"f6", x"eb", x"d4", x"e2", x"eb", x"e8", x"e6", x"e6", x"e8", x"e8", x"e7", x"e6", 
        x"e6", x"e7", x"e8", x"e5", x"e5", x"e7", x"e8", x"e8", x"e7", x"e7", x"e5", x"e4", x"e5", x"e3", x"e6", 
        x"e8", x"e7", x"e5", x"df", x"da", x"d6", x"cf", x"c7", x"be", x"b3", x"a6", x"9d", x"93", x"86", x"7e", 
        x"78", x"74", x"73", x"74", x"75", x"78", x"7d", x"81", x"83", x"82", x"83", x"86", x"85", x"86", x"88", 
        x"86", x"86", x"87", x"81", x"7b", x"75", x"6d", x"65", x"5e", x"57", x"4a", x"42", x"3a", x"30", x"38", 
        x"39", x"22", x"2c", x"2c", x"33", x"37", x"39", x"3c", x"3b", x"40", x"40", x"43", x"3e", x"1a", x"05", 
        x"22", x"3f", x"3d", x"3d", x"41", x"47", x"4e", x"56", x"61", x"6d", x"6c", x"6b", x"6e", x"72", x"73", 
        x"73", x"71", x"6c", x"69", x"64", x"5f", x"58", x"59", x"55", x"52", x"4e", x"45", x"41", x"48", x"49", 
        x"3d", x"45", x"4d", x"4e", x"4b", x"41", x"67", x"82", x"88", x"82", x"7a", x"76", x"71", x"6f", x"69", 
        x"67", x"61", x"51", x"4e", x"4f", x"4d", x"48", x"42", x"47", x"3d", x"4f", x"81", x"86", x"83", x"85", 
        x"85", x"85", x"83", x"81", x"86", x"73", x"54", x"56", x"56", x"58", x"40", x"16", x"09", x"34", x"4e", 
        x"3c", x"74", x"67", x"75", x"6f", x"69", x"7d", x"7d", x"5f", x"5f", x"5e", x"4e", x"75", x"86", x"63", 
        x"83", x"64", x"3f", x"48", x"38", x"43", x"44", x"3a", x"57", x"6a", x"61", x"74", x"68", x"48", x"5d", 
        x"6e", x"48", x"24", x"52", x"62", x"3f", x"36", x"41", x"55", x"4c", x"51", x"5e", x"4b", x"6b", x"7b", 
        x"81", x"7d", x"6d", x"5c", x"6e", x"66", x"78", x"6b", x"5e", x"4d", x"67", x"6e", x"58", x"50", x"45", 
        x"5a", x"83", x"70", x"60", x"5d", x"66", x"71", x"95", x"90", x"6f", x"72", x"77", x"6e", x"93", x"81", 
        x"73", x"68", x"6e", x"85", x"77", x"ac", x"dd", x"c4", x"9a", x"a5", x"b7", x"db", x"d3", x"dc", x"e9", 
        x"eb", x"ec", x"df", x"c1", x"ad", x"a5", x"9b", x"9b", x"c6", x"c3", x"b1", x"c8", x"be", x"94", x"cd", 
        x"ba", x"7b", x"cb", x"d6", x"d6", x"d6", x"d5", x"d6", x"d8", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", 
        x"d1", x"d2", x"d3", x"d5", x"d6", x"d6", x"d3", x"cf", x"c9", x"b7", x"a3", x"88", x"66", x"47", x"2b", 
        x"1b", x"19", x"19", x"1f", x"25", x"2c", x"3e", x"53", x"62", x"6f", x"75", x"78", x"77", x"74", x"70", 
        x"6d", x"63", x"65", x"ba", x"e1", x"db", x"dd", x"d8", x"d6", x"e0", x"d4", x"cb", x"ce", x"cd", x"ce", 
        x"d0", x"d0", x"d1", x"d1", x"d1", x"cf", x"cd", x"cf", x"d0", x"d0", x"d1", x"d2", x"d2", x"d2", x"d1", 
        x"d1", x"d3", x"d4", x"d3", x"d2", x"d2", x"d3", x"d4", x"d4", x"d4", x"d4", x"d3", x"d1", x"d2", x"d6", 
        x"d4", x"d2", x"d3", x"d5", x"d6", x"d5", x"d4", x"d3", x"d3", x"d1", x"d1", x"e0", x"c1", x"8a", x"78", 
        x"6f", x"68", x"60", x"69", x"83", x"b5", x"99", x"75", x"6d", x"6c", x"6f", x"66", x"5e", x"5f", x"67", 
        x"6c", x"69", x"65", x"68", x"6f", x"75", x"7c", x"7d", x"7b", x"7d", x"86", x"8d", x"8d", x"86", x"7d", 
        x"7e", x"88", x"8a", x"7f", x"73", x"72", x"75", x"76", x"6f", x"65", x"60", x"64", x"6c", x"6c", x"65", 
        x"5f", x"61", x"66", x"75", x"b7", x"d6", x"a2", x"98", x"9b", x"8f", x"89", x"91", x"96", x"97", x"8c", 
        x"85", x"8c", x"8f", x"89", x"79", x"77", x"80", x"84", x"81", x"77", x"7b", x"85", x"8b", x"86", x"82", 
        x"88", x"98", x"9e", x"99", x"8d", x"8b", x"93", x"9b", x"95", x"8b", x"8c", x"95", x"a4", x"9e", x"9d", 
        x"d3", x"c5", x"87", x"88", x"84", x"85", x"89", x"89", x"89", x"89", x"8a", x"92", x"96", x"98", x"9a", 
        x"9f", x"9e", x"9e", x"98", x"94", x"98", x"9b", x"9b", x"97", x"90", x"8d", x"8c", x"8a", x"85", x"83", 
        x"85", x"88", x"88", x"85", x"89", x"90", x"8d", x"92", x"c8", x"d0", x"87", x"7b", x"85", x"89", x"83", 
        x"7d", x"82", x"84", x"81", x"7e", x"7e", x"7e", x"7d", x"72", x"6e", x"70", x"73", x"76", x"76", x"7a", 
        x"8c", x"9c", x"9b", x"9c", x"93", x"8e", x"82", x"7f", x"7a", x"77", x"75", x"74", x"80", x"b6", x"dd", 
        x"c3", x"ba", x"b6", x"b6", x"c0", x"be", x"b8", x"b6", x"b9", x"bd", x"bb", x"b8", x"be", x"c4", x"bb", 
        x"b8", x"b8", x"bf", x"be", x"bb", x"be", x"c1", x"bd", x"b5", x"b6", x"ba", x"bb", x"b7", x"b5", x"b2", 
        x"b2", x"cd", x"af", x"85", x"8a", x"8f", x"92", x"8a", x"85", x"8d", x"91", x"8c", x"82", x"82", x"86", 
        x"87", x"82", x"81", x"87", x"8c", x"87", x"83", x"8b", x"94", x"91", x"85", x"86", x"8e", x"93", x"87", 
        x"ad", x"d8", x"97", x"79", x"7e", x"7f", x"7e", x"81", x"84", x"84", x"82", x"84", x"82", x"7c", x"7d", 
        x"85", x"88", x"85", x"80", x"7b", x"7d", x"7f", x"7d", x"7b", x"7d", x"83", x"82", x"9a", x"d6", x"b7", 
        x"7e", x"7d", x"76", x"79", x"80", x"7f", x"79", x"7b", x"7b", x"74", x"73", x"73", x"73", x"73", x"73", 
        x"71", x"73", x"6f", x"6a", x"6b", x"70", x"72", x"71", x"82", x"c4", x"ab", x"70", x"6f", x"70", x"67", 
        x"6a", x"6f", x"69", x"67", x"73", x"7a", x"79", x"80", x"8e", x"91", x"8f", x"9b", x"aa", x"a8", x"a7", 
        x"b8", x"c0", x"bc", x"cb", x"cc", x"c1", x"c2", x"bb", x"b9", x"bd", x"bd", x"bc", x"c2", x"c8", x"cb", 
        x"ce", x"d4", x"d5", x"d4", x"da", x"de", x"dc", x"e1", x"e4", x"e5", x"e9", x"e5", x"e5", x"ee", x"ec", 
        x"ee", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", x"f2", x"f3", x"f2", x"f2", x"f1", x"f2", x"f4", x"f3", 
        x"f3", x"f3", x"f2", x"f5", x"eb", x"d2", x"df", x"e7", x"e5", x"e4", x"e9", x"ea", x"e8", x"ea", x"e9", 
        x"e9", x"e9", x"e8", x"e5", x"e4", x"e4", x"e4", x"e5", x"e3", x"e0", x"dc", x"d9", x"d6", x"cf", x"c7", 
        x"bf", x"b6", x"ad", x"a2", x"92", x"8c", x"85", x"7f", x"7e", x"7e", x"7c", x"84", x"86", x"86", x"8a", 
        x"8e", x"8d", x"8c", x"8d", x"8e", x"8e", x"8d", x"89", x"84", x"82", x"7e", x"7a", x"71", x"6e", x"6a", 
        x"5e", x"53", x"4f", x"45", x"3d", x"36", x"2f", x"2f", x"32", x"33", x"3b", x"4d", x"63", x"68", x"70", 
        x"66", x"42", x"43", x"44", x"45", x"41", x"3e", x"3d", x"39", x"3d", x"3e", x"42", x"42", x"1d", x"0a", 
        x"3c", x"6c", x"70", x"72", x"76", x"77", x"76", x"75", x"79", x"7f", x"75", x"6a", x"64", x"63", x"5d", 
        x"58", x"57", x"53", x"51", x"50", x"52", x"50", x"52", x"51", x"4f", x"4e", x"48", x"47", x"4e", x"4f", 
        x"45", x"4a", x"4d", x"4d", x"4c", x"41", x"65", x"85", x"8a", x"84", x"79", x"74", x"70", x"70", x"6b", 
        x"67", x"61", x"50", x"4b", x"4c", x"50", x"4d", x"47", x"47", x"41", x"4f", x"80", x"87", x"84", x"82", 
        x"82", x"83", x"84", x"83", x"85", x"73", x"52", x"54", x"56", x"59", x"43", x"18", x"0a", x"36", x"50", 
        x"43", x"69", x"56", x"40", x"56", x"6f", x"69", x"7b", x"71", x"67", x"72", x"5e", x"5a", x"54", x"46", 
        x"5d", x"51", x"3a", x"43", x"49", x"36", x"3c", x"3e", x"5c", x"71", x"88", x"6c", x"50", x"4f", x"63", 
        x"66", x"64", x"39", x"3c", x"47", x"45", x"3b", x"44", x"7d", x"6d", x"4a", x"36", x"54", x"77", x"73", 
        x"6c", x"5f", x"4b", x"61", x"7f", x"68", x"67", x"59", x"51", x"6d", x"69", x"65", x"72", x"53", x"39", 
        x"3b", x"5a", x"45", x"48", x"64", x"5d", x"5f", x"7f", x"74", x"74", x"61", x"68", x"77", x"85", x"8b", 
        x"80", x"74", x"7f", x"5f", x"77", x"ae", x"d1", x"a8", x"9c", x"ab", x"ba", x"c6", x"d3", x"e0", x"e6", 
        x"e5", x"e3", x"e6", x"da", x"d2", x"d3", x"c6", x"ca", x"c9", x"af", x"a1", x"98", x"ca", x"ad", x"bd", 
        x"90", x"8d", x"cd", x"d8", x"d8", x"d5", x"d5", x"d5", x"d8", x"d1", x"cf", x"d0", x"d3", x"d5", x"d5", 
        x"d7", x"d8", x"d2", x"cc", x"bd", x"a8", x"8c", x"73", x"57", x"36", x"21", x"19", x"17", x"1e", x"22", 
        x"2c", x"3a", x"45", x"5e", x"7c", x"7e", x"7b", x"7a", x"79", x"75", x"71", x"6d", x"6b", x"6a", x"69", 
        x"69", x"5f", x"64", x"ba", x"e3", x"d9", x"db", x"db", x"d8", x"e0", x"d6", x"cc", x"ce", x"cf", x"cf", 
        x"cf", x"ce", x"ce", x"cf", x"d1", x"d0", x"cf", x"d0", x"d1", x"d0", x"d0", x"d2", x"d3", x"d2", x"d1", 
        x"d2", x"d3", x"d2", x"d1", x"d1", x"d2", x"d4", x"d4", x"d4", x"d4", x"d4", x"d5", x"d5", x"d5", x"d5", 
        x"d3", x"d2", x"d3", x"d4", x"d4", x"d4", x"d4", x"d6", x"d2", x"d0", x"ce", x"e2", x"ce", x"9d", x"86", 
        x"81", x"82", x"7d", x"77", x"79", x"9c", x"86", x"72", x"7e", x"83", x"82", x"7e", x"7b", x"7c", x"83", 
        x"84", x"7c", x"73", x"76", x"7e", x"80", x"78", x"6d", x"6a", x"68", x"6b", x"69", x"61", x"5c", x"5d", 
        x"66", x"6c", x"6a", x"64", x"66", x"6d", x"73", x"7a", x"7b", x"77", x"79", x"81", x"8a", x"88", x"7f", 
        x"78", x"7e", x"84", x"8a", x"c1", x"d7", x"9a", x"80", x"79", x"70", x"76", x"81", x"84", x"81", x"77", 
        x"79", x"84", x"89", x"88", x"81", x"8d", x"9b", x"a0", x"9b", x"8a", x"8c", x"97", x"9a", x"97", x"8e", 
        x"85", x"89", x"8b", x"85", x"78", x"77", x"82", x"8b", x"89", x"7e", x"7a", x"81", x"89", x"89", x"93", 
        x"ce", x"cf", x"99", x"9a", x"97", x"94", x"97", x"9a", x"9a", x"96", x"93", x"9a", x"9b", x"95", x"8c", 
        x"82", x"84", x"87", x"86", x"83", x"84", x"87", x"86", x"85", x"88", x"8e", x"95", x"98", x"96", x"97", 
        x"9b", x"9f", x"9e", x"99", x"96", x"99", x"9c", x"a2", x"cc", x"d1", x"86", x"77", x"72", x"76", x"73", 
        x"6b", x"6c", x"71", x"74", x"74", x"72", x"74", x"7a", x"7c", x"7c", x"7a", x"80", x"89", x"8b", x"94", 
        x"98", x"a1", x"98", x"9d", x"95", x"86", x"75", x"74", x"6b", x"60", x"65", x"69", x"73", x"ae", x"db", 
        x"bb", x"bf", x"c4", x"c7", x"c6", x"c0", x"c2", x"bc", x"b9", x"be", x"c3", x"be", x"b7", x"b7", x"b8", 
        x"bc", x"b6", x"ba", x"bc", x"bb", x"b7", x"b8", x"bd", x"bf", x"c1", x"be", x"c2", x"c1", x"be", x"b5", 
        x"b4", x"cf", x"b6", x"8e", x"98", x"94", x"87", x"82", x"88", x"8d", x"8a", x"84", x"84", x"87", x"8b", 
        x"8a", x"89", x"8f", x"95", x"8f", x"87", x"8b", x"93", x"8c", x"7f", x"7a", x"7e", x"89", x"85", x"81", 
        x"a9", x"d8", x"94", x"7b", x"82", x"85", x"87", x"88", x"87", x"85", x"85", x"86", x"80", x"78", x"79", 
        x"81", x"84", x"81", x"7c", x"79", x"80", x"83", x"7f", x"7d", x"83", x"86", x"83", x"97", x"d4", x"bb", 
        x"81", x"87", x"81", x"7e", x"80", x"81", x"7e", x"7b", x"7b", x"7c", x"7d", x"78", x"79", x"7f", x"7c", 
        x"72", x"74", x"75", x"73", x"72", x"73", x"74", x"72", x"83", x"c2", x"af", x"74", x"72", x"77", x"6e", 
        x"69", x"6e", x"70", x"6d", x"70", x"74", x"6f", x"68", x"6e", x"70", x"6e", x"6f", x"73", x"6e", x"6d", 
        x"7d", x"80", x"87", x"c7", x"cd", x"a8", x"ac", x"ab", x"ab", x"b4", x"b0", x"a7", x"b2", x"bf", x"bb", 
        x"b5", x"c1", x"c1", x"b4", x"b8", x"c2", x"bb", x"b2", x"ba", x"c2", x"c0", x"c1", x"c6", x"d2", x"d1", 
        x"d5", x"da", x"de", x"df", x"e0", x"e1", x"e2", x"e7", x"eb", x"ea", x"eb", x"ee", x"f2", x"f2", x"f0", 
        x"f2", x"f2", x"f0", x"f2", x"ec", x"d4", x"e3", x"e7", x"e7", x"e8", x"ea", x"ea", x"e8", x"e9", x"e8", 
        x"e3", x"e1", x"db", x"d9", x"d8", x"cd", x"c8", x"c3", x"b9", x"b3", x"a9", x"a0", x"99", x"93", x"8d", 
        x"8a", x"8a", x"8e", x"90", x"93", x"95", x"97", x"98", x"99", x"99", x"99", x"98", x"96", x"93", x"8e", 
        x"8c", x"84", x"7d", x"7a", x"73", x"6b", x"67", x"5c", x"53", x"4f", x"42", x"2c", x"16", x"2d", x"42", 
        x"41", x"44", x"49", x"4b", x"52", x"51", x"50", x"4f", x"4c", x"4c", x"4e", x"52", x"58", x"5a", x"5c", 
        x"48", x"42", x"4a", x"4e", x"50", x"5a", x"58", x"59", x"5e", x"62", x"66", x"6c", x"6c", x"30", x"06", 
        x"3d", x"70", x"6a", x"65", x"64", x"62", x"5f", x"5d", x"5d", x"67", x"67", x"5f", x"5a", x"5d", x"58", 
        x"57", x"58", x"56", x"54", x"54", x"56", x"55", x"54", x"53", x"4b", x"45", x"48", x"4d", x"4f", x"4d", 
        x"44", x"4b", x"50", x"51", x"4f", x"41", x"63", x"87", x"89", x"86", x"79", x"78", x"76", x"74", x"6d", 
        x"6a", x"63", x"52", x"50", x"4e", x"4f", x"4c", x"47", x"46", x"42", x"4a", x"7e", x"88", x"81", x"82", 
        x"84", x"82", x"82", x"84", x"83", x"75", x"55", x"54", x"54", x"57", x"46", x"19", x"08", x"22", x"31", 
        x"5f", x"60", x"4f", x"38", x"56", x"75", x"68", x"66", x"64", x"6a", x"a0", x"8d", x"68", x"5b", x"62", 
        x"5e", x"43", x"54", x"70", x"8f", x"57", x"4f", x"4c", x"66", x"4b", x"4b", x"32", x"28", x"35", x"47", 
        x"39", x"50", x"44", x"4c", x"4b", x"3f", x"71", x"56", x"5c", x"69", x"59", x"4a", x"5a", x"64", x"4b", 
        x"56", x"5c", x"4c", x"5d", x"66", x"69", x"7b", x"7f", x"64", x"59", x"4a", x"4f", x"46", x"51", x"55", 
        x"38", x"48", x"4c", x"40", x"45", x"60", x"72", x"87", x"71", x"78", x"6e", x"71", x"7b", x"83", x"80", 
        x"78", x"87", x"85", x"5e", x"83", x"93", x"a2", x"87", x"8b", x"93", x"8d", x"b2", x"bd", x"dd", x"ef", 
        x"e4", x"e3", x"e5", x"d7", x"c6", x"bc", x"cc", x"e0", x"d3", x"a4", x"92", x"90", x"cc", x"92", x"a1", 
        x"ac", x"ab", x"d9", x"d9", x"d7", x"d7", x"d7", x"d9", x"dc", x"d7", x"d5", x"d8", x"d4", x"ca", x"bb", 
        x"a5", x"8d", x"72", x"55", x"36", x"1e", x"12", x"12", x"24", x"21", x"28", x"3a", x"47", x"5b", x"69", 
        x"72", x"75", x"76", x"7f", x"93", x"88", x"75", x"70", x"6f", x"6c", x"6a", x"68", x"68", x"68", x"68", 
        x"69", x"62", x"66", x"bb", x"e5", x"d9", x"d9", x"d9", x"d7", x"e0", x"d6", x"cc", x"d0", x"cf", x"cf", 
        x"cf", x"ce", x"ce", x"cf", x"d1", x"d0", x"d0", x"d0", x"d1", x"d0", x"d0", x"d1", x"d2", x"d2", x"d1", 
        x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", x"d3", x"d4", x"d4", x"d3", x"d3", x"d4", x"d4", x"d4", x"d4", 
        x"d2", x"d1", x"d2", x"d3", x"d3", x"d3", x"d1", x"d4", x"d1", x"cf", x"d0", x"df", x"c1", x"8a", x"76", 
        x"72", x"72", x"74", x"73", x"86", x"b9", x"a1", x"83", x"84", x"7f", x"77", x"72", x"71", x"74", x"78", 
        x"76", x"6c", x"65", x"6c", x"74", x"72", x"6f", x"6d", x"73", x"7d", x"82", x"7e", x"78", x"75", x"79", 
        x"7f", x"81", x"7c", x"79", x"78", x"77", x"77", x"7a", x"75", x"69", x"65", x"6a", x"6a", x"5e", x"59", 
        x"5d", x"67", x"68", x"72", x"b8", x"db", x"a3", x"91", x"90", x"90", x"99", x"9e", x"9a", x"92", x"8d", 
        x"95", x"9c", x"9a", x"8b", x"7f", x"80", x"81", x"80", x"7d", x"74", x"7f", x"8a", x"87", x"82", x"7c", 
        x"7a", x"86", x"8e", x"90", x"8c", x"8f", x"98", x"9f", x"9c", x"90", x"87", x"8f", x"98", x"99", x"a0", 
        x"d6", x"d1", x"8f", x"89", x"82", x"80", x"85", x"8a", x"8c", x"8d", x"86", x"88", x"8c", x"8e", x"8f", 
        x"8d", x"93", x"9a", x"9b", x"96", x"92", x"93", x"95", x"97", x"92", x"8f", x"92", x"96", x"92", x"89", 
        x"84", x"86", x"87", x"88", x"89", x"89", x"88", x"8e", x"c1", x"d1", x"85", x"74", x"74", x"7d", x"80", 
        x"86", x"82", x"83", x"87", x"87", x"82", x"7e", x"7b", x"7d", x"7d", x"74", x"71", x"7e", x"89", x"90", 
        x"8b", x"8f", x"86", x"8f", x"8f", x"83", x"6b", x"6f", x"79", x"7a", x"74", x"6a", x"76", x"af", x"db", 
        x"be", x"bc", x"bb", x"c0", x"be", x"b4", x"b2", x"b3", x"b7", x"bd", x"be", x"bf", x"c3", x"c1", x"bf", 
        x"c6", x"c7", x"c8", x"c2", x"bd", x"bf", x"b9", x"b9", x"be", x"c2", x"be", x"b9", x"b7", x"b9", x"bb", 
        x"b9", x"cd", x"b4", x"89", x"8b", x"85", x"86", x"8e", x"96", x"96", x"8f", x"8f", x"95", x"90", x"8a", 
        x"8c", x"95", x"97", x"8f", x"85", x"83", x"8c", x"8f", x"85", x"7e", x"84", x"8a", x"8e", x"87", x"88", 
        x"ae", x"db", x"9b", x"80", x"8b", x"8e", x"87", x"7c", x"78", x"7b", x"7f", x"81", x"7e", x"7a", x"7e", 
        x"87", x"89", x"85", x"82", x"83", x"8b", x"8b", x"85", x"85", x"8b", x"8b", x"87", x"95", x"cf", x"bd", 
        x"7f", x"80", x"7a", x"76", x"78", x"7b", x"7b", x"7a", x"7b", x"7e", x"7e", x"7b", x"7e", x"84", x"83", 
        x"77", x"73", x"72", x"71", x"72", x"72", x"73", x"72", x"81", x"bf", x"b6", x"7e", x"7c", x"81", x"7e", 
        x"79", x"78", x"7c", x"79", x"74", x"77", x"7e", x"80", x"7c", x"79", x"72", x"6f", x"77", x"79", x"76", 
        x"75", x"75", x"84", x"c6", x"be", x"89", x"87", x"8f", x"87", x"80", x"85", x"88", x"88", x"93", x"9c", 
        x"9c", x"a1", x"a7", x"aa", x"af", x"b5", x"b3", x"a9", x"b1", x"bc", x"c1", x"d9", x"dd", x"d8", x"d2", 
        x"d0", x"cd", x"c9", x"c6", x"c6", x"c5", x"c4", x"ca", x"ce", x"cf", x"d2", x"d9", x"dd", x"da", x"de", 
        x"e3", x"e0", x"df", x"e8", x"e6", x"d5", x"dd", x"e5", x"e6", x"ea", x"ea", x"e5", x"df", x"d8", x"cf", 
        x"c3", x"bb", x"b1", x"ab", x"a8", x"9f", x"99", x"98", x"97", x"9d", x"a0", x"a1", x"a5", x"a6", x"a8", 
        x"a9", x"a8", x"a4", x"a1", x"a0", x"98", x"93", x"8b", x"82", x"79", x"72", x"6a", x"65", x"5e", x"55", 
        x"50", x"48", x"42", x"41", x"3d", x"3a", x"41", x"47", x"4d", x"5a", x"4b", x"1e", x"05", x"3d", x"62", 
        x"5c", x"57", x"56", x"54", x"57", x"54", x"54", x"54", x"55", x"5d", x"69", x"6f", x"77", x"82", x"8b", 
        x"77", x"68", x"72", x"74", x"6c", x"6e", x"6a", x"65", x"62", x"5b", x"53", x"4c", x"4c", x"26", x"08", 
        x"2a", x"57", x"5a", x"56", x"59", x"5a", x"5c", x"5e", x"5f", x"68", x"6f", x"68", x"5d", x"5b", x"59", 
        x"5b", x"58", x"57", x"54", x"52", x"54", x"56", x"55", x"50", x"47", x"46", x"4e", x"50", x"4e", x"4f", 
        x"48", x"4a", x"4d", x"4e", x"4e", x"41", x"60", x"86", x"89", x"88", x"7c", x"7c", x"78", x"74", x"6d", 
        x"6c", x"65", x"53", x"4f", x"4d", x"4e", x"4b", x"44", x"47", x"43", x"47", x"79", x"86", x"82", x"81", 
        x"84", x"81", x"81", x"83", x"83", x"79", x"57", x"54", x"52", x"55", x"47", x"1c", x"0a", x"04", x"05", 
        x"82", x"78", x"78", x"68", x"72", x"60", x"71", x"66", x"66", x"71", x"6c", x"5a", x"55", x"57", x"76", 
        x"59", x"5c", x"6d", x"49", x"41", x"36", x"3a", x"3b", x"40", x"3f", x"3c", x"30", x"37", x"45", x"32", 
        x"2e", x"52", x"75", x"80", x"60", x"38", x"45", x"3a", x"3b", x"4c", x"48", x"4a", x"57", x"4f", x"29", 
        x"34", x"5a", x"79", x"6b", x"55", x"45", x"5d", x"86", x"68", x"4f", x"3f", x"4e", x"3c", x"51", x"6f", 
        x"63", x"69", x"63", x"67", x"5d", x"5b", x"68", x"80", x"73", x"6a", x"61", x"77", x"81", x"6c", x"69", 
        x"6c", x"66", x"6c", x"79", x"8c", x"72", x"85", x"80", x"7d", x"91", x"96", x"91", x"7c", x"9e", x"c0", 
        x"b6", x"b0", x"c4", x"c1", x"ce", x"c8", x"d5", x"d6", x"cd", x"c0", x"b2", x"b2", x"ad", x"83", x"86", 
        x"a2", x"93", x"d8", x"df", x"de", x"de", x"dc", x"d9", x"cc", x"b7", x"a0", x"87", x"6d", x"53", x"3c", 
        x"2a", x"1f", x"1c", x"1d", x"25", x"35", x"45", x"45", x"48", x"4e", x"5c", x"66", x"6e", x"75", x"74", 
        x"6f", x"6b", x"69", x"6f", x"88", x"83", x"6f", x"6e", x"6f", x"6a", x"68", x"66", x"67", x"68", x"68", 
        x"69", x"62", x"66", x"b8", x"e4", x"d8", x"d7", x"d7", x"d5", x"df", x"d7", x"ce", x"d1", x"d0", x"d0", 
        x"cf", x"cf", x"ce", x"d0", x"d1", x"d0", x"d0", x"d0", x"d1", x"d0", x"d0", x"d1", x"d2", x"d3", x"d1", 
        x"d1", x"d2", x"d3", x"d2", x"d1", x"d2", x"d3", x"d4", x"d4", x"d3", x"d3", x"d2", x"d1", x"d2", x"d3", 
        x"d1", x"d1", x"d1", x"d2", x"d3", x"d2", x"d1", x"d2", x"d1", x"d1", x"d0", x"de", x"c5", x"91", x"7b", 
        x"76", x"74", x"71", x"76", x"83", x"af", x"9d", x"7f", x"77", x"76", x"7a", x"80", x"81", x"7b", x"76", 
        x"76", x"78", x"77", x"75", x"74", x"71", x"6d", x"6e", x"76", x"7a", x"7b", x"79", x"70", x"6e", x"75", 
        x"7f", x"7f", x"80", x"85", x"8a", x"8b", x"86", x"7e", x"7d", x"7d", x"7e", x"80", x"7f", x"73", x"70", 
        x"73", x"78", x"7a", x"80", x"bc", x"de", x"9d", x"81", x"7d", x"81", x"86", x"8b", x"86", x"7d", x"7b", 
        x"84", x"89", x"88", x"80", x"81", x"91", x"9a", x"9a", x"93", x"88", x"8e", x"98", x"96", x"8e", x"83", 
        x"82", x"8e", x"91", x"8c", x"7e", x"7a", x"80", x"87", x"86", x"7f", x"7d", x"85", x"8d", x"8c", x"94", 
        x"ce", x"d3", x"96", x"98", x"9a", x"9a", x"9b", x"9b", x"9b", x"98", x"92", x"93", x"96", x"97", x"93", 
        x"8c", x"85", x"87", x"87", x"80", x"7d", x"83", x"8c", x"92", x"92", x"8f", x"8c", x"8e", x"92", x"93", 
        x"95", x"95", x"96", x"9a", x"9b", x"96", x"8d", x"91", x"c4", x"d6", x"8a", x"7d", x"80", x"7c", x"75", 
        x"77", x"74", x"74", x"74", x"71", x"72", x"73", x"6f", x"70", x"77", x"7a", x"80", x"8b", x"91", x"9a", 
        x"94", x"9f", x"98", x"9c", x"9c", x"90", x"77", x"6e", x"6c", x"6f", x"73", x"6e", x"72", x"a9", x"db", 
        x"c1", x"bc", x"b6", x"b8", x"bd", x"bf", x"c1", x"bf", x"c3", x"c8", x"c6", x"bf", x"bb", x"c2", x"bf", 
        x"be", x"b8", x"bb", x"b9", x"b1", x"b1", x"b4", x"bd", x"c0", x"bf", x"c1", x"c2", x"c6", x"c5", x"c3", 
        x"c2", x"d3", x"bf", x"8f", x"8c", x"89", x"8b", x"8d", x"89", x"85", x"87", x"8b", x"87", x"7f", x"7d", 
        x"89", x"94", x"91", x"87", x"8c", x"92", x"97", x"90", x"86", x"85", x"8d", x"8d", x"8a", x"89", x"8e", 
        x"ac", x"d5", x"99", x"7a", x"7e", x"7f", x"7e", x"7f", x"80", x"7f", x"83", x"84", x"7e", x"7a", x"80", 
        x"89", x"8c", x"88", x"86", x"86", x"86", x"82", x"7c", x"7e", x"86", x"8b", x"87", x"93", x"ce", x"c6", 
        x"85", x"82", x"7c", x"79", x"7c", x"80", x"80", x"7d", x"7e", x"80", x"7c", x"77", x"79", x"7f", x"81", 
        x"78", x"76", x"76", x"74", x"73", x"74", x"75", x"75", x"84", x"c0", x"bc", x"82", x"7b", x"7d", x"7e", 
        x"80", x"80", x"7c", x"78", x"77", x"7e", x"87", x"89", x"82", x"7e", x"81", x"7e", x"7f", x"81", x"84", 
        x"84", x"80", x"89", x"c6", x"c5", x"94", x"89", x"91", x"92", x"86", x"83", x"8a", x"89", x"85", x"92", 
        x"95", x"87", x"88", x"92", x"91", x"86", x"86", x"8b", x"89", x"85", x"9f", x"e0", x"f3", x"f3", x"f4", 
        x"f2", x"f0", x"ee", x"eb", x"e9", x"e6", x"e3", x"e6", x"e5", x"e0", x"e0", x"e2", x"e2", x"da", x"dc", 
        x"dc", x"d3", x"d0", x"d5", x"d0", x"a2", x"86", x"8f", x"90", x"90", x"90", x"92", x"90", x"8e", x"8f", 
        x"8f", x"8f", x"8e", x"8e", x"92", x"93", x"94", x"98", x"98", x"97", x"90", x"8b", x"8c", x"85", x"7a", 
        x"71", x"6a", x"62", x"5c", x"52", x"4a", x"48", x"46", x"46", x"46", x"44", x"44", x"49", x"4c", x"4f", 
        x"55", x"58", x"5a", x"5b", x"5c", x"5d", x"60", x"60", x"5d", x"66", x"5f", x"29", x"04", x"41", x"65", 
        x"60", x"66", x"69", x"6a", x"6f", x"71", x"75", x"70", x"6a", x"79", x"9f", x"a1", x"9c", x"9a", x"96", 
        x"7d", x"5f", x"55", x"52", x"46", x"44", x"47", x"46", x"47", x"4a", x"4a", x"4d", x"51", x"2e", x"0b", 
        x"2b", x"5a", x"5f", x"5a", x"5c", x"5b", x"5c", x"5e", x"5e", x"65", x"6e", x"6a", x"5f", x"5c", x"59", 
        x"5b", x"58", x"57", x"53", x"51", x"53", x"54", x"50", x"48", x"48", x"4b", x"4f", x"51", x"51", x"51", 
        x"4a", x"4a", x"4d", x"4d", x"4c", x"41", x"5d", x"86", x"8b", x"89", x"7d", x"7d", x"7a", x"76", x"71", 
        x"6e", x"67", x"50", x"44", x"40", x"42", x"3f", x"3c", x"40", x"3f", x"41", x"73", x"85", x"81", x"81", 
        x"83", x"80", x"80", x"82", x"83", x"7c", x"5a", x"55", x"53", x"55", x"49", x"1e", x"09", x"07", x"19", 
        x"68", x"58", x"74", x"83", x"67", x"54", x"6b", x"5c", x"60", x"5e", x"6c", x"50", x"31", x"42", x"4c", 
        x"52", x"78", x"5a", x"2b", x"1f", x"2b", x"31", x"3f", x"40", x"3d", x"3c", x"4b", x"5c", x"46", x"24", 
        x"2e", x"58", x"66", x"57", x"4d", x"3f", x"2d", x"2f", x"2e", x"44", x"3c", x"35", x"41", x"42", x"2e", 
        x"33", x"3e", x"61", x"69", x"7b", x"83", x"83", x"63", x"65", x"66", x"37", x"44", x"5f", x"62", x"6b", 
        x"61", x"58", x"4c", x"53", x"61", x"52", x"56", x"67", x"60", x"50", x"51", x"6c", x"61", x"5c", x"60", 
        x"71", x"65", x"6a", x"73", x"8e", x"7f", x"89", x"98", x"a2", x"aa", x"b6", x"a4", x"7c", x"7e", x"92", 
        x"a4", x"a5", x"b1", x"9c", x"a3", x"ab", x"c0", x"9b", x"93", x"b7", x"af", x"a9", x"8f", x"98", x"88", 
        x"8c", x"94", x"d0", x"d0", x"c1", x"ae", x"92", x"76", x"5a", x"46", x"34", x"24", x"18", x"16", x"20", 
        x"2f", x"3f", x"4d", x"5a", x"66", x"6d", x"79", x"64", x"3d", x"54", x"6b", x"62", x"63", x"67", x"65", 
        x"66", x"66", x"66", x"69", x"84", x"84", x"6e", x"6b", x"6f", x"6c", x"69", x"67", x"68", x"69", x"6a", 
        x"6c", x"67", x"68", x"b6", x"e4", x"da", x"da", x"da", x"d5", x"de", x"d8", x"ce", x"d2", x"d0", x"d0", 
        x"cf", x"cf", x"cf", x"d0", x"d1", x"d1", x"d0", x"d0", x"d1", x"d1", x"d0", x"d1", x"d2", x"d3", x"d2", 
        x"d1", x"d2", x"d4", x"d3", x"d2", x"d2", x"d3", x"d4", x"d4", x"d3", x"d2", x"d2", x"d1", x"d0", x"d3", 
        x"d3", x"d1", x"d2", x"d3", x"d3", x"d3", x"d1", x"d3", x"d4", x"d4", x"cf", x"dd", x"cb", x"96", x"7d", 
        x"77", x"72", x"66", x"71", x"84", x"ac", x"9a", x"78", x"6b", x"6a", x"6f", x"71", x"6d", x"63", x"5f", 
        x"65", x"70", x"73", x"6c", x"66", x"67", x"6d", x"75", x"77", x"72", x"79", x"89", x"8f", x"89", x"83", 
        x"7b", x"78", x"83", x"8f", x"94", x"95", x"93", x"8a", x"80", x"7a", x"79", x"77", x"73", x"6e", x"72", 
        x"77", x"7a", x"79", x"7c", x"b5", x"e0", x"9d", x"82", x"84", x"8e", x"96", x"97", x"92", x"88", x"89", 
        x"91", x"92", x"90", x"86", x"86", x"8f", x"92", x"8e", x"84", x"7b", x"81", x"8c", x"8f", x"88", x"7c", 
        x"7b", x"85", x"85", x"82", x"7c", x"81", x"91", x"9c", x"9c", x"92", x"88", x"8a", x"91", x"96", x"9d", 
        x"cf", x"d3", x"99", x"98", x"97", x"90", x"8b", x"8a", x"8c", x"8b", x"88", x"89", x"8e", x"92", x"8f", 
        x"89", x"86", x"8d", x"94", x"96", x"94", x"95", x"97", x"9a", x"9d", x"9c", x"96", x"93", x"94", x"95", 
        x"95", x"90", x"8d", x"8d", x"8e", x"88", x"81", x"85", x"ba", x"d6", x"81", x"6f", x"78", x"79", x"72", 
        x"73", x"79", x"80", x"7f", x"7a", x"7d", x"85", x"88", x"84", x"87", x"90", x"96", x"99", x"94", x"9c", 
        x"92", x"9b", x"96", x"97", x"93", x"82", x"6d", x"67", x"64", x"69", x"6e", x"6a", x"6d", x"a2", x"d9", 
        x"c7", x"c2", x"c1", x"c4", x"c2", x"c1", x"c8", x"c5", x"c1", x"ba", x"b5", x"b4", x"b1", x"b1", x"b5", 
        x"bb", x"b7", x"b5", x"b7", x"b9", x"bd", x"be", x"c4", x"c8", x"c6", x"c6", x"c1", x"c5", x"c4", x"bf", 
        x"bc", x"ce", x"c2", x"87", x"82", x"82", x"83", x"81", x"7f", x"84", x"8d", x"90", x"87", x"86", x"90", 
        x"9c", x"9c", x"92", x"8c", x"93", x"95", x"91", x"88", x"84", x"85", x"85", x"7c", x"7b", x"85", x"8e", 
        x"a8", x"d4", x"9e", x"7e", x"84", x"87", x"85", x"83", x"86", x"87", x"82", x"7f", x"7d", x"7b", x"7d", 
        x"80", x"81", x"7f", x"7e", x"7c", x"7d", x"7d", x"7c", x"7c", x"82", x"87", x"82", x"8e", x"cb", x"c8", 
        x"82", x"7e", x"7c", x"7b", x"7d", x"7f", x"7c", x"79", x"79", x"7f", x"7c", x"7a", x"7d", x"85", x"86", 
        x"7f", x"7c", x"7a", x"76", x"75", x"76", x"79", x"7b", x"86", x"be", x"c0", x"83", x"7a", x"7a", x"7d", 
        x"80", x"81", x"7f", x"7b", x"77", x"7d", x"86", x"85", x"7c", x"7b", x"80", x"7e", x"7e", x"7f", x"7d", 
        x"82", x"82", x"88", x"bc", x"c8", x"9e", x"90", x"8f", x"92", x"8f", x"87", x"8c", x"95", x"90", x"8d", 
        x"95", x"93", x"89", x"89", x"90", x"89", x"80", x"83", x"86", x"7a", x"90", x"da", x"f3", x"f7", x"f4", 
        x"f2", x"f1", x"f2", x"f2", x"f2", x"f1", x"f1", x"f5", x"f5", x"f2", x"f2", x"f4", x"f4", x"f1", x"f1", 
        x"ee", x"e2", x"d8", x"cd", x"c1", x"8d", x"49", x"3e", x"3e", x"3c", x"3c", x"42", x"40", x"3f", x"44", 
        x"46", x"45", x"46", x"48", x"4e", x"51", x"50", x"4e", x"4c", x"47", x"3f", x"39", x"37", x"31", x"2b", 
        x"29", x"2a", x"2c", x"2d", x"2f", x"34", x"3d", x"46", x"4d", x"53", x"56", x"59", x"60", x"62", x"61", 
        x"63", x"63", x"63", x"62", x"64", x"68", x"6a", x"6e", x"6c", x"77", x"74", x"34", x"04", x"4e", x"7d", 
        x"76", x"77", x"73", x"70", x"73", x"72", x"72", x"5d", x"48", x"50", x"72", x"6e", x"65", x"61", x"5f", 
        x"58", x"4b", x"47", x"4a", x"46", x"48", x"50", x"51", x"54", x"56", x"55", x"5a", x"5d", x"34", x"04", 
        x"27", x"59", x"5f", x"5b", x"5d", x"5c", x"5c", x"5d", x"5d", x"61", x"69", x"6a", x"61", x"5c", x"58", 
        x"59", x"59", x"57", x"53", x"53", x"54", x"51", x"48", x"44", x"4b", x"4f", x"4f", x"51", x"53", x"52", 
        x"49", x"49", x"4f", x"4d", x"4a", x"3f", x"59", x"86", x"8d", x"8b", x"7e", x"7f", x"7d", x"78", x"75", 
        x"71", x"6a", x"51", x"3f", x"3b", x"3d", x"3c", x"3d", x"3e", x"3e", x"3f", x"72", x"85", x"80", x"80", 
        x"83", x"80", x"7f", x"80", x"82", x"7d", x"5c", x"56", x"55", x"56", x"4c", x"21", x"09", x"0b", x"32", 
        x"6b", x"67", x"75", x"7b", x"70", x"74", x"6e", x"5b", x"4e", x"63", x"82", x"5c", x"43", x"53", x"52", 
        x"52", x"61", x"43", x"32", x"47", x"34", x"33", x"34", x"35", x"3f", x"42", x"3f", x"5b", x"43", x"3a", 
        x"48", x"42", x"3a", x"41", x"49", x"3c", x"32", x"36", x"36", x"29", x"3b", x"48", x"3e", x"39", x"3f", 
        x"4f", x"58", x"66", x"63", x"59", x"7c", x"62", x"53", x"69", x"5c", x"45", x"4d", x"78", x"93", x"64", 
        x"42", x"63", x"87", x"90", x"8d", x"6b", x"5d", x"75", x"60", x"4b", x"51", x"50", x"42", x"61", x"5c", 
        x"51", x"59", x"7f", x"84", x"8e", x"95", x"86", x"8b", x"a4", x"b2", x"cc", x"d0", x"c3", x"ad", x"b5", 
        x"d1", x"de", x"d8", x"a2", x"b1", x"d2", x"ba", x"85", x"a8", x"be", x"89", x"8a", x"ae", x"95", x"64", 
        x"4e", x"6b", x"9b", x"7c", x"3b", x"2c", x"22", x"1c", x"1b", x"26", x"3b", x"4a", x"5d", x"6c", x"73", 
        x"76", x"7a", x"7b", x"7b", x"76", x"6c", x"75", x"61", x"2f", x"4b", x"6c", x"66", x"63", x"66", x"66", 
        x"65", x"67", x"66", x"6c", x"88", x"8e", x"7e", x"75", x"77", x"73", x"71", x"71", x"72", x"74", x"75", 
        x"76", x"71", x"6f", x"b6", x"e3", x"d9", x"d9", x"da", x"d6", x"de", x"d8", x"cd", x"d1", x"d0", x"d0", 
        x"d0", x"cf", x"cf", x"d0", x"d2", x"d1", x"d0", x"d0", x"d1", x"d2", x"d2", x"d2", x"d2", x"d3", x"d2", 
        x"d1", x"d2", x"d3", x"d2", x"d1", x"d2", x"d3", x"d5", x"d4", x"d3", x"d2", x"d2", x"d1", x"d1", x"d4", 
        x"d4", x"d2", x"d3", x"d4", x"d4", x"d4", x"d4", x"d6", x"d4", x"d1", x"ce", x"e1", x"d0", x"98", x"77", 
        x"6b", x"73", x"7a", x"83", x"8d", x"af", x"9e", x"84", x"86", x"8d", x"89", x"7f", x"7c", x"7a", x"7d", 
        x"7d", x"75", x"6a", x"64", x"66", x"68", x"6a", x"67", x"5f", x"5a", x"5e", x"68", x"7d", x"81", x"79", 
        x"65", x"65", x"75", x"7b", x"87", x"8c", x"8d", x"86", x"7f", x"80", x"87", x"7e", x"78", x"7d", x"82", 
        x"81", x"78", x"70", x"7f", x"bd", x"df", x"96", x"6d", x"71", x"7d", x"7b", x"78", x"74", x"75", x"83", 
        x"90", x"91", x"8d", x"89", x"8b", x"95", x"9a", x"9b", x"98", x"96", x"9a", x"9f", x"9d", x"93", x"88", 
        x"89", x"92", x"93", x"8f", x"82", x"7c", x"7e", x"80", x"7d", x"76", x"71", x"78", x"85", x"92", x"99", 
        x"ca", x"d3", x"97", x"92", x"92", x"95", x"99", x"a1", x"a8", x"a6", x"a1", x"98", x"97", x"9a", x"99", 
        x"96", x"8e", x"8b", x"8a", x"8a", x"87", x"81", x"7e", x"84", x"89", x"8b", x"8a", x"8b", x"90", x"93", 
        x"94", x"91", x"8f", x"95", x"9e", x"a3", x"a2", x"a0", x"c6", x"df", x"91", x"82", x"86", x"7d", x"74", 
        x"75", x"7b", x"7f", x"7b", x"71", x"6e", x"71", x"77", x"7c", x"83", x"8c", x"8e", x"91", x"8c", x"92", 
        x"8d", x"9a", x"97", x"99", x"97", x"91", x"7f", x"7b", x"7f", x"85", x"7e", x"71", x"74", x"a8", x"db", 
        x"c2", x"b2", x"ad", x"b8", x"be", x"bc", x"ba", x"ba", x"bf", x"b9", x"b4", x"b7", x"bb", x"c4", x"c0", 
        x"c4", x"c4", x"c0", x"be", x"be", x"c4", x"c3", x"c0", x"bd", x"ba", x"ba", x"b7", x"b9", x"b8", x"b8", 
        x"ba", x"ce", x"c4", x"89", x"8a", x"88", x"82", x"86", x"94", x"9b", x"94", x"8c", x"8e", x"93", x"95", 
        x"8e", x"87", x"82", x"82", x"89", x"86", x"82", x"87", x"8e", x"8d", x"85", x"80", x"88", x"97", x"9c", 
        x"b0", x"dc", x"a4", x"7f", x"85", x"88", x"82", x"7e", x"7e", x"7d", x"7b", x"7b", x"7e", x"84", x"8a", 
        x"8b", x"87", x"83", x"87", x"8c", x"89", x"82", x"7f", x"84", x"88", x"86", x"81", x"8c", x"c7", x"c9", 
        x"7f", x"7a", x"77", x"77", x"7a", x"7c", x"7a", x"7b", x"80", x"88", x"85", x"7e", x"7e", x"85", x"82", 
        x"7d", x"7f", x"7c", x"76", x"70", x"6e", x"6e", x"6f", x"7c", x"b6", x"c3", x"89", x"80", x"7f", x"7e", 
        x"7c", x"7e", x"85", x"86", x"7c", x"7c", x"82", x"7f", x"7b", x"79", x"7b", x"79", x"7d", x"7f", x"7f", 
        x"7c", x"79", x"7d", x"b3", x"c9", x"a1", x"95", x"8e", x"8e", x"97", x"95", x"8b", x"91", x"99", x"8f", 
        x"88", x"8e", x"8f", x"84", x"80", x"89", x"86", x"7a", x"85", x"89", x"99", x"da", x"f3", x"f3", x"f4", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f1", x"ef", x"f2", x"f4", x"f4", x"f4", x"f4", x"f5", x"f6", x"f4", 
        x"f1", x"e2", x"cf", x"b8", x"b3", x"af", x"78", x"56", x"4f", x"40", x"33", x"32", x"2e", x"2c", x"27", 
        x"22", x"1e", x"20", x"24", x"28", x"2a", x"1b", x"0a", x"08", x"0d", x"19", x"21", x"24", x"23", x"24", 
        x"27", x"2b", x"2f", x"31", x"32", x"2f", x"34", x"43", x"4f", x"4d", x"4e", x"52", x"5e", x"62", x"62", 
        x"65", x"68", x"6b", x"6d", x"6d", x"6d", x"6c", x"71", x"70", x"74", x"75", x"3a", x"06", x"48", x"6f", 
        x"66", x"68", x"68", x"65", x"67", x"66", x"69", x"55", x"3d", x"3e", x"3b", x"3c", x"42", x"49", x"4d", 
        x"51", x"54", x"50", x"4e", x"4f", x"4d", x"50", x"51", x"55", x"58", x"56", x"5a", x"5a", x"37", x"04", 
        x"23", x"55", x"5d", x"5b", x"5c", x"5a", x"59", x"5b", x"5b", x"5e", x"67", x"6d", x"65", x"5b", x"57", 
        x"59", x"59", x"55", x"53", x"54", x"53", x"4b", x"43", x"48", x"4c", x"4f", x"50", x"50", x"51", x"52", 
        x"4a", x"49", x"51", x"4d", x"48", x"3c", x"55", x"85", x"8e", x"8d", x"82", x"83", x"80", x"79", x"77", 
        x"72", x"6d", x"53", x"40", x"3e", x"41", x"40", x"40", x"3e", x"3d", x"3e", x"71", x"85", x"7d", x"7f", 
        x"82", x"81", x"80", x"7e", x"80", x"7d", x"5b", x"53", x"55", x"57", x"51", x"26", x"0a", x"08", x"34", 
        x"7f", x"7c", x"74", x"6f", x"6e", x"6f", x"54", x"66", x"82", x"6b", x"4a", x"4c", x"4d", x"3e", x"4c", 
        x"2a", x"38", x"48", x"2a", x"2e", x"32", x"2c", x"24", x"2c", x"3e", x"5c", x"3f", x"5d", x"5b", x"3f", 
        x"56", x"51", x"55", x"62", x"73", x"46", x"2c", x"34", x"4b", x"4f", x"4f", x"34", x"35", x"4c", x"4a", 
        x"46", x"54", x"63", x"65", x"44", x"3a", x"44", x"5d", x"84", x"7d", x"59", x"64", x"75", x"67", x"51", 
        x"55", x"55", x"7f", x"8f", x"80", x"70", x"5b", x"52", x"4b", x"57", x"5c", x"57", x"51", x"4d", x"5d", 
        x"5b", x"8a", x"69", x"4f", x"64", x"99", x"7c", x"62", x"72", x"77", x"8c", x"8d", x"87", x"8d", x"98", 
        x"b4", x"c8", x"c1", x"af", x"d1", x"ee", x"d7", x"b6", x"d3", x"d4", x"b7", x"b5", x"c5", x"bf", x"7d", 
        x"4b", x"aa", x"c5", x"80", x"1d", x"2e", x"3d", x"41", x"49", x"52", x"5d", x"60", x"65", x"68", x"64", 
        x"62", x"66", x"67", x"66", x"67", x"66", x"6d", x"5f", x"34", x"4d", x"71", x"70", x"65", x"65", x"69", 
        x"69", x"6a", x"67", x"6e", x"86", x"92", x"8c", x"7f", x"80", x"7b", x"7b", x"7b", x"7d", x"7d", x"7d", 
        x"7d", x"76", x"71", x"b5", x"e2", x"d8", x"d8", x"d9", x"d7", x"df", x"d8", x"cc", x"d0", x"cf", x"d0", 
        x"d0", x"cf", x"cf", x"d0", x"d2", x"d1", x"d0", x"d0", x"d1", x"d4", x"d5", x"d4", x"d3", x"d3", x"d2", 
        x"d1", x"d2", x"d2", x"d1", x"d1", x"d2", x"d4", x"d5", x"d4", x"d3", x"d2", x"d2", x"d1", x"d2", x"d5", 
        x"d3", x"d2", x"d2", x"d3", x"d4", x"d4", x"d3", x"d4", x"d1", x"d0", x"cf", x"e2", x"cf", x"9c", x"87", 
        x"7b", x"76", x"65", x"60", x"76", x"ac", x"9c", x"76", x"69", x"68", x"66", x"69", x"73", x"77", x"79", 
        x"79", x"75", x"71", x"74", x"7b", x"7e", x"7d", x"7b", x"7a", x"84", x"87", x"88", x"8b", x"84", x"7f", 
        x"7b", x"83", x"8d", x"86", x"78", x"78", x"7c", x"76", x"70", x"70", x"6c", x"64", x"62", x"65", x"6b", 
        x"71", x"6c", x"62", x"6f", x"ac", x"dd", x"a1", x"85", x"93", x"9b", x"9a", x"92", x"88", x"89", x"90", 
        x"91", x"8a", x"81", x"82", x"87", x"8e", x"8b", x"81", x"75", x"72", x"7b", x"80", x"7f", x"7b", x"78", 
        x"83", x"8e", x"8f", x"8d", x"83", x"84", x"8d", x"97", x"98", x"93", x"8a", x"8c", x"93", x"99", x"9c", 
        x"cd", x"d9", x"99", x"96", x"9b", x"9b", x"94", x"8f", x"8f", x"8e", x"8e", x"89", x"8c", x"92", x"92", 
        x"92", x"8f", x"8a", x"89", x"8e", x"91", x"90", x"91", x"9c", x"a1", x"a2", x"a0", x"9a", x"96", x"95", 
        x"99", x"9b", x"99", x"96", x"94", x"91", x"8d", x"8f", x"bd", x"dc", x"85", x"69", x"6c", x"70", x"73", 
        x"70", x"71", x"75", x"78", x"77", x"78", x"7c", x"85", x"90", x"95", x"97", x"94", x"98", x"96", x"9b", 
        x"94", x"9d", x"99", x"9b", x"93", x"8a", x"73", x"66", x"65", x"6f", x"72", x"6b", x"6b", x"a2", x"db", 
        x"c6", x"bb", x"b7", x"bb", x"c1", x"c8", x"c5", x"bc", x"bd", x"bc", x"be", x"c1", x"be", x"c1", x"be", 
        x"bc", x"b8", x"b7", x"bc", x"bc", x"bc", x"be", x"ba", x"ba", x"ba", x"ba", x"b9", x"bd", x"c4", x"c3", 
        x"bd", x"cf", x"cc", x"8f", x"89", x"85", x"88", x"90", x"92", x"8a", x"84", x"83", x"8a", x"8e", x"8a", 
        x"86", x"8a", x"8e", x"8d", x"8a", x"8a", x"90", x"97", x"95", x"8c", x"84", x"86", x"90", x"97", x"91", 
        x"a5", x"db", x"a0", x"75", x"7c", x"82", x"80", x"80", x"81", x"7f", x"80", x"83", x"85", x"85", x"83", 
        x"82", x"83", x"84", x"85", x"86", x"7f", x"79", x"7a", x"7f", x"81", x"7f", x"7e", x"8a", x"c5", x"d0", 
        x"88", x"83", x"7f", x"81", x"85", x"85", x"80", x"80", x"84", x"8a", x"89", x"84", x"86", x"8f", x"86", 
        x"7f", x"7a", x"76", x"72", x"6f", x"6f", x"71", x"72", x"7d", x"b4", x"c5", x"84", x"79", x"79", x"7c", 
        x"7f", x"80", x"7f", x"80", x"7a", x"7b", x"80", x"7e", x"7f", x"7b", x"7b", x"7c", x"7b", x"7e", x"87", 
        x"81", x"7e", x"81", x"b5", x"c9", x"9d", x"97", x"95", x"90", x"96", x"9b", x"92", x"8a", x"95", x"9b", 
        x"93", x"8b", x"91", x"94", x"87", x"84", x"89", x"85", x"83", x"86", x"99", x"d8", x"f5", x"f1", x"f2", 
        x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f5", x"f4", x"f3", x"f6", x"f2", x"f2", 
        x"f6", x"e9", x"d4", x"b5", x"ad", x"b3", x"97", x"69", x"59", x"52", x"48", x"42", x"3d", x"3a", x"34", 
        x"2e", x"26", x"26", x"27", x"21", x"1c", x"10", x"02", x"03", x"06", x"0e", x"13", x"14", x"15", x"16", 
        x"17", x"18", x"1c", x"1d", x"1c", x"19", x"27", x"4c", x"61", x"5b", x"62", x"64", x"6c", x"69", x"5e", 
        x"54", x"4f", x"4e", x"4b", x"49", x"4b", x"47", x"4a", x"49", x"4a", x"54", x"2f", x"06", x"3c", x"63", 
        x"64", x"69", x"6b", x"6d", x"6d", x"6a", x"6f", x"5c", x"42", x"42", x"40", x"42", x"48", x"4e", x"52", 
        x"53", x"57", x"59", x"50", x"52", x"50", x"51", x"53", x"55", x"55", x"56", x"5c", x"5a", x"3b", x"07", 
        x"1f", x"50", x"5d", x"5a", x"5b", x"59", x"5a", x"5e", x"5f", x"5b", x"60", x"6c", x"69", x"5e", x"57", 
        x"58", x"57", x"55", x"53", x"51", x"4b", x"45", x"45", x"4c", x"4f", x"50", x"50", x"50", x"4f", x"4f", 
        x"48", x"45", x"4c", x"48", x"44", x"39", x"4e", x"83", x"8f", x"8e", x"84", x"86", x"82", x"7a", x"78", 
        x"74", x"6e", x"55", x"40", x"40", x"42", x"3f", x"3e", x"3e", x"3e", x"3b", x"6c", x"83", x"7d", x"7d", 
        x"81", x"81", x"81", x"7e", x"80", x"7f", x"5d", x"53", x"54", x"56", x"53", x"29", x"0c", x"08", x"32", 
        x"51", x"43", x"53", x"53", x"62", x"78", x"6a", x"7b", x"6f", x"42", x"35", x"66", x"71", x"62", x"51", 
        x"35", x"3d", x"3c", x"3a", x"25", x"37", x"33", x"2c", x"2d", x"61", x"6e", x"34", x"34", x"56", x"5c", 
        x"60", x"67", x"5f", x"51", x"79", x"75", x"60", x"41", x"36", x"50", x"68", x"3a", x"40", x"4e", x"3d", 
        x"40", x"55", x"58", x"5c", x"4f", x"5c", x"60", x"69", x"6e", x"4e", x"35", x"57", x"7c", x"6f", x"69", 
        x"78", x"76", x"88", x"72", x"2d", x"4f", x"50", x"27", x"20", x"40", x"41", x"39", x"4d", x"5c", x"40", 
        x"41", x"56", x"58", x"50", x"41", x"71", x"7c", x"6b", x"69", x"6c", x"74", x"64", x"48", x"5f", x"4d", 
        x"53", x"63", x"64", x"5c", x"82", x"ad", x"d5", x"bc", x"b7", x"c0", x"c6", x"c8", x"b6", x"c5", x"a6", 
        x"77", x"e5", x"e2", x"8a", x"48", x"93", x"b4", x"aa", x"a4", x"98", x"9c", x"9f", x"95", x"85", x"81", 
        x"81", x"79", x"6d", x"6a", x"6d", x"70", x"72", x"60", x"31", x"49", x"6f", x"75", x"6d", x"6d", x"6e", 
        x"69", x"6c", x"6a", x"73", x"89", x"97", x"97", x"84", x"83", x"7c", x"7c", x"7d", x"7e", x"7c", x"79", 
        x"76", x"6b", x"68", x"ad", x"df", x"d8", x"d9", x"db", x"d8", x"df", x"d8", x"cb", x"cf", x"cf", x"d0", 
        x"d0", x"cf", x"d0", x"d1", x"d2", x"d1", x"d1", x"d0", x"d1", x"d4", x"d6", x"d5", x"d4", x"d3", x"d3", 
        x"d2", x"d3", x"d2", x"d1", x"d1", x"d3", x"d4", x"d4", x"d3", x"d3", x"d2", x"d2", x"d1", x"d2", x"d4", 
        x"d2", x"d1", x"d2", x"d3", x"d3", x"d3", x"d4", x"d2", x"d0", x"d1", x"cf", x"e0", x"d2", x"9d", x"7d", 
        x"72", x"7d", x"7d", x"81", x"8a", x"a3", x"9c", x"8f", x"87", x"82", x"83", x"88", x"8f", x"8b", x"7d", 
        x"79", x"7e", x"83", x"81", x"7c", x"6f", x"64", x"62", x"63", x"6b", x"67", x"63", x"67", x"5f", x"65", 
        x"6f", x"73", x"80", x"8b", x"7a", x"75", x"7c", x"81", x"82", x"85", x"82", x"7f", x"85", x"8f", x"94", 
        x"95", x"8a", x"7c", x"86", x"b8", x"df", x"9c", x"75", x"7f", x"83", x"79", x"6c", x"6a", x"75", x"80", 
        x"7e", x"7a", x"77", x"86", x"8c", x"8f", x"8c", x"8c", x"92", x"a0", x"aa", x"a9", x"a2", x"98", x"90", 
        x"94", x"97", x"94", x"8e", x"83", x"83", x"8c", x"8f", x"87", x"76", x"67", x"6a", x"70", x"7a", x"87", 
        x"c3", x"d5", x"92", x"90", x"95", x"94", x"8f", x"8f", x"97", x"a2", x"a5", x"9f", x"9d", x"9f", x"9d", 
        x"9c", x"94", x"8f", x"8f", x"93", x"96", x"94", x"93", x"8d", x"89", x"87", x"88", x"88", x"87", x"89", 
        x"8d", x"90", x"90", x"8e", x"8f", x"92", x"94", x"97", x"bf", x"da", x"8c", x"7b", x"80", x"82", x"89", 
        x"8a", x"86", x"83", x"80", x"7a", x"77", x"7a", x"87", x"8d", x"8b", x"89", x"86", x"8c", x"8a", x"90", 
        x"8b", x"93", x"8c", x"8e", x"89", x"85", x"76", x"6f", x"70", x"76", x"7c", x"7b", x"79", x"a6", x"dc", 
        x"c3", x"b8", x"bc", x"c1", x"bb", x"ba", x"be", x"b9", x"b8", x"b2", x"b9", x"c3", x"c0", x"bc", x"b9", 
        x"bb", x"bf", x"bd", x"be", x"bf", x"c5", x"c9", x"bf", x"b9", x"b9", x"bc", x"c2", x"bf", x"c3", x"c0", 
        x"ba", x"ca", x"c2", x"84", x"81", x"7c", x"7e", x"87", x"89", x"80", x"7d", x"83", x"8d", x"8d", x"88", 
        x"8d", x"97", x"96", x"8d", x"89", x"8a", x"93", x"92", x"83", x"78", x"7d", x"82", x"8c", x"8e", x"86", 
        x"9d", x"dc", x"a1", x"75", x"7b", x"81", x"82", x"85", x"85", x"80", x"80", x"82", x"81", x"7f", x"7c", 
        x"7c", x"7d", x"7d", x"7c", x"7d", x"7a", x"79", x"7c", x"80", x"81", x"82", x"85", x"8b", x"c0", x"cf", 
        x"87", x"80", x"80", x"86", x"8c", x"8b", x"82", x"7e", x"81", x"84", x"8b", x"8c", x"93", x"9c", x"8a", 
        x"7e", x"7c", x"79", x"76", x"74", x"72", x"70", x"6e", x"78", x"b1", x"cb", x"8a", x"7b", x"78", x"78", 
        x"79", x"77", x"78", x"80", x"7d", x"7a", x"7a", x"76", x"78", x"78", x"78", x"7a", x"7e", x"7c", x"82", 
        x"7d", x"7b", x"7d", x"b5", x"cf", x"9f", x"90", x"97", x"92", x"86", x"8d", x"98", x"91", x"8c", x"95", 
        x"97", x"8b", x"89", x"94", x"8d", x"82", x"89", x"93", x"8e", x"84", x"92", x"d0", x"f1", x"f3", x"f2", 
        x"f2", x"f1", x"ef", x"f0", x"f3", x"f6", x"f7", x"f4", x"f4", x"f5", x"f2", x"f0", x"f3", x"f2", x"ef", 
        x"f1", x"e6", x"d6", x"b6", x"aa", x"ac", x"b2", x"84", x"63", x"54", x"4a", x"42", x"3a", x"36", x"37", 
        x"35", x"2a", x"25", x"22", x"1c", x"1b", x"13", x"06", x"05", x"03", x"04", x"04", x"05", x"06", x"06", 
        x"05", x"04", x"06", x"08", x"08", x"0b", x"1e", x"40", x"48", x"40", x"58", x"63", x"71", x"73", x"6d", 
        x"65", x"62", x"61", x"5f", x"5e", x"62", x"57", x"50", x"4d", x"50", x"59", x"35", x"07", x"2d", x"49", 
        x"45", x"48", x"4e", x"56", x"5a", x"5b", x"67", x"5a", x"40", x"40", x"45", x"46", x"49", x"4d", x"54", 
        x"53", x"54", x"5b", x"4d", x"51", x"52", x"53", x"56", x"55", x"55", x"54", x"58", x"59", x"3f", x"0a", 
        x"1b", x"4e", x"60", x"5a", x"59", x"57", x"58", x"5d", x"5e", x"57", x"57", x"65", x"6b", x"61", x"57", 
        x"55", x"57", x"54", x"54", x"4d", x"44", x"43", x"4b", x"4e", x"51", x"50", x"4e", x"4f", x"50", x"4b", 
        x"48", x"44", x"49", x"44", x"41", x"38", x"4b", x"82", x"91", x"8f", x"84", x"86", x"83", x"7d", x"7b", 
        x"76", x"70", x"57", x"41", x"42", x"44", x"41", x"42", x"43", x"44", x"3c", x"69", x"83", x"7e", x"7c", 
        x"80", x"80", x"81", x"7f", x"81", x"80", x"61", x"55", x"55", x"55", x"52", x"2a", x"0c", x"06", x"2d", 
        x"6e", x"4c", x"64", x"64", x"71", x"6b", x"6f", x"55", x"40", x"4c", x"42", x"50", x"46", x"46", x"3c", 
        x"49", x"4a", x"42", x"4f", x"42", x"45", x"4c", x"39", x"33", x"62", x"62", x"30", x"39", x"47", x"57", 
        x"51", x"5a", x"77", x"7b", x"69", x"3a", x"40", x"3e", x"36", x"3c", x"3f", x"2f", x"3d", x"34", x"21", 
        x"3f", x"79", x"6f", x"4e", x"44", x"6a", x"70", x"61", x"46", x"27", x"21", x"2e", x"63", x"6f", x"5b", 
        x"69", x"82", x"7a", x"5c", x"29", x"33", x"36", x"23", x"1a", x"2c", x"3b", x"3a", x"4d", x"62", x"40", 
        x"4e", x"59", x"61", x"4d", x"46", x"55", x"80", x"85", x"77", x"76", x"71", x"46", x"3e", x"69", x"5e", 
        x"41", x"5d", x"69", x"41", x"4e", x"73", x"bd", x"84", x"3b", x"55", x"5b", x"59", x"5c", x"6b", x"64", 
        x"5f", x"ac", x"c1", x"95", x"55", x"a7", x"c4", x"c9", x"cf", x"bd", x"b0", x"c7", x"c3", x"a3", x"ae", 
        x"d2", x"c6", x"b7", x"c2", x"bd", x"95", x"79", x"5d", x"2e", x"46", x"6a", x"74", x"6e", x"70", x"75", 
        x"72", x"74", x"74", x"7c", x"93", x"98", x"9c", x"8b", x"87", x"7b", x"75", x"75", x"73", x"72", x"72", 
        x"71", x"6a", x"69", x"ab", x"e0", x"db", x"d9", x"d8", x"d5", x"dc", x"da", x"ca", x"cf", x"ce", x"d0", 
        x"ce", x"ce", x"d1", x"d1", x"d1", x"d1", x"d2", x"d3", x"d0", x"d0", x"d2", x"d4", x"d3", x"d2", x"d3", 
        x"d3", x"d4", x"d3", x"d1", x"d0", x"d3", x"d5", x"d4", x"d2", x"d0", x"d0", x"d0", x"d1", x"d2", x"d3", 
        x"d3", x"d3", x"d4", x"d5", x"d5", x"d5", x"d4", x"d2", x"d2", x"d2", x"d0", x"df", x"ce", x"92", x"81", 
        x"74", x"6a", x"5a", x"5f", x"76", x"ab", x"9f", x"76", x"66", x"64", x"6c", x"6c", x"6b", x"67", x"60", 
        x"64", x"70", x"7b", x"7c", x"80", x"7d", x"77", x"7c", x"83", x"8a", x"90", x"8e", x"87", x"8a", x"8f", 
        x"8c", x"85", x"81", x"78", x"79", x"7d", x"7f", x"7a", x"71", x"6a", x"68", x"69", x"6c", x"68", x"61", 
        x"5e", x"60", x"60", x"6b", x"a7", x"de", x"a1", x"81", x"8e", x"90", x"8e", x"8b", x"8e", x"9a", x"a1", 
        x"98", x"8b", x"86", x"8f", x"97", x"9a", x"8d", x"80", x"7b", x"80", x"84", x"81", x"77", x"70", x"76", 
        x"83", x"87", x"88", x"84", x"7e", x"82", x"8c", x"8f", x"8c", x"88", x"87", x"94", x"a3", x"a5", x"a9", 
        x"cb", x"d7", x"9d", x"98", x"9b", x"99", x"97", x"91", x"90", x"91", x"8e", x"8b", x"83", x"7d", x"7f", 
        x"83", x"83", x"85", x"87", x"8a", x"8e", x"8f", x"8e", x"8a", x"8e", x"95", x"9d", x"a2", x"9d", x"95", 
        x"95", x"99", x"9a", x"98", x"93", x"90", x"91", x"97", x"be", x"de", x"8d", x"79", x"78", x"6f", x"6b", 
        x"6e", x"6f", x"6d", x"69", x"70", x"80", x"8d", x"8b", x"8e", x"91", x"8f", x"90", x"97", x"97", x"9e", 
        x"9a", x"9f", x"95", x"9a", x"9b", x"8c", x"78", x"76", x"74", x"68", x"65", x"67", x"6b", x"a0", x"dd", 
        x"c3", x"b6", x"b9", x"bf", x"bf", x"bd", x"bc", x"ba", x"c2", x"c7", x"c5", x"c4", x"c1", x"c0", x"bd", 
        x"b8", x"b8", x"ba", x"bd", x"be", x"b5", x"ba", x"ba", x"ba", x"bc", x"bc", x"c0", x"c2", x"c2", x"bf", 
        x"b9", x"c9", x"c5", x"87", x"84", x"8c", x"94", x"8f", x"88", x"8a", x"8c", x"8a", x"84", x"85", x"8a", 
        x"8d", x"89", x"84", x"82", x"84", x"86", x"8a", x"8b", x"82", x"79", x"7e", x"89", x"8b", x"88", x"85", 
        x"9a", x"d9", x"a7", x"7c", x"7e", x"7f", x"81", x"80", x"7a", x"78", x"79", x"7b", x"7d", x"7a", x"7a", 
        x"7e", x"7e", x"7f", x"7d", x"7c", x"80", x"80", x"86", x"8b", x"88", x"87", x"87", x"8d", x"bb", x"d4", 
        x"87", x"7d", x"7c", x"7d", x"85", x"87", x"82", x"7e", x"82", x"86", x"8e", x"9a", x"99", x"a0", x"8e", 
        x"7f", x"7b", x"79", x"76", x"78", x"79", x"71", x"6e", x"79", x"b0", x"ce", x"87", x"79", x"79", x"7b", 
        x"7d", x"7c", x"7a", x"7a", x"78", x"7a", x"7f", x"7b", x"7a", x"7a", x"7a", x"7e", x"7d", x"78", x"7a", 
        x"80", x"7f", x"81", x"b2", x"cd", x"a2", x"88", x"91", x"99", x"92", x"88", x"91", x"9b", x"95", x"8f", 
        x"94", x"95", x"8a", x"86", x"8c", x"89", x"7f", x"80", x"8d", x"8e", x"93", x"ce", x"f4", x"f5", x"f4", 
        x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f5", x"f5", x"f4", x"f5", x"f3", x"f2", x"f2", x"f2", x"f1", 
        x"f2", x"e9", x"d7", x"bb", x"b3", x"b4", x"b5", x"a0", x"73", x"62", x"5e", x"54", x"51", x"4a", x"40", 
        x"35", x"2d", x"2b", x"2c", x"27", x"1f", x"14", x"05", x"03", x"04", x"06", x"07", x"07", x"08", x"04", 
        x"06", x"04", x"05", x"05", x"05", x"0c", x"28", x"41", x"3e", x"39", x"4f", x"58", x"69", x"72", x"6d", 
        x"69", x"6a", x"6c", x"6c", x"6c", x"6d", x"6e", x"6c", x"6b", x"6e", x"71", x"42", x"0a", x"2a", x"4f", 
        x"52", x"54", x"56", x"55", x"51", x"4e", x"50", x"47", x"32", x"2e", x"2f", x"31", x"34", x"3a", x"49", 
        x"4f", x"55", x"62", x"58", x"54", x"58", x"5c", x"60", x"5e", x"5c", x"5a", x"5c", x"60", x"43", x"0f", 
        x"19", x"4b", x"5b", x"56", x"5a", x"58", x"5a", x"5e", x"5a", x"59", x"5b", x"5e", x"6a", x"64", x"54", 
        x"57", x"5a", x"55", x"52", x"46", x"44", x"4c", x"4e", x"4e", x"4e", x"4e", x"4f", x"50", x"50", x"4e", 
        x"4d", x"43", x"48", x"46", x"42", x"3a", x"48", x"7f", x"93", x"91", x"87", x"8b", x"84", x"7e", x"7d", 
        x"77", x"70", x"59", x"40", x"3f", x"3f", x"3e", x"3e", x"3d", x"3d", x"3a", x"63", x"7e", x"7e", x"7f", 
        x"80", x"7d", x"7d", x"7f", x"80", x"80", x"61", x"53", x"53", x"52", x"51", x"2d", x"0c", x"09", x"2a", 
        x"46", x"74", x"89", x"74", x"55", x"4e", x"64", x"64", x"5a", x"5a", x"6f", x"5b", x"32", x"26", x"2f", 
        x"48", x"42", x"3d", x"2a", x"23", x"2c", x"32", x"2b", x"53", x"91", x"6c", x"52", x"4a", x"4c", x"55", 
        x"69", x"56", x"53", x"76", x"6b", x"32", x"2d", x"3f", x"58", x"33", x"25", x"40", x"47", x"3b", x"2f", 
        x"6a", x"7e", x"47", x"52", x"54", x"3c", x"39", x"75", x"66", x"35", x"2c", x"37", x"4a", x"67", x"51", 
        x"6a", x"5a", x"53", x"61", x"2e", x"2e", x"3e", x"31", x"2c", x"2e", x"34", x"4f", x"37", x"4f", x"67", 
        x"6e", x"56", x"36", x"3a", x"62", x"5f", x"7e", x"8c", x"7a", x"79", x"72", x"53", x"39", x"66", x"7f", 
        x"47", x"61", x"6a", x"73", x"9f", x"7a", x"c2", x"8e", x"2c", x"55", x"50", x"2b", x"47", x"3b", x"33", 
        x"54", x"72", x"74", x"61", x"50", x"8e", x"92", x"93", x"a1", x"a5", x"a4", x"af", x"b6", x"a1", x"a5", 
        x"c2", x"be", x"bd", x"b3", x"b1", x"9f", x"90", x"7c", x"36", x"49", x"71", x"74", x"6f", x"7b", x"7c", 
        x"7c", x"7f", x"7b", x"80", x"96", x"98", x"93", x"84", x"82", x"75", x"72", x"75", x"74", x"72", x"72", 
        x"72", x"68", x"65", x"a8", x"e1", x"d9", x"d7", x"d9", x"d3", x"da", x"d9", x"ca", x"cf", x"cf", x"d0", 
        x"ce", x"cf", x"d1", x"d1", x"d1", x"d1", x"d2", x"d4", x"d0", x"d0", x"d1", x"d2", x"d2", x"d0", x"d2", 
        x"d3", x"d4", x"d3", x"d1", x"d1", x"d3", x"d5", x"d5", x"d3", x"d2", x"d1", x"d1", x"d0", x"cf", x"d2", 
        x"d3", x"d3", x"d4", x"d5", x"d5", x"d5", x"d5", x"d2", x"d1", x"d1", x"d0", x"e2", x"d9", x"a6", x"84", 
        x"77", x"80", x"79", x"84", x"87", x"9d", x"95", x"81", x"8d", x"93", x"97", x"94", x"8d", x"86", x"89", 
        x"8d", x"8f", x"8b", x"80", x"7f", x"7a", x"78", x"7d", x"78", x"6b", x"68", x"69", x"6b", x"72", x"76", 
        x"6d", x"62", x"61", x"62", x"6d", x"73", x"76", x"73", x"6f", x"71", x"79", x"83", x"8b", x"8c", x"87", 
        x"82", x"83", x"85", x"88", x"b4", x"e5", x"ab", x"8c", x"93", x"8b", x"7e", x"70", x"72", x"78", x"7e", 
        x"76", x"6b", x"6c", x"7b", x"83", x"85", x"7e", x"7a", x"7f", x"8b", x"90", x"92", x"8f", x"8c", x"92", 
        x"9e", x"a3", x"a1", x"95", x"88", x"88", x"90", x"99", x"9d", x"95", x"81", x"79", x"76", x"75", x"87", 
        x"c0", x"d6", x"88", x"83", x"8b", x"8d", x"8f", x"8b", x"8a", x"90", x"91", x"93", x"93", x"94", x"9c", 
        x"a5", x"a8", x"a4", x"99", x"91", x"94", x"99", x"98", x"96", x"92", x"8f", x"8d", x"8e", x"8b", x"86", 
        x"83", x"81", x"81", x"86", x"89", x"89", x"8a", x"8b", x"b1", x"de", x"8e", x"76", x"7b", x"7a", x"77", 
        x"7a", x"85", x"88", x"89", x"94", x"9b", x"9b", x"92", x"93", x"95", x"94", x"90", x"91", x"8c", x"92", 
        x"8e", x"92", x"88", x"8b", x"89", x"7a", x"61", x"65", x"70", x"70", x"70", x"6d", x"69", x"98", x"d8", 
        x"cf", x"c5", x"c3", x"c0", x"bc", x"be", x"c3", x"be", x"bc", x"b9", x"b9", x"bb", x"b8", x"b0", x"b4", 
        x"b9", x"bd", x"bc", x"ba", x"c0", x"bd", x"bc", x"ba", x"bc", x"c8", x"cd", x"c7", x"c4", x"c3", x"bf", 
        x"ba", x"cc", x"cc", x"90", x"8e", x"8b", x"82", x"81", x"89", x"8c", x"83", x"7c", x"7f", x"82", x"8a", 
        x"90", x"8c", x"86", x"88", x"96", x"9b", x"96", x"8d", x"84", x"83", x"8b", x"85", x"83", x"85", x"88", 
        x"99", x"d5", x"ab", x"79", x"77", x"7a", x"80", x"83", x"80", x"80", x"80", x"80", x"83", x"7f", x"80", 
        x"85", x"85", x"85", x"81", x"82", x"85", x"82", x"86", x"88", x"84", x"84", x"82", x"86", x"b5", x"d5", 
        x"88", x"7f", x"7d", x"80", x"85", x"88", x"81", x"84", x"8b", x"93", x"97", x"a0", x"9b", x"a4", x"95", 
        x"87", x"7d", x"77", x"72", x"72", x"74", x"6f", x"6e", x"79", x"ad", x"cc", x"85", x"79", x"7b", x"7a", 
        x"7d", x"80", x"7f", x"7d", x"79", x"7a", x"80", x"7b", x"79", x"78", x"79", x"80", x"83", x"81", x"81", 
        x"7c", x"78", x"7a", x"a9", x"cc", x"a6", x"8e", x"89", x"8e", x"94", x"91", x"8e", x"92", x"9e", x"9a", 
        x"91", x"93", x"92", x"85", x"7f", x"8b", x"8f", x"85", x"83", x"87", x"97", x"d2", x"f3", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f5", x"f5", x"f5", x"f4", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"e8", x"d5", x"bb", x"b2", x"b5", x"ba", x"b7", x"91", x"69", x"67", x"62", x"56", x"50", x"4b", 
        x"46", x"40", x"3b", x"36", x"2f", x"27", x"1a", x"06", x"02", x"03", x"05", x"06", x"09", x"0b", x"07", 
        x"08", x"07", x"0a", x"08", x"05", x"19", x"2f", x"39", x"3a", x"33", x"4d", x"5d", x"67", x"6e", x"6c", 
        x"6b", x"6b", x"6e", x"6c", x"69", x"6a", x"6d", x"6d", x"6c", x"6c", x"70", x"49", x"0b", x"1a", x"39", 
        x"39", x"37", x"3f", x"45", x"44", x"45", x"4c", x"47", x"30", x"27", x"28", x"2a", x"2b", x"2f", x"38", 
        x"37", x"37", x"47", x"3c", x"36", x"3c", x"43", x"46", x"41", x"3a", x"36", x"2c", x"25", x"1a", x"08", 
        x"11", x"33", x"41", x"41", x"47", x"47", x"49", x"52", x"53", x"53", x"52", x"54", x"65", x"65", x"58", 
        x"5b", x"60", x"5a", x"4d", x"40", x"46", x"4f", x"4d", x"4e", x"4e", x"4d", x"4e", x"50", x"51", x"51", 
        x"51", x"43", x"43", x"45", x"43", x"3a", x"43", x"7c", x"93", x"92", x"88", x"8b", x"85", x"80", x"80", 
        x"7a", x"75", x"60", x"42", x"3f", x"3d", x"3d", x"3e", x"40", x"41", x"3e", x"62", x"80", x"7e", x"7e", 
        x"81", x"7f", x"7f", x"82", x"84", x"83", x"65", x"55", x"54", x"53", x"54", x"30", x"0e", x"08", x"26", 
        x"69", x"87", x"67", x"67", x"85", x"75", x"77", x"6d", x"66", x"71", x"87", x"87", x"6c", x"37", x"4a", 
        x"84", x"7b", x"69", x"4a", x"17", x"2b", x"3e", x"37", x"2b", x"49", x"40", x"59", x"3b", x"2f", x"3e", 
        x"3e", x"2d", x"45", x"67", x"77", x"47", x"3e", x"3f", x"2b", x"37", x"43", x"6b", x"53", x"48", x"4c", 
        x"73", x"59", x"4f", x"6b", x"4f", x"3f", x"51", x"6b", x"39", x"36", x"2c", x"2b", x"45", x"5b", x"4b", 
        x"5d", x"3c", x"2e", x"42", x"35", x"44", x"45", x"1f", x"2c", x"30", x"32", x"49", x"46", x"50", x"7a", 
        x"5a", x"3f", x"33", x"5d", x"67", x"5c", x"75", x"7b", x"62", x"61", x"68", x"59", x"43", x"5c", x"85", 
        x"5b", x"5a", x"64", x"8b", x"99", x"79", x"d2", x"9b", x"3e", x"58", x"51", x"37", x"62", x"62", x"58", 
        x"5a", x"81", x"7f", x"68", x"4b", x"81", x"8b", x"83", x"85", x"8b", x"8e", x"90", x"95", x"8f", x"98", 
        x"a0", x"a0", x"a7", x"a7", x"a5", x"9c", x"b3", x"98", x"34", x"43", x"72", x"74", x"70", x"7c", x"7a", 
        x"77", x"75", x"72", x"76", x"89", x"8c", x"8b", x"80", x"7f", x"79", x"75", x"76", x"74", x"6f", x"72", 
        x"71", x"69", x"64", x"a7", x"e0", x"d6", x"d4", x"d8", x"d4", x"db", x"da", x"ca", x"cf", x"ce", x"cf", 
        x"cf", x"cf", x"d1", x"d2", x"d1", x"d1", x"d1", x"d3", x"d0", x"d0", x"d0", x"d1", x"d1", x"cf", x"d2", 
        x"d4", x"d4", x"d2", x"d1", x"d1", x"d1", x"d1", x"d3", x"d2", x"d3", x"d4", x"d5", x"d2", x"d0", x"d2", 
        x"d3", x"d3", x"d3", x"d4", x"d4", x"d5", x"d7", x"d2", x"d1", x"d2", x"cf", x"db", x"cf", x"96", x"80", 
        x"76", x"74", x"61", x"67", x"78", x"a6", x"9b", x"75", x"72", x"72", x"71", x"69", x"66", x"69", x"72", 
        x"74", x"71", x"6e", x"6e", x"77", x"7e", x"7b", x"77", x"75", x"7b", x"80", x"7f", x"89", x"8f", x"91", 
        x"86", x"76", x"74", x"79", x"7c", x"7d", x"7b", x"75", x"70", x"70", x"73", x"76", x"76", x"6f", x"67", 
        x"65", x"68", x"6d", x"75", x"a8", x"e1", x"a9", x"89", x"8e", x"86", x"81", x"86", x"91", x"98", x"9b", 
        x"90", x"83", x"87", x"8f", x"93", x"90", x"85", x"80", x"86", x"90", x"90", x"8c", x"80", x"78", x"7a", 
        x"82", x"86", x"84", x"7c", x"75", x"79", x"83", x"8a", x"8b", x"85", x"7a", x"7c", x"89", x"91", x"9b", 
        x"c4", x"db", x"9f", x"98", x"a1", x"a0", x"9e", x"98", x"94", x"99", x"9d", x"9d", x"99", x"91", x"87", 
        x"84", x"81", x"81", x"7e", x"7c", x"84", x"8d", x"8c", x"8e", x"8d", x"8b", x"8b", x"90", x"93", x"92", 
        x"94", x"94", x"94", x"9c", x"a1", x"9e", x"97", x"91", x"b4", x"e0", x"94", x"7d", x"81", x"80", x"7f", 
        x"78", x"78", x"81", x"8a", x"8d", x"8b", x"8d", x"84", x"87", x"88", x"89", x"86", x"8d", x"8c", x"99", 
        x"97", x"9d", x"98", x"98", x"97", x"90", x"7f", x"7b", x"75", x"70", x"77", x"76", x"72", x"9d", x"d9", 
        x"c8", x"b7", x"b5", x"b5", x"b1", x"b3", x"b8", x"b8", x"bd", x"bb", x"b4", x"b6", x"b9", x"b9", x"bb", 
        x"ba", x"c0", x"c5", x"c3", x"bf", x"be", x"bb", x"bd", x"be", x"be", x"bf", x"bd", x"bd", x"ba", x"b4", 
        x"b1", x"c4", x"c5", x"81", x"7a", x"7e", x"81", x"87", x"8a", x"8a", x"87", x"86", x"8d", x"95", x"99", 
        x"93", x"8c", x"8a", x"8e", x"94", x"8f", x"87", x"86", x"86", x"83", x"80", x"79", x"79", x"81", x"89", 
        x"9b", x"d6", x"b2", x"83", x"82", x"86", x"8b", x"8f", x"8a", x"88", x"87", x"86", x"85", x"7e", x"7e", 
        x"85", x"87", x"84", x"7d", x"7e", x"7f", x"7e", x"84", x"89", x"85", x"83", x"80", x"82", x"b2", x"da", 
        x"8d", x"83", x"80", x"81", x"83", x"8a", x"88", x"90", x"98", x"9b", x"99", x"9c", x"96", x"9e", x"91", 
        x"83", x"7f", x"7b", x"76", x"74", x"75", x"71", x"6f", x"77", x"a8", x"cc", x"84", x"78", x"7c", x"79", 
        x"76", x"76", x"78", x"78", x"75", x"75", x"7a", x"78", x"77", x"79", x"7b", x"7c", x"7b", x"7b", x"80", 
        x"7f", x"7b", x"7c", x"a5", x"cd", x"a6", x"95", x"8d", x"85", x"8b", x"96", x"93", x"8b", x"91", x"97", 
        x"8f", x"8a", x"90", x"8f", x"86", x"80", x"85", x"8e", x"8b", x"85", x"8b", x"ca", x"f2", x"f2", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f5", x"f5", x"f5", x"f4", x"f2", x"f2", x"f1", x"ef", 
        x"f2", x"e8", x"d6", x"be", x"b3", x"b5", x"b1", x"b6", x"ac", x"7e", x"68", x"68", x"61", x"5b", x"50", 
        x"45", x"3c", x"37", x"34", x"34", x"31", x"22", x"09", x"04", x"05", x"08", x"07", x"07", x"08", x"07", 
        x"07", x"06", x"09", x"07", x"0b", x"2d", x"3a", x"41", x"47", x"36", x"48", x"5f", x"67", x"6b", x"6b", 
        x"6d", x"6c", x"70", x"70", x"6c", x"69", x"69", x"69", x"69", x"6c", x"70", x"4b", x"0d", x"18", x"3d", 
        x"44", x"40", x"40", x"3c", x"3d", x"3f", x"42", x"38", x"20", x"17", x"1a", x"17", x"14", x"18", x"21", 
        x"22", x"21", x"25", x"1a", x"10", x"0f", x"11", x"13", x"12", x"11", x"15", x"12", x"0f", x"0d", x"08", 
        x"08", x"14", x"1f", x"1f", x"24", x"28", x"2a", x"30", x"35", x"38", x"36", x"36", x"40", x"3f", x"37", 
        x"43", x"49", x"40", x"37", x"37", x"43", x"4a", x"49", x"48", x"49", x"49", x"4a", x"4c", x"4c", x"4a", 
        x"46", x"3b", x"3d", x"43", x"43", x"3a", x"46", x"7c", x"90", x"93", x"8e", x"8e", x"8b", x"86", x"83", 
        x"7b", x"77", x"62", x"42", x"41", x"42", x"44", x"40", x"40", x"42", x"3c", x"5b", x"82", x"81", x"7d", 
        x"7e", x"7e", x"7f", x"80", x"80", x"81", x"64", x"51", x"52", x"54", x"56", x"32", x"0e", x"07", x"23", 
        x"7a", x"6b", x"51", x"51", x"70", x"77", x"78", x"6f", x"83", x"7c", x"70", x"67", x"64", x"53", x"62", 
        x"74", x"63", x"7e", x"4f", x"24", x"26", x"49", x"60", x"40", x"31", x"27", x"3c", x"38", x"3d", x"4b", 
        x"45", x"40", x"51", x"4a", x"47", x"46", x"5c", x"5d", x"23", x"33", x"49", x"70", x"5c", x"48", x"64", 
        x"50", x"37", x"64", x"6f", x"3c", x"20", x"3d", x"56", x"48", x"58", x"3d", x"23", x"35", x"48", x"49", 
        x"51", x"69", x"5d", x"4e", x"3d", x"38", x"2c", x"14", x"25", x"26", x"25", x"3e", x"42", x"51", x"54", 
        x"40", x"27", x"3c", x"6b", x"5a", x"57", x"57", x"5b", x"55", x"59", x"6a", x"5e", x"61", x"67", x"61", 
        x"54", x"60", x"5f", x"85", x"8f", x"7e", x"d4", x"a8", x"4d", x"5b", x"57", x"4c", x"6e", x"8f", x"9a", 
        x"5b", x"6e", x"7c", x"66", x"4d", x"84", x"8e", x"7b", x"7e", x"87", x"7d", x"87", x"85", x"7f", x"8d", 
        x"80", x"7e", x"7c", x"9c", x"9d", x"6d", x"8b", x"81", x"32", x"45", x"74", x"77", x"71", x"7a", x"79", 
        x"76", x"72", x"72", x"77", x"79", x"72", x"7e", x"82", x"81", x"7b", x"78", x"7a", x"71", x"71", x"72", 
        x"73", x"6c", x"68", x"a7", x"de", x"d4", x"d5", x"d7", x"d5", x"dc", x"dc", x"cb", x"cf", x"cd", x"cd", 
        x"cf", x"d0", x"d1", x"d1", x"d2", x"d1", x"d1", x"d1", x"d0", x"d1", x"d0", x"d0", x"d1", x"cf", x"cf", 
        x"cf", x"d1", x"d1", x"d2", x"d3", x"d1", x"d0", x"d4", x"d2", x"d3", x"d5", x"d6", x"d2", x"d0", x"d1", 
        x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"d5", x"d6", x"d6", x"d4", x"ce", x"de", x"d6", x"9c", x"84", 
        x"79", x"81", x"7c", x"7c", x"7e", x"a0", x"97", x"78", x"7b", x"7e", x"81", x"7f", x"80", x"84", x"85", 
        x"80", x"7a", x"79", x"7f", x"85", x"82", x"7d", x"72", x"6a", x"6e", x"73", x"75", x"74", x"68", x"62", 
        x"5f", x"5f", x"65", x"69", x"69", x"66", x"65", x"66", x"6a", x"6f", x"72", x"74", x"75", x"75", x"78", 
        x"7b", x"7f", x"81", x"81", x"a8", x"e2", x"b2", x"8f", x"90", x"88", x"7f", x"7f", x"84", x"83", x"82", 
        x"7a", x"72", x"79", x"81", x"85", x"81", x"79", x"78", x"7f", x"87", x"8a", x"86", x"80", x"83", x"8f", 
        x"9c", x"a0", x"9f", x"96", x"8a", x"88", x"8d", x"91", x"91", x"8e", x"85", x"85", x"8f", x"93", x"98", 
        x"c3", x"db", x"91", x"83", x"89", x"89", x"8b", x"8c", x"8c", x"8d", x"90", x"8d", x"8d", x"8c", x"89", 
        x"8d", x"94", x"99", x"98", x"97", x"9a", x"9e", x"a0", x"a0", x"9f", x"9b", x"97", x"9a", x"9f", x"9f", 
        x"9e", x"97", x"8c", x"88", x"88", x"85", x"83", x"85", x"af", x"df", x"8a", x"67", x"6b", x"6e", x"74", 
        x"76", x"75", x"7f", x"8b", x"8d", x"8e", x"96", x"97", x"9a", x"95", x"98", x"98", x"9d", x"92", x"9c", 
        x"9a", x"99", x"90", x"8a", x"88", x"88", x"7d", x"77", x"6d", x"66", x"6b", x"69", x"68", x"98", x"dc", 
        x"cd", x"ba", x"b9", x"bd", x"c0", x"c4", x"c3", x"c4", x"c8", x"c7", x"c1", x"c0", x"bf", x"c0", x"c4", 
        x"c2", x"bd", x"bb", x"b8", x"b9", x"b9", x"b1", x"b4", x"bb", x"be", x"c1", x"b9", x"b8", x"bb", x"bc", 
        x"ba", x"ca", x"cd", x"8d", x"84", x"87", x"8c", x"91", x"90", x"8b", x"8c", x"8f", x"8f", x"8d", x"88", 
        x"82", x"81", x"83", x"85", x"84", x"82", x"82", x"89", x"8a", x"82", x"7e", x"7e", x"83", x"8c", x"94", 
        x"a3", x"dc", x"b9", x"87", x"86", x"89", x"8d", x"90", x"8a", x"86", x"84", x"82", x"80", x"7a", x"7c", 
        x"86", x"8b", x"88", x"82", x"81", x"83", x"87", x"8f", x"91", x"8a", x"85", x"83", x"84", x"b1", x"dd", 
        x"8d", x"81", x"81", x"81", x"84", x"8d", x"91", x"98", x"9d", x"a0", x"9c", x"9e", x"9b", x"a3", x"97", 
        x"85", x"82", x"7d", x"77", x"73", x"73", x"71", x"6e", x"73", x"a2", x"cc", x"82", x"72", x"76", x"74", 
        x"73", x"77", x"79", x"79", x"74", x"71", x"76", x"75", x"72", x"77", x"7e", x"83", x"80", x"7a", x"77", 
        x"79", x"77", x"78", x"9f", x"cb", x"a4", x"92", x"97", x"8c", x"88", x"91", x"96", x"92", x"8d", x"95", 
        x"97", x"8a", x"84", x"8a", x"90", x"86", x"7e", x"87", x"92", x"8f", x"8a", x"c0", x"ee", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f4", x"f4", x"f3", x"f2", x"f2", x"f1", x"f0", 
        x"f3", x"ea", x"d9", x"c2", x"b5", x"b5", x"b8", x"bf", x"c2", x"9d", x"74", x"6a", x"60", x"55", x"4e", 
        x"49", x"45", x"42", x"40", x"3d", x"36", x"27", x"0a", x"02", x"04", x"09", x"08", x"07", x"07", x"07", 
        x"07", x"08", x"08", x"08", x"1b", x"3f", x"42", x"45", x"46", x"37", x"47", x"5d", x"67", x"6b", x"6a", 
        x"6c", x"6d", x"70", x"6e", x"6b", x"68", x"67", x"67", x"69", x"69", x"6d", x"4a", x"10", x"17", x"39", 
        x"40", x"34", x"2d", x"31", x"33", x"2e", x"24", x"1b", x"13", x"15", x"13", x"0e", x"07", x"09", x"10", 
        x"10", x"0f", x"0e", x"12", x"17", x"1b", x"1b", x"1b", x"1c", x"1b", x"1d", x"1d", x"1b", x"13", x"0a", 
        x"07", x"0b", x"12", x"0f", x"0e", x"11", x"0c", x"0a", x"0c", x"0d", x"0e", x"12", x"18", x"19", x"1d", 
        x"38", x"3e", x"27", x"26", x"2b", x"2e", x"2e", x"2d", x"2e", x"30", x"32", x"35", x"38", x"38", x"34", 
        x"33", x"2e", x"33", x"39", x"36", x"30", x"41", x"7d", x"93", x"96", x"91", x"8c", x"8d", x"89", x"84", 
        x"7c", x"78", x"65", x"40", x"3c", x"3e", x"3f", x"3b", x"3c", x"40", x"39", x"51", x"7d", x"7e", x"7a", 
        x"7d", x"7e", x"80", x"80", x"7f", x"81", x"67", x"4f", x"51", x"52", x"56", x"36", x"11", x"08", x"1f", 
        x"67", x"55", x"63", x"65", x"57", x"5f", x"59", x"42", x"48", x"50", x"65", x"5b", x"45", x"4e", x"64", 
        x"59", x"64", x"5c", x"39", x"54", x"4b", x"3f", x"3f", x"49", x"3c", x"30", x"48", x"43", x"3d", x"57", 
        x"58", x"48", x"5b", x"4e", x"38", x"27", x"28", x"38", x"3d", x"4a", x"4a", x"79", x"79", x"3d", x"39", 
        x"22", x"33", x"5f", x"48", x"2b", x"2b", x"2b", x"43", x"7d", x"6f", x"6a", x"55", x"47", x"6a", x"60", 
        x"3c", x"5e", x"58", x"44", x"31", x"42", x"34", x"21", x"21", x"2a", x"2e", x"26", x"26", x"2a", x"30", 
        x"50", x"39", x"3d", x"30", x"47", x"76", x"75", x"7c", x"75", x"73", x"7b", x"69", x"51", x"64", x"6e", 
        x"7c", x"89", x"8a", x"b0", x"95", x"73", x"b6", x"79", x"42", x"63", x"62", x"53", x"70", x"85", x"96", 
        x"5d", x"83", x"7c", x"50", x"55", x"89", x"8d", x"7d", x"83", x"89", x"7e", x"8c", x"8c", x"81", x"97", 
        x"96", x"9c", x"98", x"ae", x"a7", x"8d", x"b2", x"99", x"36", x"40", x"6f", x"73", x"75", x"93", x"93", 
        x"97", x"98", x"94", x"98", x"82", x"70", x"88", x"95", x"94", x"7b", x"67", x"68", x"68", x"8f", x"7b", 
        x"76", x"6f", x"6c", x"a7", x"dc", x"d5", x"d9", x"d6", x"d3", x"db", x"db", x"cc", x"d0", x"ce", x"ce", 
        x"cf", x"d0", x"d0", x"d1", x"d2", x"d1", x"d0", x"d0", x"d0", x"d2", x"d0", x"d0", x"d1", x"d0", x"d0", 
        x"d2", x"d4", x"d3", x"d1", x"d0", x"cc", x"cb", x"d5", x"d4", x"d2", x"d3", x"d4", x"d2", x"d0", x"d2", 
        x"d3", x"d3", x"d3", x"d4", x"d4", x"d4", x"d5", x"d6", x"d6", x"d2", x"d0", x"df", x"d6", x"9b", x"89", 
        x"79", x"79", x"6f", x"6b", x"74", x"a2", x"9e", x"7d", x"75", x"6e", x"74", x"81", x"88", x"81", x"76", 
        x"72", x"74", x"7b", x"84", x"84", x"81", x"7b", x"78", x"7b", x"83", x"88", x"8d", x"87", x"75", x"6e", 
        x"73", x"7c", x"7f", x"7b", x"73", x"6c", x"68", x"6a", x"71", x"75", x"75", x"6c", x"63", x"60", x"64", 
        x"6c", x"70", x"6b", x"6c", x"9d", x"df", x"b2", x"8b", x"8c", x"85", x"85", x"8e", x"97", x"98", x"95", 
        x"8d", x"86", x"8d", x"95", x"96", x"8f", x"84", x"83", x"88", x"8b", x"8c", x"85", x"7a", x"75", x"78", 
        x"80", x"83", x"80", x"79", x"76", x"7e", x"8a", x"92", x"93", x"8f", x"82", x"7d", x"85", x"8e", x"95", 
        x"bf", x"dd", x"a0", x"95", x"a4", x"a7", x"a5", x"9e", x"94", x"8e", x"90", x"8f", x"8f", x"8f", x"8a", 
        x"89", x"8b", x"8e", x"8f", x"8b", x"84", x"81", x"85", x"8f", x"96", x"96", x"92", x"91", x"93", x"92", 
        x"92", x"91", x"91", x"95", x"99", x"9b", x"9f", x"a0", x"ba", x"e2", x"95", x"77", x"7b", x"7c", x"85", 
        x"8d", x"95", x"90", x"8f", x"90", x"91", x"92", x"88", x"81", x"72", x"73", x"7a", x"7f", x"6e", x"6f", 
        x"6b", x"6b", x"6e", x"72", x"75", x"7a", x"73", x"75", x"7b", x"7f", x"7c", x"72", x"6c", x"94", x"d9", 
        x"d2", x"c0", x"bf", x"bf", x"bc", x"c1", x"c4", x"be", x"b9", x"b2", x"b8", x"bf", x"bf", x"ba", x"bb", 
        x"bd", x"c0", x"be", x"ba", x"bc", x"be", x"c0", x"ca", x"ca", x"c4", x"c8", x"c6", x"c1", x"c1", x"c0", 
        x"bc", x"ca", x"cf", x"8f", x"86", x"8d", x"8c", x"87", x"80", x"82", x"89", x"8c", x"89", x"89", x"8c", 
        x"90", x"91", x"90", x"8d", x"89", x"8d", x"94", x"97", x"8d", x"80", x"7f", x"83", x"8a", x"8d", x"8a", 
        x"95", x"d4", x"b9", x"7e", x"7a", x"7e", x"81", x"86", x"87", x"87", x"86", x"85", x"84", x"80", x"84", 
        x"8d", x"8f", x"8b", x"84", x"82", x"86", x"8c", x"91", x"8e", x"85", x"80", x"84", x"85", x"ab", x"db", 
        x"8b", x"79", x"7a", x"83", x"8f", x"96", x"9b", x"9d", x"a2", x"a0", x"9b", x"a0", x"9d", x"a3", x"97", 
        x"84", x"7f", x"7b", x"78", x"76", x"74", x"71", x"6a", x"6e", x"9e", x"d0", x"86", x"73", x"78", x"7a", 
        x"7a", x"7a", x"7a", x"7b", x"77", x"75", x"7c", x"7e", x"7f", x"80", x"82", x"81", x"7c", x"7c", x"7e", 
        x"7b", x"76", x"76", x"9d", x"cf", x"a6", x"88", x"94", x"98", x"96", x"91", x"98", x"9c", x"92", x"8f", 
        x"97", x"96", x"8a", x"84", x"88", x"8f", x"8a", x"81", x"83", x"8a", x"91", x"c3", x"ef", x"f3", x"f1", 
        x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f3", x"f2", x"f1", x"ef", x"ed", 
        x"f2", x"e9", x"db", x"c7", x"b8", x"b8", x"ba", x"b3", x"b9", x"b5", x"86", x"69", x"65", x"5f", x"58", 
        x"50", x"4b", x"48", x"47", x"44", x"3d", x"30", x"0e", x"03", x"03", x"0b", x"0a", x"0a", x"08", x"09", 
        x"0a", x"0a", x"09", x"12", x"31", x"3b", x"39", x"3b", x"41", x"36", x"41", x"57", x"66", x"6d", x"6a", 
        x"6a", x"6c", x"70", x"6d", x"6a", x"69", x"68", x"69", x"6a", x"68", x"6c", x"4e", x"15", x"0e", x"18", 
        x"16", x"0e", x"08", x"08", x"08", x"09", x"0b", x"10", x"0b", x"09", x"08", x"09", x"08", x"0d", x"14", 
        x"15", x"13", x"16", x"1c", x"1d", x"1b", x"1a", x"19", x"1a", x"1b", x"1b", x"18", x"1a", x"10", x"06", 
        x"07", x"0d", x"17", x"19", x"18", x"18", x"13", x"12", x"15", x"12", x"0f", x"11", x"11", x"0d", x"10", 
        x"2f", x"2d", x"08", x"08", x"09", x"08", x"0b", x"0a", x"10", x"11", x"11", x"13", x"17", x"19", x"17", 
        x"23", x"24", x"20", x"23", x"20", x"1e", x"2f", x"6e", x"8f", x"91", x"8b", x"89", x"8c", x"89", x"84", 
        x"7c", x"7a", x"6b", x"43", x"42", x"46", x"49", x"47", x"47", x"48", x"42", x"55", x"81", x"81", x"7d", 
        x"7e", x"7e", x"7f", x"7e", x"7d", x"81", x"6a", x"4f", x"53", x"53", x"56", x"38", x"11", x"08", x"1c", 
        x"58", x"53", x"63", x"6a", x"55", x"61", x"4e", x"38", x"2b", x"3f", x"8c", x"6c", x"36", x"33", x"47", 
        x"55", x"79", x"50", x"4c", x"52", x"65", x"3b", x"18", x"32", x"2a", x"21", x"2e", x"21", x"1e", x"40", 
        x"55", x"69", x"6f", x"46", x"35", x"3f", x"4a", x"3e", x"3d", x"44", x"46", x"65", x"72", x"4c", x"54", 
        x"35", x"43", x"4b", x"45", x"44", x"34", x"4a", x"5f", x"63", x"65", x"70", x"6a", x"47", x"5a", x"53", 
        x"38", x"3f", x"40", x"43", x"46", x"5d", x"4f", x"34", x"24", x"32", x"3f", x"36", x"30", x"33", x"2f", 
        x"51", x"5e", x"61", x"6e", x"6b", x"71", x"7b", x"87", x"63", x"5b", x"66", x"5f", x"62", x"6f", x"82", 
        x"a7", x"91", x"7e", x"91", x"95", x"6e", x"8d", x"68", x"49", x"60", x"79", x"7d", x"81", x"79", x"82", 
        x"5f", x"86", x"79", x"5e", x"55", x"85", x"8f", x"80", x"85", x"88", x"82", x"8b", x"8a", x"7f", x"94", 
        x"98", x"9d", x"98", x"9a", x"a5", x"a4", x"bd", x"9c", x"37", x"41", x"70", x"73", x"77", x"a2", x"9f", 
        x"96", x"9e", x"a0", x"a5", x"8d", x"89", x"9e", x"9b", x"9c", x"7b", x"5e", x"62", x"5d", x"9e", x"7c", 
        x"76", x"72", x"6c", x"a5", x"dd", x"d6", x"d9", x"d6", x"d2", x"da", x"db", x"cc", x"d0", x"ce", x"ce", 
        x"d0", x"d1", x"d0", x"d1", x"d2", x"d1", x"d0", x"ce", x"cf", x"d2", x"d0", x"d0", x"d3", x"d3", x"d2", 
        x"d2", x"d6", x"d3", x"d0", x"d1", x"d0", x"ce", x"d4", x"d3", x"d2", x"d2", x"d3", x"d3", x"d2", x"d2", 
        x"d3", x"d3", x"d4", x"d5", x"d5", x"d5", x"d2", x"d4", x"d6", x"d4", x"d0", x"de", x"d6", x"9e", x"83", 
        x"71", x"77", x"6f", x"74", x"7c", x"a5", x"a1", x"7d", x"7b", x"7c", x"7e", x"7b", x"7e", x"81", x"7c", 
        x"7d", x"7e", x"7c", x"80", x"7d", x"7a", x"7b", x"77", x"77", x"7a", x"79", x"78", x"73", x"6f", x"74", 
        x"7a", x"7c", x"7b", x"76", x"71", x"6f", x"70", x"75", x"7a", x"7d", x"7c", x"73", x"6f", x"73", x"7a", 
        x"82", x"84", x"7c", x"78", x"a0", x"e1", x"b3", x"86", x"82", x"7d", x"7f", x"8b", x"8d", x"89", x"81", 
        x"7a", x"78", x"7d", x"84", x"86", x"84", x"7e", x"82", x"8a", x"8c", x"8c", x"88", x"81", x"81", x"86", 
        x"8f", x"96", x"96", x"8f", x"88", x"8c", x"94", x"97", x"95", x"90", x"85", x"7f", x"83", x"8a", x"91", 
        x"bc", x"dc", x"9c", x"85", x"8c", x"8d", x"8c", x"8a", x"85", x"88", x"8e", x"94", x"96", x"96", x"90", 
        x"89", x"8b", x"8d", x"90", x"91", x"8f", x"90", x"95", x"9b", x"9e", x"9f", x"9b", x"94", x"8f", x"90", 
        x"94", x"95", x"94", x"93", x"90", x"90", x"94", x"95", x"b0", x"e0", x"94", x"6e", x"6e", x"74", x"83", 
        x"88", x"8f", x"87", x"85", x"82", x"84", x"86", x"77", x"74", x"6e", x"6d", x"74", x"82", x"83", x"7f", 
        x"79", x"75", x"77", x"7a", x"7f", x"87", x"7d", x"73", x"71", x"75", x"75", x"70", x"6d", x"91", x"d3", 
        x"c6", x"b4", x"bd", x"c3", x"bb", x"ba", x"b9", x"ba", x"bc", x"b9", x"ba", x"bf", x"c4", x"c8", x"c4", 
        x"bb", x"bb", x"bf", x"bf", x"be", x"c1", x"bd", x"c3", x"c6", x"bf", x"bc", x"b9", x"ba", x"bd", x"bd", 
        x"b8", x"c3", x"ce", x"92", x"88", x"8a", x"87", x"85", x"89", x"8e", x"8d", x"8c", x"8f", x"90", x"93", 
        x"93", x"8f", x"8c", x"8c", x"8c", x"8e", x"8d", x"8a", x"7f", x"76", x"7b", x"87", x"8d", x"8b", x"87", 
        x"92", x"d3", x"be", x"83", x"80", x"84", x"85", x"8a", x"8d", x"90", x"8d", x"87", x"85", x"80", x"84", 
        x"89", x"86", x"82", x"7d", x"79", x"7c", x"81", x"83", x"83", x"81", x"7f", x"84", x"88", x"a7", x"db", 
        x"90", x"7e", x"83", x"91", x"9c", x"9e", x"9b", x"9c", x"a0", x"a0", x"9b", x"9d", x"99", x"9c", x"92", 
        x"82", x"7a", x"76", x"75", x"75", x"75", x"74", x"6c", x"6f", x"9d", x"d4", x"8b", x"74", x"76", x"78", 
        x"78", x"76", x"78", x"7b", x"77", x"72", x"75", x"78", x"7e", x"7d", x"81", x"82", x"7f", x"7d", x"7b", 
        x"7d", x"79", x"79", x"9e", x"d3", x"ae", x"88", x"8d", x"96", x"98", x"90", x"92", x"9a", x"98", x"92", 
        x"90", x"90", x"90", x"8b", x"82", x"83", x"8b", x"8d", x"82", x"7d", x"86", x"c1", x"f1", x"f2", x"f1", 
        x"f1", x"f2", x"f2", x"f3", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f1", x"f1", x"f2", x"f0", 
        x"f4", x"ea", x"da", x"c6", x"b4", x"b6", x"bd", x"b5", x"b4", x"bb", x"9c", x"72", x"5f", x"5c", x"57", 
        x"53", x"50", x"4e", x"4e", x"49", x"42", x"36", x"11", x"03", x"03", x"0c", x"0b", x"0b", x"0b", x"09", 
        x"0b", x"0a", x"0a", x"1f", x"3a", x"3b", x"3d", x"40", x"46", x"3a", x"43", x"58", x"66", x"6c", x"6c", 
        x"6b", x"6c", x"71", x"70", x"6d", x"69", x"65", x"66", x"69", x"68", x"6d", x"52", x"17", x"07", x"0f", 
        x"14", x"1a", x"1f", x"1e", x"1a", x"1b", x"21", x"2a", x"24", x"1a", x"12", x"12", x"0c", x"0b", x"0a", 
        x"08", x"06", x"11", x"17", x"17", x"16", x"1a", x"19", x"18", x"19", x"1a", x"18", x"1c", x"13", x"07", 
        x"06", x"0b", x"16", x"1c", x"1b", x"18", x"14", x"17", x"1a", x"15", x"0e", x"10", x"13", x"11", x"0e", 
        x"28", x"31", x"0d", x"10", x"12", x"11", x"11", x"0f", x"10", x"0e", x"08", x"06", x"09", x"0b", x"08", 
        x"15", x"17", x"0e", x"11", x"12", x"13", x"21", x"5d", x"8b", x"8d", x"88", x"87", x"8a", x"87", x"7f", 
        x"76", x"71", x"60", x"36", x"36", x"3c", x"41", x"41", x"3e", x"38", x"36", x"47", x"75", x"78", x"75", 
        x"75", x"76", x"77", x"76", x"78", x"80", x"69", x"4d", x"55", x"56", x"58", x"3a", x"13", x"08", x"1a", 
        x"58", x"6d", x"70", x"68", x"5b", x"42", x"53", x"66", x"29", x"20", x"61", x"54", x"49", x"40", x"32", 
        x"3a", x"44", x"2f", x"3a", x"45", x"47", x"2d", x"36", x"31", x"23", x"19", x"13", x"10", x"10", x"26", 
        x"2d", x"3e", x"4c", x"45", x"4c", x"63", x"98", x"65", x"32", x"2d", x"29", x"31", x"78", x"6d", x"80", 
        x"53", x"32", x"4e", x"56", x"57", x"4d", x"4b", x"4d", x"53", x"35", x"3b", x"63", x"62", x"50", x"58", 
        x"47", x"2b", x"3d", x"5d", x"6b", x"7f", x"59", x"32", x"2c", x"36", x"4a", x"3c", x"35", x"3f", x"33", 
        x"40", x"58", x"77", x"8d", x"6f", x"55", x"5f", x"86", x"62", x"61", x"80", x"6f", x"66", x"55", x"78", 
        x"b6", x"93", x"65", x"55", x"75", x"52", x"78", x"73", x"45", x"5c", x"87", x"94", x"88", x"7d", x"71", 
        x"4c", x"74", x"78", x"6f", x"51", x"8c", x"96", x"7c", x"87", x"8a", x"80", x"8d", x"88", x"7e", x"96", 
        x"98", x"9e", x"93", x"9c", x"ba", x"a5", x"be", x"a1", x"39", x"42", x"6f", x"74", x"75", x"a9", x"b1", 
        x"9b", x"9b", x"9e", x"a1", x"8d", x"9b", x"a2", x"8c", x"95", x"7b", x"5e", x"62", x"53", x"9a", x"7b", 
        x"76", x"77", x"6b", x"a4", x"de", x"d3", x"d5", x"d4", x"d4", x"dc", x"dc", x"cc", x"d0", x"cc", x"cc", 
        x"d0", x"d1", x"d0", x"d1", x"d2", x"d1", x"cf", x"cd", x"ce", x"d2", x"d0", x"d1", x"d4", x"d4", x"d2", 
        x"d2", x"d6", x"d3", x"d1", x"d4", x"d6", x"d4", x"d4", x"d4", x"d3", x"d2", x"d2", x"d1", x"d2", x"d3", 
        x"d3", x"d4", x"d4", x"d5", x"d5", x"d5", x"d6", x"d4", x"d4", x"d4", x"d0", x"dd", x"d9", x"a3", x"91", 
        x"83", x"84", x"71", x"67", x"69", x"96", x"91", x"69", x"69", x"6a", x"6a", x"68", x"6f", x"75", x"75", 
        x"7c", x"7d", x"78", x"7c", x"7a", x"7b", x"83", x"85", x"85", x"7d", x"77", x"7b", x"85", x"84", x"83", 
        x"7d", x"74", x"72", x"71", x"73", x"74", x"73", x"6d", x"68", x"64", x"63", x"61", x"62", x"63", x"63", 
        x"66", x"69", x"64", x"65", x"97", x"e1", x"b4", x"83", x"81", x"84", x"8c", x"90", x"93", x"93", x"8f", 
        x"91", x"97", x"9c", x"9a", x"97", x"8d", x"82", x"84", x"8b", x"8d", x"8a", x"80", x"73", x"71", x"78", 
        x"80", x"84", x"7e", x"73", x"6a", x"6d", x"77", x"7e", x"80", x"7f", x"7c", x"7b", x"82", x"8d", x"94", 
        x"bc", x"dd", x"a2", x"8e", x"9b", x"a3", x"a8", x"a8", x"a1", x"9c", x"9a", x"98", x"95", x"95", x"94", 
        x"8d", x"89", x"8b", x"8e", x"8e", x"8c", x"85", x"7f", x"84", x"83", x"84", x"86", x"80", x"7e", x"89", 
        x"96", x"99", x"9a", x"99", x"94", x"91", x"94", x"99", x"b3", x"e2", x"9e", x"7f", x"82", x"84", x"8e", 
        x"8d", x"8e", x"85", x"81", x"76", x"70", x"73", x"77", x"78", x"74", x"6c", x"64", x"6b", x"72", x"75", 
        x"73", x"6e", x"69", x"66", x"6d", x"7e", x"7c", x"6f", x"67", x"6a", x"6a", x"6c", x"71", x"90", x"d2", 
        x"cf", x"bb", x"bf", x"c5", x"c3", x"c3", x"b7", x"b9", x"be", x"c0", x"c2", x"be", x"b7", x"b8", x"b9", 
        x"b6", x"b4", x"b3", x"b1", x"b7", x"c7", x"c1", x"be", x"bd", x"bc", x"c0", x"c1", x"be", x"c0", x"c0", 
        x"bc", x"c7", x"d5", x"96", x"87", x"89", x"8c", x"8c", x"88", x"84", x"84", x"85", x"87", x"86", x"88", 
        x"88", x"84", x"84", x"8c", x"96", x"94", x"8a", x"84", x"82", x"88", x"93", x"91", x"8d", x"86", x"87", 
        x"97", x"d5", x"bd", x"80", x"7e", x"83", x"82", x"83", x"84", x"85", x"84", x"7f", x"7c", x"79", x"81", 
        x"8a", x"88", x"84", x"81", x"80", x"84", x"86", x"83", x"84", x"88", x"89", x"8e", x"90", x"a9", x"dd", 
        x"98", x"86", x"93", x"9c", x"9c", x"9b", x"92", x"95", x"97", x"9a", x"95", x"95", x"8f", x"93", x"8f", 
        x"85", x"7e", x"78", x"78", x"77", x"76", x"75", x"6c", x"6d", x"98", x"d2", x"8d", x"76", x"78", x"77", 
        x"77", x"75", x"73", x"76", x"75", x"74", x"7d", x"80", x"81", x"7c", x"7f", x"7f", x"7c", x"7b", x"79", 
        x"7a", x"7b", x"7e", x"9f", x"d2", x"b4", x"91", x"8d", x"93", x"9a", x"96", x"90", x"91", x"99", x"99", 
        x"8f", x"83", x"87", x"92", x"8a", x"7c", x"7d", x"8d", x"90", x"85", x"80", x"b9", x"f1", x"f4", x"f1", 
        x"f2", x"f2", x"f3", x"f3", x"f4", x"f4", x"f3", x"f3", x"f4", x"f4", x"f3", x"f1", x"f1", x"f2", x"ef", 
        x"f4", x"ec", x"de", x"cc", x"b9", x"b4", x"b4", x"b4", x"bb", x"c3", x"b6", x"89", x"68", x"67", x"61", 
        x"5b", x"55", x"4f", x"4b", x"47", x"43", x"3a", x"14", x"05", x"05", x"10", x"0f", x"0f", x"10", x"0e", 
        x"0e", x"0b", x"10", x"31", x"43", x"40", x"3a", x"3d", x"40", x"38", x"43", x"5b", x"65", x"6a", x"6d", 
        x"6e", x"6d", x"72", x"74", x"72", x"6d", x"67", x"68", x"6b", x"69", x"70", x"58", x"18", x"0a", x"22", 
        x"30", x"35", x"3f", x"45", x"4e", x"55", x"53", x"45", x"27", x"12", x"12", x"16", x"10", x"0e", x"0a", 
        x"09", x"0a", x"13", x"18", x"15", x"15", x"1a", x"1c", x"1c", x"1b", x"1d", x"1b", x"1f", x"14", x"06", 
        x"08", x"0e", x"17", x"1a", x"18", x"15", x"14", x"17", x"18", x"13", x"0f", x"0f", x"11", x"11", x"09", 
        x"1e", x"35", x"11", x"14", x"19", x"17", x"11", x"13", x"13", x"10", x"0b", x"09", x"0d", x"0e", x"0b", 
        x"17", x"1c", x"12", x"14", x"12", x"0f", x"16", x"4d", x"85", x"8c", x"8c", x"8e", x"8d", x"84", x"7d", 
        x"7b", x"76", x"64", x"33", x"2d", x"2b", x"2c", x"2d", x"2b", x"25", x"28", x"39", x"66", x"6a", x"6c", 
        x"6a", x"69", x"68", x"66", x"67", x"71", x"61", x"43", x"49", x"48", x"4d", x"37", x"15", x"08", x"12", 
        x"4e", x"55", x"66", x"62", x"3f", x"4b", x"41", x"4d", x"56", x"52", x"2b", x"27", x"4a", x"6f", x"5e", 
        x"30", x"30", x"4c", x"2e", x"2e", x"3f", x"3a", x"34", x"2a", x"2a", x"38", x"41", x"24", x"19", x"23", 
        x"1d", x"2f", x"38", x"49", x"50", x"41", x"5c", x"5f", x"77", x"62", x"55", x"41", x"6b", x"6a", x"46", 
        x"5b", x"46", x"82", x"76", x"62", x"75", x"57", x"70", x"67", x"36", x"46", x"5a", x"3b", x"3f", x"65", 
        x"67", x"61", x"4b", x"54", x"68", x"6c", x"34", x"2d", x"4a", x"48", x"48", x"35", x"4c", x"5c", x"78", 
        x"68", x"4c", x"52", x"65", x"6c", x"6b", x"63", x"6b", x"67", x"5e", x"7d", x"7a", x"6a", x"61", x"68", 
        x"6b", x"67", x"65", x"69", x"71", x"56", x"7d", x"67", x"5a", x"55", x"7e", x"a0", x"9b", x"96", x"7c", 
        x"4e", x"6e", x"7f", x"75", x"52", x"89", x"91", x"7f", x"83", x"8b", x"81", x"87", x"95", x"94", x"90", 
        x"96", x"a0", x"98", x"ae", x"c9", x"a9", x"bc", x"9c", x"39", x"40", x"6e", x"6f", x"71", x"a8", x"b8", 
        x"9c", x"9a", x"9c", x"a1", x"89", x"93", x"98", x"8d", x"9a", x"74", x"5c", x"64", x"55", x"9c", x"81", 
        x"76", x"76", x"6d", x"a2", x"de", x"d4", x"d4", x"d6", x"d2", x"d9", x"dc", x"cd", x"d0", x"ce", x"ce", 
        x"d0", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"d0", x"cf", x"d0", x"d0", x"d1", x"d3", x"d1", x"d1", 
        x"d4", x"d5", x"d2", x"d0", x"d3", x"d3", x"d1", x"d3", x"d3", x"d3", x"d1", x"d1", x"d1", x"d2", x"d2", 
        x"d2", x"d2", x"d3", x"d4", x"d5", x"d6", x"d5", x"d6", x"d5", x"d3", x"cf", x"dd", x"da", x"9f", x"82", 
        x"6b", x"6d", x"6f", x"77", x"84", x"a9", x"aa", x"8e", x"91", x"92", x"91", x"98", x"9f", x"9d", x"98", 
        x"92", x"8b", x"84", x"85", x"89", x"87", x"82", x"76", x"72", x"79", x"71", x"66", x"66", x"65", x"68", 
        x"64", x"60", x"62", x"6f", x"76", x"76", x"78", x"76", x"73", x"71", x"73", x"7a", x"81", x"87", x"82", 
        x"79", x"74", x"73", x"7a", x"a5", x"e2", x"b3", x"7e", x"82", x"88", x"8d", x"8b", x"83", x"78", x"72", 
        x"76", x"7d", x"7e", x"79", x"74", x"73", x"7c", x"86", x"8d", x"90", x"8b", x"81", x"80", x"87", x"8c", 
        x"91", x"93", x"8d", x"88", x"8c", x"95", x"9e", x"a0", x"9d", x"97", x"88", x"82", x"84", x"8c", x"94", 
        x"bb", x"e2", x"a5", x"89", x"8a", x"89", x"8a", x"8c", x"89", x"7f", x"7a", x"7e", x"84", x"86", x"87", 
        x"88", x"89", x"8e", x"97", x"9a", x"95", x"90", x"89", x"90", x"9c", x"a4", x"a7", x"a5", x"9f", x"98", 
        x"95", x"96", x"95", x"94", x"92", x"8d", x"88", x"88", x"a9", x"e1", x"9f", x"77", x"7f", x"7a", x"72", 
        x"64", x"68", x"6e", x"72", x"6f", x"6b", x"6a", x"6c", x"77", x"7c", x"77", x"72", x"72", x"71", x"70", 
        x"78", x"80", x"84", x"82", x"83", x"88", x"88", x"83", x"81", x"7d", x"72", x"6e", x"70", x"92", x"d3", 
        x"d1", x"c0", x"bf", x"b7", x"b6", x"bb", x"b9", x"ba", x"bc", x"bb", x"bf", x"c5", x"c4", x"bd", x"bb", 
        x"b9", x"bd", x"c5", x"c5", x"c0", x"bf", x"bf", x"bf", x"c1", x"bf", x"bb", x"bf", x"bf", x"bf", x"bd", 
        x"b9", x"c0", x"d4", x"95", x"82", x"82", x"83", x"83", x"81", x"7e", x"7f", x"87", x"90", x"8e", x"8c", 
        x"8c", x"8e", x"93", x"98", x"96", x"8e", x"83", x"86", x"86", x"81", x"83", x"80", x"7d", x"7d", x"84", 
        x"93", x"cf", x"c1", x"80", x"7b", x"7d", x"7f", x"87", x"8a", x"89", x"87", x"86", x"84", x"81", x"84", 
        x"88", x"89", x"89", x"8d", x"8e", x"89", x"85", x"82", x"81", x"85", x"85", x"83", x"82", x"a3", x"db", 
        x"9c", x"91", x"91", x"9c", x"94", x"97", x"92", x"95", x"95", x"9b", x"98", x"9a", x"94", x"9b", x"95", 
        x"8b", x"83", x"7b", x"79", x"7a", x"7b", x"7a", x"77", x"79", x"9a", x"d7", x"8f", x"71", x"72", x"75", 
        x"76", x"73", x"75", x"7a", x"7d", x"78", x"74", x"73", x"77", x"7b", x"7f", x"80", x"7f", x"7e", x"7d", 
        x"79", x"7a", x"7c", x"99", x"cf", x"b7", x"99", x"96", x"92", x"96", x"9b", x"95", x"8b", x"8c", x"95", 
        x"98", x"8c", x"83", x"87", x"8f", x"8c", x"82", x"7e", x"86", x"8c", x"8c", x"b5", x"ef", x"f5", x"f3", 
        x"f2", x"f2", x"f2", x"f4", x"f5", x"f6", x"f6", x"f4", x"f2", x"f0", x"f2", x"f3", x"f2", x"f3", x"f2", 
        x"f1", x"ec", x"de", x"c8", x"b5", x"b9", x"bb", x"b9", x"bb", x"ba", x"bd", x"a4", x"71", x"65", x"62", 
        x"58", x"53", x"54", x"56", x"51", x"4b", x"3d", x"15", x"07", x"09", x"13", x"14", x"0f", x"10", x"0e", 
        x"0e", x"0e", x"26", x"3c", x"37", x"3a", x"37", x"3a", x"41", x"39", x"42", x"57", x"64", x"6d", x"6a", 
        x"6b", x"69", x"6e", x"6f", x"71", x"70", x"69", x"69", x"69", x"66", x"70", x"5c", x"1a", x"0b", x"30", 
        x"56", x"58", x"4a", x"3d", x"38", x"3a", x"44", x"53", x"3b", x"26", x"1a", x"1a", x"0a", x"0b", x"0b", 
        x"08", x"0c", x"18", x"19", x"14", x"17", x"19", x"1c", x"1b", x"18", x"17", x"1a", x"1e", x"13", x"07", 
        x"07", x"0a", x"13", x"13", x"12", x"13", x"15", x"18", x"19", x"14", x"0f", x"11", x"17", x"0f", x"07", 
        x"1d", x"3b", x"19", x"1b", x"1c", x"19", x"13", x"14", x"13", x"11", x"0d", x"0b", x"0d", x"0d", x"08", 
        x"0e", x"1c", x"15", x"18", x"13", x"0c", x"0f", x"45", x"86", x"8b", x"89", x"8d", x"8b", x"7f", x"79", 
        x"75", x"72", x"66", x"32", x"25", x"1f", x"0e", x"0b", x"0a", x"0a", x"0b", x"11", x"48", x"51", x"52", 
        x"51", x"58", x"62", x"5f", x"5d", x"66", x"54", x"2c", x"2e", x"33", x"39", x"2d", x"16", x"09", x"0f", 
        x"2f", x"3b", x"5a", x"6e", x"58", x"75", x"41", x"48", x"7b", x"5e", x"3a", x"2b", x"32", x"36", x"26", 
        x"25", x"2f", x"2c", x"40", x"46", x"38", x"47", x"3a", x"2b", x"28", x"45", x"6a", x"2f", x"17", x"1c", 
        x"24", x"3b", x"38", x"23", x"21", x"29", x"59", x"4e", x"52", x"35", x"38", x"3f", x"4f", x"7d", x"45", 
        x"70", x"74", x"8c", x"72", x"64", x"56", x"5b", x"65", x"56", x"46", x"50", x"73", x"3d", x"28", x"5f", 
        x"77", x"7c", x"72", x"74", x"80", x"69", x"40", x"38", x"42", x"50", x"3b", x"3a", x"4d", x"49", x"68", 
        x"65", x"76", x"59", x"59", x"6b", x"81", x"7b", x"5b", x"45", x"6d", x"7b", x"86", x"a5", x"b0", x"9a", 
        x"93", x"8e", x"98", x"9c", x"81", x"79", x"89", x"5d", x"6b", x"55", x"5b", x"79", x"7a", x"81", x"6c", 
        x"57", x"63", x"6e", x"5b", x"4f", x"85", x"92", x"81", x"83", x"8a", x"85", x"90", x"a1", x"99", x"87", 
        x"90", x"b4", x"a5", x"a9", x"bc", x"9e", x"b2", x"98", x"3c", x"42", x"6f", x"70", x"71", x"a6", x"b7", 
        x"9a", x"97", x"9c", x"9d", x"87", x"95", x"9f", x"96", x"a3", x"74", x"57", x"61", x"55", x"9a", x"82", 
        x"78", x"78", x"70", x"a4", x"df", x"d6", x"d6", x"d8", x"d2", x"d8", x"dc", x"cd", x"cf", x"cf", x"cf", 
        x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d1", x"d0", x"d0", x"d2", x"d2", x"d1", x"d1", 
        x"d5", x"d5", x"d2", x"d1", x"d2", x"d2", x"d1", x"d3", x"d4", x"d4", x"d2", x"d1", x"d1", x"d1", x"d0", 
        x"d0", x"d0", x"d1", x"d2", x"d4", x"d4", x"d4", x"d4", x"d1", x"cf", x"cd", x"dd", x"db", x"a6", x"92", 
        x"7d", x"76", x"6d", x"64", x"6a", x"9c", x"9c", x"6e", x"74", x"82", x"84", x"87", x"8c", x"8f", x"8e", 
        x"8e", x"8c", x"8c", x"8e", x"95", x"94", x"8a", x"85", x"84", x"94", x"9b", x"90", x"92", x"8d", x"87", 
        x"7a", x"73", x"75", x"80", x"82", x"7b", x"77", x"71", x"6b", x"68", x"6b", x"6c", x"6d", x"6e", x"66", 
        x"5d", x"59", x"5c", x"66", x"98", x"e0", x"b4", x"7d", x"85", x"91", x"95", x"8f", x"8c", x"8b", x"8f", 
        x"97", x"9a", x"9a", x"9a", x"8e", x"8a", x"92", x"95", x"93", x"91", x"8c", x"80", x"7d", x"86", x"8c", 
        x"8e", x"8b", x"80", x"78", x"77", x"7a", x"7e", x"7f", x"80", x"7b", x"71", x"73", x"7c", x"86", x"8e", 
        x"b6", x"e0", x"a4", x"8c", x"93", x"97", x"9a", x"9b", x"9a", x"99", x"9a", x"a3", x"a8", x"a6", x"a1", 
        x"9f", x"95", x"91", x"94", x"94", x"93", x"95", x"93", x"8a", x"8a", x"8c", x"8a", x"88", x"85", x"81", 
        x"7f", x"81", x"83", x"84", x"85", x"84", x"84", x"86", x"a6", x"d9", x"98", x"6e", x"7f", x"85", x"82", 
        x"77", x"76", x"7d", x"87", x"8e", x"8e", x"8b", x"7d", x"7d", x"7d", x"7f", x"84", x"81", x"77", x"6d", 
        x"6f", x"74", x"7a", x"7d", x"7f", x"7f", x"71", x"65", x"67", x"6e", x"6e", x"6e", x"6c", x"89", x"cc", 
        x"d4", x"c6", x"ca", x"c6", x"c1", x"be", x"c0", x"c8", x"ce", x"c8", x"c1", x"bd", x"b9", x"b7", x"be", 
        x"bd", x"b8", x"bb", x"c0", x"c2", x"c0", x"ba", x"b3", x"b6", x"bb", x"ba", x"bd", x"c0", x"bf", x"c0", 
        x"c1", x"c7", x"d6", x"98", x"8e", x"94", x"8e", x"8c", x"8e", x"92", x"99", x"99", x"91", x"8e", x"8f", 
        x"90", x"8d", x"8b", x"8a", x"86", x"85", x"81", x"84", x"80", x"76", x"76", x"76", x"7b", x"83", x"87", 
        x"91", x"cf", x"c9", x"8b", x"88", x"8b", x"8b", x"8e", x"8e", x"8d", x"89", x"87", x"85", x"80", x"80", 
        x"83", x"85", x"87", x"89", x"87", x"7e", x"7b", x"7c", x"7f", x"85", x"8a", x"88", x"86", x"a7", x"e0", 
        x"a4", x"97", x"95", x"a0", x"95", x"97", x"93", x"97", x"96", x"99", x"98", x"9b", x"93", x"98", x"92", 
        x"89", x"7d", x"75", x"72", x"72", x"74", x"72", x"70", x"75", x"98", x"db", x"97", x"78", x"78", x"79", 
        x"7a", x"79", x"75", x"75", x"77", x"78", x"79", x"79", x"7a", x"7c", x"7d", x"7c", x"7a", x"79", x"79", 
        x"7c", x"78", x"74", x"92", x"cd", x"b8", x"95", x"9b", x"97", x"91", x"94", x"99", x"98", x"8f", x"90", 
        x"98", x"98", x"8d", x"82", x"82", x"8f", x"92", x"86", x"81", x"87", x"8d", x"b5", x"ec", x"f2", x"f1", 
        x"f1", x"f0", x"f1", x"f2", x"f3", x"f4", x"f5", x"f4", x"f1", x"ef", x"ef", x"f1", x"f1", x"f0", x"f1", 
        x"ee", x"eb", x"df", x"cb", x"ba", x"ba", x"bb", x"b8", x"be", x"bf", x"bf", x"b6", x"88", x"63", x"62", 
        x"63", x"5c", x"58", x"52", x"4e", x"4a", x"3f", x"17", x"06", x"08", x"12", x"13", x"11", x"14", x"16", 
        x"10", x"12", x"32", x"43", x"3d", x"43", x"42", x"43", x"48", x"3c", x"42", x"57", x"66", x"70", x"6c", 
        x"6d", x"6a", x"6d", x"70", x"70", x"6f", x"6b", x"67", x"67", x"67", x"6d", x"5d", x"23", x"0b", x"1f", 
        x"38", x"39", x"3a", x"41", x"41", x"3e", x"39", x"3c", x"24", x"17", x"18", x"19", x"08", x"0c", x"0d", 
        x"08", x"0b", x"14", x"16", x"14", x"19", x"19", x"1c", x"1c", x"1a", x"19", x"1a", x"1b", x"10", x"06", 
        x"06", x"09", x"13", x"13", x"12", x"14", x"15", x"16", x"16", x"14", x"11", x"12", x"12", x"09", x"04", 
        x"19", x"3d", x"1f", x"1f", x"1d", x"1b", x"16", x"15", x"14", x"13", x"0f", x"0c", x"0c", x"0d", x"0a", 
        x"0b", x"19", x"14", x"17", x"13", x"0d", x"10", x"43", x"86", x"8b", x"88", x"8c", x"8d", x"85", x"7e", 
        x"72", x"6f", x"6a", x"34", x"22", x"1c", x"09", x"02", x"03", x"03", x"03", x"08", x"43", x"50", x"4f", 
        x"4e", x"53", x"5d", x"58", x"55", x"5a", x"46", x"18", x"19", x"1f", x"25", x"1f", x"0f", x"07", x"0b", 
        x"36", x"3e", x"49", x"5e", x"56", x"46", x"49", x"6b", x"69", x"42", x"67", x"62", x"41", x"36", x"1d", 
        x"1f", x"21", x"10", x"1f", x"37", x"3e", x"3a", x"3f", x"2e", x"1a", x"1d", x"3f", x"2f", x"1a", x"21", 
        x"37", x"49", x"3a", x"20", x"24", x"27", x"48", x"4d", x"63", x"41", x"31", x"2f", x"2c", x"45", x"56", 
        x"4b", x"5f", x"8e", x"7d", x"6b", x"44", x"4f", x"51", x"65", x"3b", x"4e", x"63", x"57", x"4e", x"76", 
        x"82", x"53", x"65", x"72", x"78", x"5d", x"2b", x"2f", x"49", x"61", x"4c", x"37", x"27", x"39", x"56", 
        x"5c", x"75", x"64", x"82", x"79", x"5b", x"5e", x"73", x"6c", x"78", x"77", x"94", x"a9", x"ab", x"a0", 
        x"a1", x"9d", x"ae", x"99", x"95", x"9a", x"93", x"7a", x"70", x"a0", x"ae", x"a2", x"98", x"a1", x"74", 
        x"49", x"6f", x"73", x"5a", x"54", x"84", x"93", x"84", x"8b", x"94", x"8c", x"8f", x"98", x"8e", x"83", 
        x"a1", x"c1", x"a4", x"a1", x"aa", x"9c", x"bb", x"9c", x"3c", x"40", x"70", x"6f", x"70", x"ad", x"bb", 
        x"9b", x"90", x"90", x"97", x"85", x"95", x"a6", x"93", x"a7", x"7a", x"54", x"60", x"53", x"95", x"80", 
        x"7a", x"7a", x"72", x"a4", x"de", x"d6", x"d5", x"d8", x"d3", x"da", x"dd", x"cc", x"cf", x"d0", x"d0", 
        x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d2", x"d1", x"d1", x"d3", x"d2", x"d1", x"d2", 
        x"d4", x"d4", x"d2", x"d1", x"d2", x"d3", x"d2", x"d3", x"d5", x"d5", x"d4", x"d2", x"d1", x"d1", x"d0", 
        x"d0", x"d0", x"d1", x"d2", x"d3", x"d4", x"d4", x"d6", x"d5", x"d4", x"d2", x"e0", x"db", x"a3", x"86", 
        x"6e", x"72", x"75", x"7a", x"83", x"a3", x"a3", x"86", x"90", x"96", x"92", x"96", x"97", x"90", x"8d", 
        x"91", x"95", x"95", x"8f", x"89", x"77", x"66", x"6d", x"6f", x"75", x"7d", x"6d", x"5d", x"5b", x"5c", 
        x"5a", x"5f", x"67", x"70", x"70", x"6a", x"69", x"6a", x"6c", x"6d", x"6f", x"78", x"7c", x"79", x"78", 
        x"77", x"7a", x"80", x"81", x"a0", x"e2", x"bb", x"89", x"8e", x"91", x"91", x"8c", x"82", x"7c", x"7e", 
        x"82", x"83", x"81", x"7a", x"70", x"6f", x"7b", x"81", x"81", x"82", x"7c", x"77", x"7e", x"8a", x"90", 
        x"92", x"8f", x"88", x"84", x"88", x"90", x"98", x"9c", x"9d", x"9c", x"93", x"8c", x"8d", x"96", x"97", 
        x"b6", x"df", x"aa", x"8a", x"8d", x"92", x"97", x"96", x"94", x"8f", x"86", x"83", x"84", x"84", x"82", 
        x"83", x"80", x"80", x"87", x"8e", x"90", x"90", x"8c", x"8b", x"8c", x"8e", x"92", x"95", x"97", x"98", 
        x"95", x"95", x"9d", x"a4", x"a7", x"a6", x"a2", x"98", x"ac", x"e2", x"a5", x"73", x"77", x"7c", x"7f", 
        x"77", x"6d", x"69", x"6b", x"6f", x"71", x"71", x"6b", x"63", x"60", x"66", x"71", x"75", x"72", x"70", 
        x"6d", x"6a", x"6f", x"76", x"7f", x"88", x"80", x"76", x"72", x"79", x"7f", x"84", x"83", x"97", x"d1", 
        x"d4", x"bc", x"ba", x"bf", x"c5", x"c2", x"ba", x"ba", x"bc", x"ba", x"b9", x"b9", x"b4", x"b2", x"ba", 
        x"bd", x"be", x"c0", x"bf", x"bb", x"c4", x"c5", x"c0", x"bf", x"c2", x"c4", x"c5", x"c9", x"c9", x"c3", 
        x"bd", x"c3", x"db", x"a0", x"8d", x"8b", x"87", x"88", x"8f", x"93", x"90", x"89", x"83", x"83", x"8b", 
        x"93", x"8f", x"89", x"87", x"8b", x"92", x"93", x"91", x"88", x"7f", x"85", x"8d", x"98", x"9f", x"98", 
        x"96", x"ce", x"cb", x"89", x"85", x"86", x"83", x"80", x"7f", x"7f", x"7b", x"7a", x"79", x"75", x"75", 
        x"7a", x"7e", x"84", x"8b", x"8a", x"82", x"80", x"7f", x"7e", x"83", x"89", x"8b", x"89", x"a6", x"e0", 
        x"a6", x"95", x"91", x"9a", x"8e", x"91", x"8f", x"93", x"94", x"94", x"95", x"99", x"91", x"96", x"94", 
        x"8d", x"7d", x"78", x"77", x"78", x"79", x"77", x"70", x"70", x"92", x"d7", x"99", x"79", x"78", x"79", 
        x"7d", x"7e", x"79", x"75", x"73", x"75", x"76", x"77", x"7b", x"7d", x"7d", x"7c", x"7c", x"7c", x"7e", 
        x"81", x"7f", x"7a", x"8f", x"ca", x"b8", x"93", x"9c", x"9d", x"94", x"8b", x"91", x"9c", x"9a", x"8e", 
        x"89", x"90", x"95", x"8f", x"83", x"7f", x"87", x"8d", x"86", x"83", x"84", x"ae", x"ea", x"f4", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f4", x"f3", x"f2", x"f1", x"ef", x"ed", x"ee", x"f1", x"ef", x"f0", 
        x"ef", x"eb", x"de", x"c9", x"b9", x"b8", x"ba", x"b6", x"bd", x"bf", x"b6", x"b7", x"ac", x"79", x"5e", 
        x"5b", x"57", x"58", x"55", x"5a", x"56", x"4c", x"1d", x"05", x"07", x"17", x"1a", x"16", x"15", x"13", 
        x"0e", x"1c", x"3d", x"46", x"41", x"3e", x"38", x"38", x"41", x"38", x"3d", x"56", x"65", x"6f", x"6b", 
        x"6d", x"6a", x"6b", x"71", x"70", x"70", x"6e", x"68", x"67", x"69", x"70", x"63", x"25", x"0d", x"25", 
        x"3a", x"37", x"36", x"36", x"37", x"35", x"32", x"36", x"23", x"16", x"19", x"18", x"09", x"0b", x"0d", 
        x"08", x"08", x"11", x"17", x"18", x"1d", x"1c", x"1e", x"1f", x"1d", x"1a", x"1a", x"1a", x"10", x"06", 
        x"05", x"09", x"12", x"14", x"13", x"14", x"14", x"14", x"13", x"12", x"13", x"11", x"0d", x"08", x"07", 
        x"17", x"35", x"1b", x"1a", x"16", x"15", x"13", x"12", x"12", x"11", x"0e", x"08", x"07", x"08", x"09", 
        x"07", x"16", x"12", x"15", x"10", x"0d", x"10", x"41", x"87", x"8c", x"88", x"8a", x"8d", x"8a", x"86", 
        x"79", x"6f", x"6b", x"3d", x"2a", x"21", x"0b", x"03", x"04", x"04", x"04", x"08", x"45", x"55", x"53", 
        x"52", x"54", x"5d", x"5a", x"57", x"5c", x"4e", x"1e", x"1d", x"20", x"22", x"20", x"12", x"07", x"09", 
        x"7b", x"8c", x"54", x"40", x"62", x"58", x"51", x"6d", x"6d", x"62", x"42", x"33", x"32", x"53", x"3f", 
        x"30", x"1d", x"20", x"20", x"49", x"91", x"7a", x"69", x"4d", x"32", x"2a", x"27", x"4d", x"6d", x"5d", 
        x"51", x"4f", x"54", x"35", x"3b", x"31", x"30", x"4a", x"75", x"6f", x"43", x"3a", x"38", x"36", x"76", 
        x"32", x"44", x"7d", x"85", x"65", x"6e", x"6d", x"42", x"2b", x"35", x"67", x"5e", x"64", x"85", x"83", 
        x"5f", x"41", x"4e", x"4f", x"7f", x"5a", x"41", x"59", x"3d", x"2b", x"3d", x"3a", x"45", x"50", x"64", 
        x"58", x"71", x"88", x"8b", x"54", x"6b", x"64", x"5e", x"65", x"67", x"67", x"82", x"a1", x"aa", x"bc", 
        x"a4", x"93", x"a3", x"87", x"84", x"90", x"7e", x"8e", x"89", x"91", x"d8", x"bc", x"9f", x"bb", x"83", 
        x"45", x"92", x"98", x"8d", x"5b", x"83", x"98", x"94", x"93", x"94", x"95", x"9c", x"8e", x"86", x"7e", 
        x"8f", x"98", x"8e", x"aa", x"bf", x"9c", x"af", x"94", x"38", x"3a", x"6e", x"6d", x"70", x"b0", x"b5", 
        x"91", x"93", x"98", x"9e", x"8c", x"9c", x"b2", x"8c", x"9f", x"76", x"4f", x"60", x"52", x"94", x"85", 
        x"7f", x"79", x"72", x"a3", x"db", x"d3", x"d3", x"d4", x"d4", x"dc", x"df", x"cd", x"cf", x"d0", x"d2", 
        x"d2", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d2", x"d2", x"d3", x"d3", x"d4", x"d3", x"d2", x"d2", 
        x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", x"d3", x"d5", x"d6", x"d6", x"d4", x"d2", x"d1", x"d1", x"d3", 
        x"d4", x"d3", x"d3", x"d3", x"d4", x"d5", x"d7", x"d7", x"d3", x"d0", x"cd", x"dc", x"da", x"a3", x"93", 
        x"81", x"78", x"6b", x"61", x"6b", x"a0", x"9f", x"71", x"70", x"75", x"71", x"77", x"83", x"88", x"87", 
        x"87", x"87", x"89", x"87", x"88", x"81", x"70", x"7a", x"81", x"87", x"8f", x"85", x"7d", x"7f", x"81", 
        x"80", x"82", x"89", x"92", x"86", x"7a", x"77", x"77", x"7a", x"7b", x"7c", x"75", x"6a", x"64", x"65", 
        x"67", x"67", x"69", x"6e", x"98", x"e0", x"b6", x"7e", x"84", x"88", x"85", x"81", x"7a", x"7c", x"87", 
        x"90", x"93", x"92", x"8d", x"8a", x"8f", x"9d", x"a3", x"a1", x"9d", x"95", x"89", x"85", x"8b", x"90", 
        x"93", x"8f", x"88", x"80", x"7c", x"80", x"86", x"87", x"83", x"7e", x"73", x"69", x"68", x"77", x"84", 
        x"af", x"de", x"a2", x"84", x"8a", x"91", x"95", x"95", x"96", x"95", x"90", x"91", x"98", x"9e", x"a0", 
        x"a1", x"a1", x"9b", x"96", x"95", x"98", x"99", x"97", x"94", x"90", x"8e", x"8f", x"93", x"95", x"96", 
        x"93", x"8c", x"84", x"7f", x"80", x"80", x"7f", x"7e", x"9d", x"d8", x"9d", x"5f", x"5b", x"6d", x"7c", 
        x"76", x"70", x"6c", x"69", x"69", x"71", x"7a", x"7d", x"7d", x"7c", x"7a", x"78", x"7d", x"85", x"85", 
        x"81", x"7c", x"7a", x"79", x"7d", x"86", x"82", x"78", x"6e", x"6a", x"67", x"65", x"64", x"8a", x"d2", 
        x"d3", x"ba", x"b4", x"b3", x"bc", x"c3", x"c4", x"c0", x"bd", x"b8", x"bd", x"c4", x"c4", x"c2", x"c5", 
        x"c6", x"c8", x"cd", x"cd", x"c3", x"bd", x"be", x"bc", x"bb", x"c0", x"c1", x"bc", x"bb", x"bc", x"bc", 
        x"b8", x"be", x"d5", x"95", x"7b", x"7e", x"82", x"84", x"87", x"87", x"85", x"84", x"84", x"87", x"8f", 
        x"93", x"90", x"8c", x"8c", x"8f", x"93", x"90", x"8a", x"84", x"7f", x"84", x"8b", x"90", x"8f", x"85", 
        x"86", x"c4", x"c7", x"7b", x"73", x"77", x"79", x"7d", x"7f", x"80", x"81", x"81", x"7c", x"78", x"7a", 
        x"7f", x"81", x"87", x"8e", x"89", x"7f", x"7b", x"79", x"7a", x"7f", x"83", x"85", x"85", x"9f", x"db", 
        x"a7", x"93", x"90", x"98", x"8e", x"90", x"91", x"95", x"96", x"94", x"94", x"97", x"90", x"98", x"99", 
        x"8f", x"7a", x"76", x"73", x"71", x"73", x"72", x"6c", x"6a", x"8c", x"d3", x"9a", x"76", x"73", x"71", 
        x"74", x"77", x"7b", x"7b", x"79", x"7a", x"79", x"79", x"80", x"81", x"81", x"7f", x"7b", x"79", x"78", 
        x"7f", x"81", x"7e", x"90", x"cb", x"b9", x"8e", x"8f", x"9b", x"9d", x"8f", x"86", x"8b", x"98", x"98", 
        x"8b", x"7e", x"81", x"8e", x"91", x"83", x"80", x"8e", x"91", x"8b", x"81", x"a6", x"e7", x"f6", x"f4", 
        x"f4", x"f5", x"f5", x"f4", x"f4", x"f3", x"f3", x"f1", x"f1", x"f1", x"ef", x"ef", x"f1", x"f1", x"f2", 
        x"f0", x"eb", x"de", x"cc", x"be", x"bf", x"c0", x"b7", x"b6", x"b7", x"b5", x"bc", x"b9", x"8e", x"69", 
        x"60", x"64", x"62", x"5c", x"5c", x"55", x"4b", x"20", x"05", x"04", x"13", x"17", x"12", x"13", x"12", 
        x"17", x"31", x"44", x"42", x"40", x"3c", x"38", x"3b", x"46", x"3e", x"3e", x"57", x"64", x"6e", x"6b", 
        x"6c", x"69", x"68", x"6e", x"72", x"72", x"6f", x"6a", x"6a", x"69", x"6e", x"62", x"23", x"0a", x"20", 
        x"3a", x"39", x"38", x"3c", x"38", x"35", x"33", x"39", x"2d", x"1f", x"1e", x"1b", x"0a", x"09", x"0b", 
        x"06", x"05", x"11", x"1d", x"1f", x"20", x"1d", x"1e", x"20", x"1d", x"1a", x"1a", x"1b", x"12", x"07", 
        x"06", x"08", x"11", x"13", x"11", x"12", x"12", x"13", x"12", x"13", x"12", x"0d", x"08", x"09", x"0b", 
        x"17", x"32", x"1e", x"1b", x"15", x"15", x"15", x"15", x"17", x"17", x"13", x"0b", x"06", x"05", x"06", 
        x"07", x"19", x"14", x"15", x"10", x"0e", x"10", x"3f", x"8a", x"8f", x"89", x"8a", x"8a", x"85", x"84", 
        x"7f", x"73", x"6c", x"3f", x"2b", x"1f", x"09", x"04", x"05", x"03", x"02", x"05", x"42", x"55", x"4e", 
        x"4e", x"51", x"5b", x"5c", x"5a", x"5d", x"54", x"23", x"21", x"22", x"20", x"1d", x"0f", x"07", x"07", 
        x"58", x"70", x"52", x"31", x"4e", x"62", x"57", x"70", x"7f", x"4f", x"2c", x"35", x"50", x"35", x"32", 
        x"32", x"2e", x"3c", x"37", x"32", x"50", x"48", x"4b", x"6d", x"73", x"3e", x"38", x"60", x"87", x"73", 
        x"43", x"39", x"33", x"28", x"3d", x"55", x"29", x"35", x"5b", x"59", x"43", x"3a", x"32", x"26", x"73", 
        x"70", x"69", x"76", x"7e", x"7d", x"8c", x"59", x"2f", x"1e", x"3e", x"5c", x"5e", x"58", x"6e", x"71", 
        x"57", x"43", x"3b", x"5a", x"7e", x"4d", x"3c", x"58", x"48", x"3e", x"38", x"40", x"57", x"41", x"4d", 
        x"54", x"60", x"81", x"77", x"5b", x"5b", x"6d", x"6e", x"6c", x"68", x"70", x"98", x"b0", x"a8", x"a7", 
        x"9f", x"ac", x"ce", x"be", x"98", x"a9", x"8b", x"94", x"b6", x"99", x"b2", x"b9", x"8f", x"a8", x"7c", 
        x"46", x"7d", x"b1", x"a6", x"51", x"7f", x"97", x"98", x"90", x"95", x"b6", x"c6", x"bb", x"a0", x"8e", 
        x"ab", x"c0", x"bd", x"b9", x"b5", x"8d", x"9a", x"91", x"3d", x"3b", x"6a", x"71", x"70", x"a0", x"a2", 
        x"8c", x"8b", x"91", x"9b", x"87", x"86", x"98", x"89", x"9e", x"73", x"55", x"67", x"55", x"97", x"88", 
        x"7f", x"7b", x"74", x"a4", x"db", x"d3", x"d4", x"d4", x"d4", x"dc", x"de", x"cd", x"cf", x"d0", x"d1", 
        x"d1", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", x"d2", x"d3", x"d3", x"d3", x"d2", x"d2", x"d3", 
        x"d3", x"d2", x"d2", x"d3", x"d2", x"d3", x"d4", x"d6", x"d6", x"d4", x"d2", x"d1", x"d2", x"d3", x"d5", 
        x"d5", x"d3", x"d2", x"d2", x"d1", x"d2", x"d5", x"d5", x"d4", x"d4", x"d2", x"e0", x"de", x"a5", x"88", 
        x"70", x"6f", x"6f", x"74", x"83", x"aa", x"ad", x"8d", x"89", x"8a", x"8b", x"90", x"92", x"93", x"94", 
        x"8e", x"85", x"83", x"85", x"8a", x"88", x"7a", x"7a", x"7c", x"78", x"72", x"67", x"62", x"6a", x"6f", 
        x"70", x"6e", x"73", x"7e", x"72", x"6a", x"6c", x"71", x"75", x"75", x"73", x"72", x"6e", x"6f", x"77", 
        x"80", x"83", x"83", x"7f", x"9a", x"e0", x"c0", x"90", x"92", x"91", x"8c", x"86", x"83", x"87", x"90", 
        x"92", x"8f", x"89", x"7b", x"79", x"7a", x"7e", x"81", x"82", x"7e", x"78", x"75", x"7b", x"85", x"8b", 
        x"8f", x"8d", x"89", x"82", x"7e", x"85", x"91", x"97", x"94", x"92", x"8e", x"88", x"88", x"93", x"97", 
        x"b8", x"e7", x"b3", x"94", x"95", x"95", x"93", x"92", x"93", x"93", x"92", x"92", x"91", x"90", x"8d", 
        x"8c", x"8c", x"88", x"83", x"84", x"8a", x"8c", x"8d", x"90", x"8f", x"8e", x"91", x"96", x"99", x"97", 
        x"94", x"91", x"8f", x"8f", x"93", x"98", x"9b", x"9a", x"af", x"e2", x"af", x"7c", x"78", x"79", x"7c", 
        x"78", x"78", x"78", x"74", x"6e", x"6f", x"73", x"71", x"74", x"77", x"74", x"6a", x"67", x"6c", x"6c", 
        x"6c", x"6c", x"72", x"71", x"71", x"76", x"76", x"75", x"77", x"7a", x"7a", x"73", x"6c", x"86", x"c7", 
        x"d4", x"c9", x"cc", x"ca", x"c9", x"c6", x"c2", x"c8", x"c9", x"c1", x"be", x"bf", x"bb", x"be", x"c6", 
        x"c4", x"bb", x"b7", x"b8", x"b7", x"b5", x"bb", x"be", x"ba", x"bc", x"c2", x"c1", x"c3", x"c2", x"c1", 
        x"c0", x"c6", x"da", x"9d", x"8a", x"91", x"91", x"91", x"8d", x"8a", x"8a", x"8e", x"90", x"89", x"84", 
        x"82", x"83", x"86", x"88", x"8a", x"86", x"7e", x"7c", x"7e", x"80", x"83", x"87", x"86", x"84", x"7f", 
        x"87", x"c3", x"c8", x"80", x"78", x"7b", x"7a", x"7c", x"7f", x"81", x"83", x"81", x"7c", x"76", x"77", 
        x"7c", x"7e", x"81", x"84", x"7e", x"76", x"74", x"74", x"76", x"7f", x"87", x"86", x"87", x"9e", x"d8", 
        x"aa", x"95", x"90", x"99", x"91", x"96", x"98", x"9d", x"9c", x"9d", x"9a", x"99", x"94", x"9a", x"9b", 
        x"8e", x"7e", x"7c", x"75", x"70", x"72", x"74", x"72", x"6e", x"8d", x"d5", x"a0", x"7a", x"77", x"77", 
        x"7a", x"7d", x"7f", x"7c", x"79", x"79", x"7a", x"7c", x"7e", x"7d", x"7e", x"7f", x"7f", x"7d", x"7b", 
        x"7d", x"7e", x"7b", x"90", x"d1", x"c5", x"94", x"89", x"8d", x"97", x"96", x"8b", x"84", x"8a", x"93", 
        x"97", x"8e", x"85", x"88", x"92", x"8e", x"85", x"82", x"89", x"8e", x"90", x"b0", x"e7", x"f4", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f4", x"f0", x"f0", x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f0", x"ec", x"de", x"cb", x"bc", x"b9", x"b7", x"b6", x"b8", x"b8", x"b5", x"b5", x"b9", x"ab", x"80", 
        x"5e", x"5e", x"5d", x"5c", x"5e", x"5c", x"4e", x"24", x"08", x"04", x"15", x"1b", x"1c", x"1c", x"15", 
        x"21", x"3b", x"42", x"40", x"42", x"42", x"3f", x"3e", x"41", x"36", x"37", x"57", x"65", x"6f", x"6d", 
        x"6d", x"6b", x"6a", x"6b", x"72", x"73", x"6d", x"6d", x"6b", x"67", x"6b", x"61", x"28", x"0c", x"1f", 
        x"3f", x"41", x"38", x"35", x"36", x"38", x"3a", x"3f", x"30", x"1e", x"1c", x"19", x"0c", x"09", x"0c", 
        x"07", x"05", x"10", x"20", x"20", x"20", x"1d", x"1d", x"21", x"1e", x"1c", x"1a", x"1a", x"13", x"08", 
        x"07", x"0a", x"13", x"15", x"10", x"0f", x"10", x"11", x"12", x"14", x"0e", x"07", x"04", x"09", x"09", 
        x"11", x"31", x"1f", x"1a", x"14", x"13", x"12", x"12", x"0f", x"0e", x"0d", x"0a", x"07", x"08", x"0b", 
        x"0b", x"1d", x"17", x"14", x"0e", x"0d", x"0e", x"3a", x"88", x"8f", x"8b", x"8f", x"8f", x"87", x"80", 
        x"7d", x"79", x"71", x"3e", x"26", x"1d", x"09", x"04", x"04", x"02", x"02", x"04", x"40", x"56", x"4f", 
        x"4f", x"51", x"5a", x"5b", x"58", x"58", x"54", x"22", x"1e", x"1f", x"1f", x"1d", x"11", x"09", x"08", 
        x"32", x"60", x"57", x"36", x"2d", x"3a", x"4a", x"65", x"6a", x"3a", x"65", x"5a", x"52", x"35", x"3b", 
        x"2d", x"2e", x"30", x"29", x"30", x"27", x"27", x"34", x"47", x"65", x"56", x"54", x"28", x"30", x"3d", 
        x"56", x"4c", x"17", x"1d", x"36", x"6d", x"42", x"4f", x"65", x"43", x"39", x"35", x"2c", x"24", x"51", 
        x"66", x"76", x"a0", x"a5", x"8a", x"86", x"4b", x"27", x"2b", x"37", x"57", x"76", x"5f", x"4a", x"47", 
        x"51", x"4e", x"5b", x"7e", x"76", x"37", x"31", x"43", x"57", x"54", x"40", x"50", x"54", x"47", x"62", 
        x"74", x"78", x"6d", x"58", x"66", x"5c", x"67", x"6b", x"6b", x"73", x"5c", x"6c", x"95", x"8b", x"a2", 
        x"b5", x"b1", x"d0", x"dc", x"a8", x"9a", x"bf", x"bb", x"be", x"99", x"90", x"a3", x"a8", x"af", x"70", 
        x"48", x"8d", x"c0", x"81", x"4c", x"8b", x"94", x"88", x"8b", x"a3", x"bf", x"c1", x"af", x"96", x"97", 
        x"bd", x"c9", x"c3", x"b3", x"9f", x"9a", x"a5", x"9c", x"3b", x"3b", x"6e", x"72", x"6b", x"9c", x"af", 
        x"ac", x"a3", x"9e", x"9f", x"8d", x"82", x"8c", x"8d", x"99", x"70", x"56", x"66", x"52", x"97", x"86", 
        x"7c", x"7d", x"76", x"a6", x"db", x"d4", x"d6", x"d6", x"d3", x"da", x"dd", x"cd", x"cf", x"cf", x"d0", 
        x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d0", x"d1", x"d2", x"d3", x"d3", x"d2", x"d2", x"d2", x"d3", 
        x"d2", x"d1", x"d2", x"d3", x"d2", x"d3", x"d5", x"d5", x"d5", x"d3", x"d1", x"d1", x"d2", x"d3", x"d3", 
        x"d3", x"d2", x"d1", x"d1", x"d0", x"d1", x"d3", x"d3", x"d3", x"d4", x"d1", x"de", x"dc", x"a1", x"8d", 
        x"7a", x"73", x"6b", x"64", x"6e", x"a2", x"a6", x"77", x"6f", x"79", x"83", x"8b", x"8d", x"8c", x"86", 
        x"80", x"7f", x"88", x"8d", x"90", x"94", x"91", x"8d", x"8f", x"8c", x"86", x"80", x"81", x"88", x"8a", 
        x"86", x"7c", x"7e", x"86", x"7f", x"7a", x"7f", x"81", x"80", x"7a", x"75", x"70", x"6c", x"6e", x"74", 
        x"79", x"79", x"74", x"73", x"96", x"de", x"be", x"89", x"87", x"84", x"7c", x"78", x"7c", x"83", x"8a", 
        x"8d", x"8b", x"85", x"7e", x"86", x"8f", x"96", x"98", x"97", x"92", x"8d", x"8c", x"90", x"94", x"94", 
        x"95", x"93", x"8d", x"86", x"83", x"89", x"93", x"98", x"97", x"92", x"88", x"7e", x"75", x"7d", x"84", 
        x"ae", x"e1", x"a2", x"80", x"80", x"85", x"8b", x"8d", x"8d", x"8c", x"8b", x"8c", x"8e", x"92", x"95", 
        x"96", x"94", x"95", x"94", x"98", x"9e", x"9f", x"a1", x"a2", x"9f", x"9b", x"98", x"96", x"95", x"93", 
        x"91", x"91", x"93", x"93", x"91", x"91", x"94", x"93", x"a5", x"dc", x"af", x"7a", x"70", x"69", x"66", 
        x"66", x"69", x"70", x"75", x"76", x"74", x"74", x"73", x"72", x"75", x"79", x"79", x"7a", x"7c", x"76", 
        x"71", x"71", x"7a", x"7f", x"83", x"8b", x"86", x"7f", x"78", x"77", x"79", x"76", x"72", x"8d", x"ce", 
        x"d6", x"c0", x"c1", x"c5", x"c6", x"be", x"b7", x"b9", x"ba", x"b8", x"be", x"c1", x"ba", x"b5", x"bb", 
        x"bb", x"b8", x"bb", x"be", x"bb", x"ba", x"c3", x"cb", x"c7", x"c5", x"c8", x"c4", x"c4", x"c5", x"c3", 
        x"be", x"c5", x"db", x"9b", x"86", x"8b", x"85", x"82", x"7e", x"7b", x"81", x"86", x"81", x"7d", x"7d", 
        x"82", x"88", x"8d", x"8f", x"8c", x"87", x"82", x"83", x"8a", x"90", x"90", x"8b", x"84", x"80", x"7e", 
        x"87", x"c2", x"cb", x"83", x"7a", x"7c", x"79", x"78", x"79", x"7b", x"74", x"76", x"79", x"76", x"74", 
        x"79", x"7f", x"83", x"83", x"7e", x"7a", x"7c", x"7f", x"85", x"8c", x"8e", x"8c", x"8c", x"9f", x"db", 
        x"b1", x"97", x"92", x"99", x"92", x"95", x"98", x"99", x"98", x"98", x"92", x"92", x"8f", x"94", x"95", 
        x"89", x"76", x"74", x"6f", x"6f", x"73", x"76", x"75", x"6f", x"8b", x"d4", x"a2", x"79", x"76", x"75", 
        x"79", x"7a", x"7b", x"78", x"75", x"75", x"79", x"7d", x"7c", x"79", x"78", x"7b", x"7e", x"7e", x"7c", 
        x"7a", x"7c", x"7b", x"8c", x"cb", x"c5", x"9a", x"8f", x"87", x"87", x"90", x"92", x"8b", x"86", x"8b", 
        x"97", x"99", x"8d", x"86", x"8d", x"92", x"91", x"8a", x"80", x"7f", x"86", x"ab", x"e6", x"f6", x"f4", 
        x"f3", x"f3", x"f3", x"f4", x"f4", x"f4", x"f4", x"f2", x"f0", x"f2", x"f3", x"f3", x"f1", x"ef", x"f1", 
        x"ef", x"ed", x"e0", x"cd", x"bd", x"be", x"ba", x"b7", x"b7", x"b8", x"b9", x"bc", x"be", x"bb", x"99", 
        x"6d", x"65", x"68", x"66", x"61", x"5d", x"52", x"29", x"0b", x"06", x"19", x"1f", x"1a", x"16", x"15", 
        x"2e", x"47", x"47", x"45", x"42", x"42", x"40", x"3d", x"3e", x"37", x"3c", x"59", x"64", x"6f", x"6c", 
        x"6b", x"6b", x"6a", x"68", x"6f", x"73", x"6e", x"6e", x"6c", x"66", x"68", x"61", x"2a", x"0c", x"1e", 
        x"41", x"40", x"34", x"33", x"36", x"38", x"36", x"34", x"27", x"16", x"19", x"18", x"0e", x"0a", x"0d", 
        x"09", x"06", x"0f", x"20", x"20", x"21", x"21", x"21", x"23", x"21", x"1f", x"19", x"18", x"13", x"07", 
        x"07", x"0a", x"14", x"17", x"11", x"0f", x"10", x"11", x"11", x"10", x"09", x"07", x"07", x"0b", x"0b", 
        x"11", x"32", x"20", x"19", x"13", x"12", x"11", x"10", x"0d", x"09", x"06", x"05", x"03", x"03", x"05", 
        x"06", x"1a", x"15", x"10", x"0a", x"0a", x"0b", x"34", x"85", x"90", x"8d", x"93", x"94", x"8e", x"85", 
        x"7e", x"79", x"73", x"45", x"2c", x"22", x"0c", x"03", x"03", x"02", x"03", x"05", x"40", x"57", x"53", 
        x"52", x"53", x"5d", x"5d", x"58", x"58", x"58", x"25", x"1b", x"1d", x"1f", x"1d", x"13", x"0a", x"07", 
        x"39", x"57", x"46", x"37", x"30", x"43", x"6a", x"55", x"2f", x"36", x"76", x"42", x"23", x"44", x"5a", 
        x"35", x"1d", x"22", x"32", x"71", x"70", x"4c", x"24", x"27", x"45", x"4d", x"66", x"34", x"27", x"3a", 
        x"6d", x"57", x"21", x"2d", x"2e", x"55", x"72", x"66", x"77", x"5f", x"4a", x"44", x"31", x"32", x"39", 
        x"71", x"65", x"7e", x"95", x"61", x"63", x"47", x"27", x"31", x"5b", x"79", x"8e", x"8c", x"47", x"3d", 
        x"81", x"5f", x"58", x"91", x"7a", x"56", x"60", x"6c", x"5e", x"5e", x"5b", x"5e", x"51", x"5b", x"73", 
        x"75", x"76", x"62", x"7a", x"74", x"4c", x"42", x"60", x"85", x"91", x"72", x"5c", x"76", x"8b", x"a3", 
        x"90", x"b0", x"dc", x"de", x"ab", x"b1", x"b5", x"b9", x"8d", x"74", x"89", x"7d", x"9f", x"a5", x"7d", 
        x"5c", x"83", x"90", x"6d", x"4f", x"85", x"8f", x"86", x"91", x"a4", x"af", x"b0", x"9d", x"9b", x"98", 
        x"b4", x"ae", x"b6", x"af", x"a3", x"a7", x"b2", x"b5", x"45", x"38", x"6d", x"6b", x"6c", x"bd", x"d8", 
        x"c9", x"c6", x"c0", x"bc", x"b9", x"b9", x"c5", x"c2", x"b3", x"77", x"58", x"62", x"4e", x"97", x"88", 
        x"7d", x"7c", x"75", x"a3", x"d9", x"d3", x"d5", x"d5", x"d2", x"d9", x"dd", x"cd", x"d0", x"d0", x"d0", 
        x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"d1", x"d3", x"d3", x"d2", x"d1", x"d2", x"d3", 
        x"d2", x"d0", x"d2", x"d3", x"d2", x"d3", x"d4", x"d3", x"d3", x"d3", x"d2", x"d1", x"d1", x"d2", x"d2", 
        x"d2", x"d2", x"d2", x"d2", x"d3", x"d4", x"d5", x"d4", x"d3", x"d5", x"d3", x"e0", x"df", x"a2", x"86", 
        x"71", x"6d", x"67", x"6a", x"78", x"a5", x"a9", x"82", x"77", x"79", x"7b", x"7b", x"76", x"72", x"70", 
        x"6d", x"70", x"79", x"7b", x"7b", x"81", x"89", x"82", x"80", x"80", x"84", x"85", x"8b", x"8e", x"81", 
        x"70", x"67", x"70", x"7a", x"7d", x"7e", x"83", x"84", x"7e", x"77", x"74", x"75", x"77", x"7d", x"82", 
        x"87", x"88", x"82", x"7c", x"97", x"dd", x"c7", x"9a", x"93", x"8b", x"83", x"85", x"8a", x"8d", x"8c", 
        x"89", x"83", x"7c", x"7e", x"84", x"8b", x"8d", x"89", x"83", x"80", x"7d", x"7e", x"84", x"89", x"8c", 
        x"8f", x"8d", x"86", x"83", x"87", x"8c", x"90", x"91", x"92", x"91", x"8c", x"83", x"82", x"94", x"97", 
        x"b5", x"e5", x"b8", x"9b", x"98", x"95", x"96", x"96", x"95", x"94", x"91", x"8e", x"8a", x"8b", x"8f", 
        x"90", x"8c", x"8c", x"85", x"81", x"7f", x"7c", x"7f", x"84", x"85", x"87", x"89", x"85", x"86", x"8d", 
        x"93", x"95", x"96", x"94", x"90", x"8f", x"90", x"91", x"a6", x"dc", x"af", x"7c", x"7a", x"7d", x"7c", 
        x"7a", x"78", x"7c", x"82", x"86", x"84", x"81", x"79", x"72", x"6f", x"71", x"74", x"77", x"78", x"75", 
        x"6e", x"68", x"68", x"68", x"6e", x"7c", x"7a", x"71", x"66", x"61", x"64", x"63", x"62", x"83", x"ca", 
        x"d7", x"be", x"b7", x"b8", x"bd", x"bd", x"c0", x"c3", x"c1", x"bb", x"c0", x"c7", x"c4", x"bf", x"bd", 
        x"b7", x"b5", x"bc", x"c2", x"c1", x"bd", x"be", x"c0", x"bd", x"bf", x"c3", x"bd", x"b8", x"b8", x"bb", 
        x"b9", x"c0", x"d7", x"96", x"7a", x"7e", x"83", x"8d", x"8e", x"86", x"84", x"86", x"86", x"8b", x"91", 
        x"90", x"8b", x"8a", x"8c", x"88", x"88", x"85", x"82", x"83", x"86", x"84", x"7e", x"7a", x"7c", x"7d", 
        x"83", x"bc", x"cb", x"82", x"76", x"78", x"7a", x"7e", x"7f", x"7d", x"7c", x"80", x"81", x"7c", x"79", 
        x"7e", x"85", x"87", x"84", x"80", x"80", x"85", x"87", x"8d", x"90", x"8d", x"8c", x"8b", x"9c", x"dd", 
        x"b4", x"95", x"90", x"96", x"8e", x"8f", x"93", x"93", x"92", x"94", x"90", x"92", x"92", x"95", x"98", 
        x"90", x"81", x"7e", x"75", x"73", x"74", x"76", x"77", x"72", x"8c", x"d4", x"a5", x"7c", x"7a", x"7d", 
        x"7d", x"79", x"7a", x"78", x"74", x"70", x"74", x"7b", x"7f", x"79", x"77", x"7a", x"7f", x"7e", x"7a", 
        x"75", x"77", x"77", x"86", x"c6", x"c3", x"9b", x"96", x"8d", x"84", x"87", x"90", x"94", x"8c", x"8a", 
        x"8f", x"95", x"96", x"92", x"8b", x"88", x"8b", x"94", x"91", x"88", x"81", x"a4", x"e3", x"f7", x"f3", 
        x"f2", x"f2", x"f2", x"f4", x"f5", x"f5", x"f1", x"f2", x"f2", x"f0", x"f1", x"f2", x"f2", x"f0", x"f1", 
        x"ef", x"ee", x"e3", x"d0", x"be", x"b7", x"ba", x"bb", x"bb", x"be", x"bc", x"b9", x"b5", x"b6", x"b0", 
        x"84", x"63", x"64", x"62", x"5f", x"5e", x"59", x"30", x"0b", x"05", x"19", x"1f", x"1e", x"1a", x"25", 
        x"40", x"4a", x"46", x"42", x"40", x"3f", x"41", x"44", x"48", x"3e", x"3d", x"5a", x"66", x"71", x"6e", 
        x"6c", x"6d", x"6e", x"69", x"6a", x"70", x"72", x"6e", x"6b", x"66", x"65", x"62", x"2d", x"0b", x"1c", 
        x"3e", x"3f", x"39", x"39", x"37", x"34", x"31", x"30", x"27", x"17", x"1c", x"1a", x"0f", x"08", x"0c", 
        x"09", x"08", x"0d", x"1e", x"1f", x"21", x"23", x"21", x"20", x"1c", x"1d", x"18", x"19", x"15", x"0a", 
        x"08", x"09", x"11", x"17", x"13", x"13", x"15", x"16", x"11", x"08", x"04", x"08", x"0b", x"0b", x"0a", 
        x"11", x"2f", x"1d", x"16", x"13", x"13", x"12", x"12", x"10", x"08", x"04", x"03", x"03", x"04", x"06", 
        x"04", x"19", x"15", x"10", x"0b", x"0d", x"0f", x"33", x"85", x"91", x"8c", x"91", x"92", x"91", x"8c", 
        x"86", x"79", x"71", x"42", x"25", x"1d", x"0b", x"04", x"04", x"01", x"03", x"04", x"3c", x"54", x"53", 
        x"50", x"50", x"5b", x"5c", x"58", x"5a", x"59", x"25", x"17", x"19", x"1e", x"1a", x"10", x"0c", x"0a", 
        x"32", x"4a", x"45", x"2f", x"36", x"5c", x"6d", x"66", x"48", x"4a", x"65", x"2c", x"1f", x"47", x"51", 
        x"26", x"10", x"1a", x"30", x"63", x"60", x"39", x"21", x"21", x"32", x"3f", x"4e", x"5c", x"45", x"55", 
        x"72", x"34", x"1c", x"39", x"44", x"36", x"53", x"56", x"48", x"55", x"50", x"42", x"46", x"4a", x"34", 
        x"6d", x"5c", x"6a", x"7d", x"46", x"43", x"32", x"2f", x"39", x"6d", x"7e", x"89", x"79", x"37", x"36", 
        x"62", x"48", x"4f", x"6d", x"81", x"5e", x"47", x"55", x"6a", x"6a", x"5f", x"6f", x"6a", x"61", x"55", 
        x"58", x"70", x"5a", x"57", x"5a", x"60", x"57", x"7c", x"7a", x"79", x"8d", x"72", x"69", x"8b", x"a1", 
        x"9f", x"b2", x"c3", x"b2", x"98", x"aa", x"91", x"be", x"93", x"6a", x"8f", x"71", x"70", x"92", x"6e", 
        x"4c", x"7c", x"76", x"7a", x"52", x"7d", x"87", x"89", x"97", x"a4", x"b0", x"9e", x"9e", x"9f", x"8f", 
        x"b7", x"c1", x"b7", x"a2", x"c0", x"b5", x"c5", x"c3", x"48", x"3b", x"6f", x"6e", x"6b", x"b3", x"ba", 
        x"b0", x"a4", x"a3", x"b6", x"b5", x"b0", x"cf", x"d9", x"cf", x"84", x"52", x"5e", x"51", x"a2", x"8e", 
        x"7d", x"7e", x"74", x"9f", x"da", x"d4", x"d7", x"d6", x"d2", x"d8", x"de", x"cd", x"d0", x"d1", x"d0", 
        x"d1", x"d1", x"d2", x"d0", x"cf", x"d0", x"d1", x"d1", x"d1", x"d2", x"d3", x"d2", x"d2", x"d2", x"d2", 
        x"d2", x"d1", x"d1", x"d1", x"d1", x"d3", x"d5", x"d2", x"d4", x"d4", x"d3", x"d2", x"d1", x"d3", x"d3", 
        x"d3", x"d3", x"d4", x"d4", x"d6", x"d7", x"d5", x"d5", x"d6", x"d7", x"d2", x"de", x"de", x"ac", x"8f", 
        x"7a", x"7a", x"6f", x"6f", x"78", x"9d", x"9d", x"7d", x"78", x"80", x"7d", x"74", x"6d", x"6d", x"78", 
        x"7e", x"80", x"81", x"7e", x"7b", x"7c", x"83", x"8a", x"93", x"96", x"96", x"93", x"8c", x"8d", x"80", 
        x"76", x"75", x"82", x"8c", x"83", x"7d", x"77", x"72", x"71", x"6c", x"69", x"6f", x"74", x"78", x"76", 
        x"73", x"70", x"6c", x"6b", x"8d", x"db", x"bf", x"85", x"7e", x"7e", x"82", x"8c", x"94", x"98", x"95", 
        x"8f", x"87", x"83", x"88", x"91", x"97", x"98", x"97", x"93", x"8c", x"8a", x"8d", x"93", x"97", x"97", 
        x"93", x"8c", x"83", x"80", x"85", x"8a", x"8e", x"8e", x"8d", x"8b", x"82", x"7a", x"7c", x"86", x"89", 
        x"ac", x"e2", x"ab", x"8d", x"8f", x"90", x"91", x"90", x"92", x"92", x"95", x"9b", x"9d", x"9c", x"99", 
        x"96", x"93", x"95", x"96", x"98", x"9a", x"9b", x"9e", x"a0", x"9f", x"9f", x"a0", x"9d", x"98", x"98", 
        x"99", x"98", x"96", x"91", x"8d", x"8b", x"8a", x"8a", x"9d", x"d7", x"ad", x"73", x"70", x"75", x"78", 
        x"77", x"73", x"6d", x"6a", x"6d", x"72", x"74", x"71", x"6d", x"6d", x"6d", x"70", x"74", x"79", x"7c", 
        x"79", x"73", x"6f", x"70", x"75", x"7f", x"7f", x"7c", x"78", x"76", x"72", x"6d", x"6d", x"89", x"cd", 
        x"d5", x"bd", x"b9", x"b8", x"b8", x"b3", x"b2", x"bd", x"c2", x"bf", x"bc", x"bc", x"b7", x"b4", x"b9", 
        x"bc", x"ba", x"bb", x"be", x"c1", x"be", x"bf", x"c1", x"bf", x"bc", x"bc", x"bb", x"bb", x"bb", x"bd", 
        x"bf", x"c1", x"d7", x"9f", x"87", x"8f", x"93", x"95", x"8d", x"86", x"84", x"85", x"8b", x"90", x"91", 
        x"8b", x"83", x"7f", x"7e", x"83", x"88", x"89", x"85", x"80", x"7c", x"7c", x"7f", x"86", x"8f", x"8c", 
        x"8b", x"be", x"d0", x"8e", x"7f", x"85", x"8c", x"8d", x"88", x"82", x"81", x"82", x"81", x"7f", x"7e", 
        x"7d", x"7e", x"7e", x"80", x"82", x"84", x"89", x"8a", x"8c", x"8c", x"88", x"8b", x"89", x"98", x"d8", 
        x"b5", x"8d", x"8a", x"90", x"8b", x"8e", x"92", x"93", x"93", x"91", x"8e", x"95", x"90", x"97", x"9b", 
        x"93", x"7f", x"7b", x"73", x"70", x"74", x"76", x"76", x"75", x"8e", x"d5", x"a9", x"76", x"75", x"73", 
        x"78", x"7c", x"7d", x"7e", x"78", x"6e", x"73", x"7c", x"80", x"7f", x"7c", x"7a", x"7a", x"7a", x"79", 
        x"7a", x"7b", x"7b", x"87", x"c5", x"c3", x"8a", x"8c", x"8f", x"89", x"84", x"87", x"8f", x"92", x"90", 
        x"8e", x"8e", x"94", x"9b", x"95", x"88", x"81", x"87", x"91", x"90", x"89", x"a0", x"e0", x"f3", x"f2", 
        x"f1", x"f1", x"f2", x"f4", x"f4", x"f3", x"f0", x"f0", x"f0", x"ef", x"f0", x"f2", x"f2", x"f1", x"f0", 
        x"f1", x"ef", x"e5", x"d0", x"bc", x"b7", x"b9", x"b8", x"b7", x"b9", x"bb", x"bf", x"be", x"b6", x"b6", 
        x"9f", x"70", x"6a", x"6a", x"63", x"60", x"5b", x"33", x"0d", x"07", x"19", x"22", x"1e", x"1c", x"36", 
        x"48", x"45", x"46", x"48", x"4a", x"46", x"41", x"40", x"43", x"3c", x"39", x"58", x"63", x"71", x"71", 
        x"6e", x"6d", x"6e", x"6d", x"6a", x"6b", x"72", x"71", x"6c", x"66", x"67", x"67", x"30", x"0b", x"16", 
        x"3b", x"3f", x"3b", x"3a", x"36", x"36", x"35", x"34", x"2d", x"1d", x"1c", x"1a", x"10", x"09", x"0c", 
        x"0a", x"07", x"08", x"16", x"1c", x"1f", x"24", x"21", x"1f", x"1e", x"1e", x"1c", x"1d", x"18", x"0a", 
        x"06", x"07", x"0e", x"16", x"12", x"11", x"15", x"16", x"10", x"06", x"06", x"0a", x"0e", x"0c", x"0a", 
        x"0f", x"2a", x"1e", x"15", x"18", x"16", x"17", x"17", x"13", x"0a", x"07", x"07", x"06", x"06", x"05", 
        x"04", x"17", x"18", x"0e", x"0b", x"0d", x"11", x"30", x"85", x"94", x"8d", x"90", x"91", x"8c", x"8c", 
        x"86", x"7d", x"78", x"48", x"26", x"1f", x"0f", x"05", x"04", x"04", x"04", x"03", x"34", x"53", x"4c", 
        x"4a", x"4e", x"59", x"5a", x"5a", x"5b", x"59", x"2b", x"1f", x"20", x"21", x"1c", x"13", x"0d", x"0b", 
        x"7e", x"70", x"3b", x"19", x"2b", x"57", x"65", x"90", x"80", x"32", x"37", x"34", x"33", x"58", x"4a", 
        x"23", x"22", x"18", x"35", x"57", x"66", x"39", x"17", x"2a", x"61", x"79", x"48", x"7e", x"78", x"58", 
        x"72", x"3c", x"15", x"3d", x"5b", x"26", x"27", x"45", x"40", x"40", x"50", x"3b", x"59", x"68", x"35", 
        x"40", x"48", x"71", x"7d", x"4b", x"3a", x"23", x"31", x"2f", x"3e", x"5a", x"55", x"5b", x"5d", x"53", 
        x"55", x"5f", x"74", x"67", x"67", x"4f", x"65", x"68", x"7a", x"74", x"66", x"6a", x"61", x"53", x"6e", 
        x"6b", x"6f", x"56", x"44", x"61", x"66", x"5f", x"7a", x"75", x"68", x"7b", x"84", x"87", x"8b", x"87", 
        x"90", x"a0", x"9d", x"90", x"ac", x"b8", x"b0", x"cd", x"ae", x"94", x"73", x"8e", x"83", x"7e", x"72", 
        x"50", x"5f", x"90", x"a7", x"58", x"74", x"8c", x"96", x"ae", x"aa", x"a2", x"98", x"99", x"98", x"9c", 
        x"be", x"b5", x"9a", x"a7", x"c5", x"c1", x"cd", x"bc", x"49", x"3b", x"6c", x"6d", x"6d", x"ad", x"b6", 
        x"b5", x"a1", x"a3", x"bc", x"bb", x"ad", x"be", x"cc", x"d0", x"81", x"4d", x"60", x"53", x"a3", x"89", 
        x"7e", x"80", x"75", x"9d", x"db", x"d4", x"d5", x"d4", x"d2", x"d6", x"de", x"ce", x"d0", x"d1", x"d0", 
        x"d1", x"d1", x"d2", x"d0", x"ce", x"ce", x"d1", x"d2", x"d1", x"d2", x"d2", x"d2", x"d1", x"d1", x"d1", 
        x"d2", x"d2", x"d1", x"d0", x"d1", x"d3", x"d5", x"d4", x"d5", x"d5", x"d3", x"d1", x"d1", x"d2", x"d4", 
        x"d3", x"d3", x"d4", x"d6", x"d6", x"d5", x"d4", x"d6", x"d6", x"d5", x"d0", x"de", x"df", x"a1", x"84", 
        x"73", x"71", x"6f", x"71", x"7e", x"ac", x"af", x"8b", x"70", x"6d", x"70", x"6e", x"6f", x"73", x"75", 
        x"6f", x"68", x"65", x"65", x"66", x"66", x"66", x"6f", x"78", x"7e", x"7f", x"81", x"80", x"7e", x"6e", 
        x"68", x"6e", x"81", x"8f", x"7f", x"78", x"71", x"6d", x"70", x"70", x"74", x"7d", x"81", x"81", x"7c", 
        x"78", x"75", x"77", x"76", x"8f", x"db", x"c4", x"8b", x"87", x"84", x"88", x"8c", x"8f", x"8f", x"8a", 
        x"82", x"7c", x"7b", x"80", x"88", x"8b", x"8a", x"87", x"81", x"76", x"78", x"7b", x"7f", x"83", x"84", 
        x"80", x"7b", x"7a", x"7f", x"88", x"92", x"9a", x"9b", x"98", x"92", x"89", x"83", x"86", x"90", x"93", 
        x"af", x"e3", x"b4", x"98", x"9b", x"9b", x"9d", x"9c", x"9c", x"9b", x"9a", x"98", x"95", x"93", x"91", 
        x"90", x"8d", x"8d", x"8e", x"90", x"92", x"93", x"93", x"92", x"90", x"8e", x"8c", x"8d", x"8d", x"8d", 
        x"8e", x"8d", x"8b", x"8a", x"8b", x"91", x"98", x"95", x"9c", x"d6", x"b2", x"74", x"6d", x"73", x"7b", 
        x"80", x"81", x"7b", x"76", x"77", x"7e", x"82", x"85", x"86", x"88", x"88", x"81", x"7d", x"7d", x"7e", 
        x"7e", x"7d", x"7a", x"7d", x"7e", x"81", x"7c", x"77", x"75", x"76", x"76", x"75", x"75", x"8b", x"c8", 
        x"cd", x"b5", x"b8", x"bf", x"c2", x"c0", x"bd", x"c1", x"c5", x"c3", x"c6", x"ca", x"c6", x"c0", x"c0", 
        x"c1", x"c3", x"c5", x"c8", x"cb", x"c1", x"bb", x"b8", x"b8", x"b7", x"b6", x"b6", x"b6", x"b4", x"b7", 
        x"bc", x"be", x"d5", x"9e", x"82", x"89", x"8b", x"88", x"7f", x"7d", x"80", x"82", x"8a", x"8f", x"8d", 
        x"86", x"82", x"81", x"83", x"8d", x"91", x"8f", x"89", x"82", x"7e", x"82", x"8b", x"94", x"97", x"8e", 
        x"88", x"ba", x"d0", x"8d", x"7d", x"84", x"86", x"82", x"7c", x"79", x"79", x"7b", x"7c", x"7a", x"79", 
        x"7b", x"7f", x"82", x"84", x"87", x"89", x"8d", x"90", x"8f", x"91", x"90", x"92", x"8e", x"99", x"d6", 
        x"b7", x"8b", x"8d", x"91", x"8b", x"8e", x"91", x"92", x"92", x"90", x"8d", x"96", x"8e", x"98", x"9c", 
        x"95", x"7c", x"79", x"72", x"6e", x"72", x"74", x"71", x"6f", x"88", x"d3", x"b1", x"7b", x"7a", x"76", 
        x"75", x"75", x"77", x"7c", x"7a", x"6d", x"6d", x"74", x"79", x"7e", x"7f", x"7c", x"79", x"78", x"77", 
        x"77", x"75", x"71", x"7a", x"bd", x"c6", x"8d", x"85", x"8a", x"8b", x"86", x"83", x"87", x"90", x"94", 
        x"94", x"8d", x"8a", x"8f", x"93", x"91", x"8b", x"83", x"7f", x"81", x"86", x"a2", x"e2", x"f5", x"f1", 
        x"f1", x"f1", x"f3", x"f4", x"f4", x"f2", x"f1", x"f0", x"ef", x"f0", x"f2", x"f3", x"f1", x"f3", x"f0", 
        x"f4", x"f1", x"e6", x"d1", x"bc", x"b3", x"b5", x"b9", x"bd", x"bc", x"b8", x"b8", x"b8", x"b5", x"ba", 
        x"b9", x"86", x"69", x"65", x"5f", x"61", x"5c", x"39", x"11", x"08", x"16", x"20", x"1c", x"23", x"44", 
        x"4b", x"43", x"44", x"49", x"47", x"43", x"3f", x"3f", x"42", x"41", x"3e", x"5a", x"62", x"71", x"72", 
        x"6f", x"6c", x"6c", x"6f", x"6c", x"6a", x"6f", x"72", x"6d", x"67", x"65", x"64", x"32", x"0e", x"15", 
        x"3c", x"42", x"3d", x"3a", x"38", x"3b", x"3b", x"37", x"2d", x"19", x"15", x"16", x"11", x"0b", x"0e", 
        x"0b", x"08", x"0e", x"1b", x"22", x"24", x"29", x"24", x"21", x"20", x"1e", x"1d", x"1c", x"16", x"09", 
        x"05", x"08", x"10", x"15", x"12", x"14", x"15", x"0f", x"09", x"07", x"09", x"0c", x"10", x"0e", x"0d", 
        x"0f", x"27", x"1f", x"12", x"17", x"15", x"15", x"11", x"0e", x"05", x"04", x"06", x"05", x"08", x"07", 
        x"05", x"13", x"16", x"0c", x"0c", x"0d", x"11", x"2b", x"81", x"94", x"8c", x"8f", x"90", x"88", x"89", 
        x"81", x"79", x"77", x"4f", x"2c", x"24", x"11", x"04", x"03", x"04", x"04", x"03", x"2f", x"53", x"4c", 
        x"4b", x"4e", x"59", x"59", x"59", x"57", x"59", x"2f", x"23", x"23", x"22", x"20", x"1a", x"17", x"1d", 
        x"77", x"57", x"2e", x"28", x"2e", x"28", x"33", x"76", x"78", x"3d", x"47", x"3b", x"2c", x"44", x"4b", 
        x"3c", x"2a", x"1e", x"2a", x"46", x"5f", x"3b", x"1a", x"4d", x"66", x"4d", x"4c", x"60", x"6d", x"5e", 
        x"52", x"38", x"1a", x"26", x"3f", x"49", x"32", x"3a", x"54", x"3c", x"3f", x"4c", x"50", x"44", x"3b", 
        x"4c", x"40", x"5e", x"7c", x"50", x"26", x"1b", x"28", x"2c", x"41", x"45", x"32", x"69", x"74", x"75", 
        x"83", x"89", x"75", x"6b", x"69", x"7d", x"91", x"6b", x"70", x"54", x"39", x"5f", x"73", x"70", x"64", 
        x"62", x"7a", x"88", x"74", x"68", x"56", x"63", x"4e", x"5a", x"6e", x"7b", x"8a", x"79", x"71", x"60", 
        x"4e", x"65", x"7a", x"79", x"96", x"b0", x"a4", x"9f", x"ab", x"b5", x"73", x"88", x"a8", x"79", x"4f", 
        x"40", x"65", x"a4", x"98", x"4c", x"6f", x"95", x"99", x"a5", x"99", x"95", x"9e", x"99", x"95", x"ae", 
        x"af", x"84", x"ab", x"b3", x"b8", x"b6", x"b7", x"b6", x"4d", x"3a", x"6c", x"71", x"6b", x"b3", x"bf", 
        x"b6", x"c3", x"c3", x"b1", x"a9", x"9f", x"a7", x"c6", x"ce", x"81", x"49", x"5c", x"55", x"9d", x"7e", 
        x"7f", x"7c", x"74", x"9c", x"dc", x"d4", x"d3", x"d4", x"d2", x"d5", x"dd", x"ce", x"d0", x"cf", x"d0", 
        x"d2", x"d2", x"d3", x"d1", x"ce", x"ce", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d1", x"d0", x"d1", 
        x"d2", x"d1", x"d0", x"d0", x"d2", x"d3", x"d4", x"d6", x"d6", x"d5", x"d2", x"d1", x"d1", x"d2", x"d5", 
        x"d2", x"d1", x"d4", x"d7", x"d5", x"d2", x"d5", x"d8", x"d6", x"d6", x"d2", x"de", x"e0", x"b1", x"96", 
        x"8c", x"8c", x"83", x"7e", x"77", x"98", x"9f", x"7c", x"69", x"7b", x"8a", x"8c", x"85", x"83", x"84", 
        x"80", x"7a", x"7a", x"7e", x"82", x"86", x"86", x"86", x"85", x"86", x"8b", x"93", x"96", x"98", x"8f", 
        x"8a", x"85", x"88", x"86", x"79", x"76", x"75", x"76", x"79", x"78", x"76", x"70", x"6b", x"67", x"61", 
        x"5d", x"5d", x"60", x"66", x"8d", x"da", x"b9", x"71", x"69", x"74", x"7d", x"84", x"87", x"88", x"86", 
        x"83", x"80", x"80", x"8d", x"92", x"94", x"92", x"8f", x"8a", x"86", x"8e", x"98", x"a4", x"aa", x"a8", 
        x"a0", x"99", x"8d", x"87", x"8a", x"8d", x"90", x"90", x"8e", x"8b", x"81", x"75", x"75", x"7e", x"85", 
        x"a9", x"e0", x"a7", x"84", x"81", x"7f", x"82", x"86", x"86", x"83", x"84", x"85", x"86", x"89", x"8f", 
        x"95", x"99", x"98", x"97", x"96", x"95", x"93", x"90", x"94", x"98", x"9b", x"9d", x"a0", x"a2", x"a4", 
        x"9f", x"9c", x"a0", x"a1", x"a1", x"a0", x"9f", x"9b", x"a3", x"d8", x"b9", x"7d", x"75", x"73", x"75", 
        x"77", x"7d", x"7b", x"75", x"6f", x"6b", x"69", x"6a", x"6b", x"70", x"74", x"72", x"6d", x"69", x"63", 
        x"62", x"66", x"6b", x"71", x"72", x"78", x"79", x"78", x"77", x"74", x"72", x"71", x"70", x"7f", x"bc", 
        x"d7", x"c8", x"c7", x"c7", x"c9", x"c9", x"c9", x"c9", x"c7", x"bf", x"bc", x"be", x"bc", x"bb", x"be", 
        x"c2", x"c2", x"bf", x"bf", x"c3", x"bc", x"b7", x"b6", x"b6", x"b4", x"b2", x"b4", x"bc", x"be", x"bf", 
        x"be", x"be", x"d7", x"a9", x"8f", x"8e", x"88", x"86", x"89", x"92", x"99", x"96", x"8d", x"8c", x"8b", 
        x"8e", x"91", x"8f", x"8a", x"89", x"88", x"86", x"82", x"81", x"85", x"88", x"85", x"84", x"82", x"7b", 
        x"7a", x"b2", x"d3", x"8a", x"7a", x"81", x"81", x"7d", x"7d", x"80", x"81", x"85", x"86", x"7f", x"7b", 
        x"81", x"87", x"8a", x"8b", x"8d", x"8c", x"8e", x"91", x"8c", x"8f", x"8d", x"8e", x"8d", x"97", x"d3", 
        x"ba", x"8a", x"8a", x"8c", x"88", x"8b", x"8e", x"91", x"91", x"91", x"8d", x"94", x"8d", x"96", x"9a", 
        x"94", x"7b", x"79", x"73", x"70", x"76", x"7a", x"7a", x"78", x"8d", x"d3", x"b3", x"79", x"79", x"78", 
        x"77", x"77", x"74", x"76", x"79", x"75", x"78", x"79", x"78", x"7a", x"7a", x"79", x"79", x"78", x"77", 
        x"7c", x"7c", x"79", x"80", x"bd", x"c6", x"91", x"84", x"87", x"8f", x"92", x"8d", x"86", x"85", x"90", 
        x"9d", x"9c", x"91", x"87", x"83", x"88", x"8f", x"8f", x"87", x"7f", x"7c", x"94", x"db", x"f5", x"f1", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f1", x"f1", x"f2", x"f3", x"f3", x"f1", x"ef", x"ed", 
        x"f1", x"ef", x"e5", x"d1", x"bd", x"be", x"bd", x"b7", x"b5", x"b3", x"b5", x"bb", x"bb", x"b3", x"b2", 
        x"b9", x"9e", x"76", x"68", x"6c", x"6a", x"64", x"3f", x"11", x"06", x"18", x"25", x"20", x"32", x"4c", 
        x"4a", x"44", x"44", x"49", x"47", x"44", x"43", x"44", x"46", x"43", x"3d", x"58", x"61", x"70", x"70", 
        x"6f", x"6e", x"70", x"6e", x"6b", x"69", x"6a", x"6d", x"6d", x"68", x"66", x"69", x"39", x"11", x"13", 
        x"35", x"3a", x"37", x"3d", x"3a", x"3a", x"3b", x"3b", x"2c", x"11", x"12", x"16", x"13", x"0c", x"0e", 
        x"0b", x"08", x"08", x"11", x"1a", x"1c", x"21", x"1c", x"19", x"1b", x"1b", x"1b", x"1c", x"17", x"09", 
        x"04", x"08", x"11", x"15", x"14", x"15", x"11", x"08", x"04", x"08", x"09", x"0c", x"0f", x"0f", x"0f", 
        x"10", x"24", x"1f", x"11", x"16", x"13", x"11", x"0d", x"0e", x"07", x"05", x"05", x"06", x"0a", x"0b", 
        x"06", x"13", x"1c", x"10", x"0e", x"0e", x"14", x"28", x"7c", x"94", x"8c", x"8e", x"91", x"8a", x"8c", 
        x"86", x"7c", x"78", x"50", x"29", x"1d", x"0a", x"03", x"03", x"03", x"04", x"03", x"2d", x"53", x"50", 
        x"4e", x"4f", x"5a", x"5c", x"59", x"55", x"58", x"2f", x"1e", x"1e", x"20", x"21", x"1c", x"25", x"37", 
        x"2e", x"38", x"33", x"4a", x"37", x"33", x"67", x"52", x"77", x"90", x"63", x"3a", x"43", x"52", x"59", 
        x"54", x"38", x"29", x"28", x"28", x"4a", x"4e", x"26", x"5b", x"48", x"3a", x"65", x"88", x"54", x"39", 
        x"3f", x"25", x"2a", x"3a", x"3a", x"34", x"2e", x"46", x"5e", x"50", x"38", x"4d", x"56", x"5e", x"3f", 
        x"3e", x"46", x"6c", x"83", x"54", x"36", x"46", x"5a", x"56", x"31", x"23", x"2d", x"62", x"4b", x"5f", 
        x"82", x"74", x"6c", x"77", x"77", x"77", x"74", x"6b", x"6d", x"49", x"5e", x"77", x"5d", x"45", x"4c", 
        x"56", x"59", x"71", x"83", x"83", x"75", x"88", x"6f", x"49", x"4c", x"6b", x"7e", x"76", x"8a", x"7e", 
        x"4f", x"5f", x"87", x"72", x"75", x"8c", x"94", x"9a", x"92", x"8e", x"6e", x"51", x"5d", x"65", x"54", 
        x"3f", x"6c", x"79", x"6a", x"4b", x"78", x"93", x"8a", x"87", x"89", x"8b", x"8e", x"96", x"9c", x"84", 
        x"7f", x"a9", x"c1", x"c2", x"d5", x"c4", x"c8", x"ad", x"42", x"37", x"6c", x"6f", x"6d", x"bb", x"d5", 
        x"c8", x"c4", x"c7", x"c0", x"b1", x"ad", x"b8", x"ae", x"aa", x"75", x"4c", x"55", x"52", x"a0", x"86", 
        x"7f", x"7e", x"74", x"9a", x"dc", x"d5", x"d2", x"d6", x"d3", x"d4", x"dc", x"cf", x"d0", x"ce", x"d0", 
        x"d2", x"d2", x"d3", x"d1", x"cf", x"cf", x"d1", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d1", x"d2", 
        x"d2", x"d1", x"d0", x"d1", x"d3", x"d3", x"d4", x"d5", x"d5", x"d4", x"d2", x"d1", x"d1", x"d1", x"d3", 
        x"d1", x"d1", x"d4", x"d6", x"d4", x"d2", x"d2", x"d4", x"d2", x"d3", x"d1", x"dd", x"e0", x"a3", x"7e", 
        x"68", x"67", x"62", x"6d", x"7e", x"ab", x"b5", x"86", x"79", x"9c", x"af", x"a0", x"7b", x"62", x"64", 
        x"65", x"66", x"67", x"68", x"65", x"5f", x"5c", x"59", x"5a", x"62", x"71", x"7e", x"7e", x"7d", x"73", 
        x"6c", x"6d", x"77", x"7f", x"76", x"74", x"77", x"7b", x"7e", x"7d", x"7d", x"7d", x"7c", x"78", x"75", 
        x"75", x"78", x"7d", x"7e", x"93", x"da", x"c7", x"8e", x"92", x"93", x"99", x"99", x"9b", x"98", x"8e", 
        x"84", x"7f", x"80", x"8a", x"8e", x"91", x"8f", x"84", x"78", x"71", x"73", x"77", x"7c", x"81", x"82", 
        x"7e", x"79", x"6f", x"6d", x"76", x"80", x"89", x"8d", x"8d", x"8b", x"85", x"7e", x"7a", x"80", x"88", 
        x"a7", x"df", x"b2", x"90", x"95", x"92", x"90", x"96", x"9f", x"a1", x"a3", x"a3", x"a0", x"9a", x"94", 
        x"91", x"90", x"8f", x"8e", x"8d", x"8c", x"8c", x"8b", x"85", x"84", x"88", x"8a", x"8c", x"8b", x"8a", 
        x"87", x"88", x"8a", x"8b", x"8b", x"8a", x"89", x"84", x"92", x"d0", x"b2", x"6f", x"69", x"6b", x"6d", 
        x"6f", x"77", x"7d", x"80", x"7f", x"7d", x"7a", x"7a", x"76", x"76", x"7d", x"83", x"84", x"84", x"7d", 
        x"7a", x"7a", x"7a", x"7d", x"80", x"8c", x"8c", x"8a", x"89", x"80", x"75", x"6f", x"6c", x"80", x"c1", 
        x"d6", x"c0", x"c1", x"c2", x"c1", x"b9", x"b1", x"b5", x"b7", x"b2", x"b3", x"b7", x"b6", x"b1", x"b4", 
        x"bd", x"c7", x"c6", x"c3", x"c4", x"c6", x"c0", x"be", x"c3", x"c7", x"c7", x"c7", x"c9", x"c8", x"c8", 
        x"c7", x"c4", x"d9", x"a7", x"84", x"83", x"82", x"88", x"8d", x"8e", x"8b", x"86", x"86", x"84", x"85", 
        x"8a", x"8e", x"8d", x"87", x"7f", x"7b", x"7f", x"85", x"8e", x"95", x"91", x"8c", x"86", x"82", x"7e", 
        x"7d", x"af", x"d2", x"91", x"7e", x"81", x"7e", x"7b", x"7b", x"7a", x"7d", x"83", x"82", x"7c", x"7a", 
        x"84", x"8c", x"8e", x"8e", x"8e", x"8b", x"89", x"8d", x"86", x"88", x"88", x"8a", x"8b", x"94", x"cc", 
        x"ba", x"84", x"89", x"8d", x"8d", x"91", x"94", x"97", x"95", x"96", x"91", x"96", x"8f", x"97", x"9b", 
        x"96", x"7d", x"7a", x"73", x"6d", x"6f", x"72", x"73", x"72", x"85", x"cb", x"b6", x"79", x"78", x"77", 
        x"7b", x"7f", x"77", x"72", x"72", x"73", x"79", x"7b", x"7e", x"80", x"80", x"7f", x"7e", x"7a", x"74", 
        x"75", x"7a", x"7d", x"84", x"bb", x"ca", x"9a", x"8d", x"8a", x"8c", x"97", x"9f", x"9d", x"95", x"8f", 
        x"96", x"9e", x"9c", x"98", x"8e", x"84", x"7f", x"82", x"8d", x"8f", x"85", x"94", x"d7", x"f6", x"f2", 
        x"f1", x"f1", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f1", x"f1", x"ee", 
        x"f0", x"ed", x"e2", x"cd", x"b9", x"ad", x"ae", x"b4", x"bb", x"bc", x"b7", x"b4", x"b7", x"b4", x"b1", 
        x"b7", x"bb", x"97", x"6d", x"6b", x"68", x"65", x"47", x"16", x"0a", x"16", x"22", x"24", x"39", x"47", 
        x"42", x"42", x"42", x"43", x"44", x"42", x"40", x"3f", x"41", x"40", x"38", x"56", x"62", x"72", x"72", 
        x"70", x"6f", x"6f", x"6f", x"6d", x"6b", x"6b", x"6d", x"6f", x"6c", x"69", x"6a", x"3c", x"11", x"0f", 
        x"33", x"3e", x"3b", x"3e", x"3b", x"38", x"36", x"39", x"2f", x"15", x"18", x"17", x"13", x"09", x"0c", 
        x"0a", x"08", x"07", x"10", x"1a", x"1d", x"21", x"1e", x"1b", x"1a", x"19", x"1a", x"1c", x"18", x"0b", 
        x"04", x"07", x"0e", x"13", x"11", x"0f", x"0a", x"05", x"06", x"0a", x"0b", x"0c", x"0f", x"0f", x"0f", 
        x"10", x"22", x"24", x"15", x"15", x"0d", x"0a", x"0a", x"10", x"0c", x"06", x"04", x"05", x"08", x"09", 
        x"05", x"0f", x"1a", x"0f", x"0f", x"0d", x"12", x"25", x"79", x"97", x"8f", x"91", x"96", x"90", x"8f", 
        x"89", x"84", x"80", x"59", x"2e", x"24", x"12", x"05", x"04", x"03", x"04", x"04", x"28", x"53", x"4f", 
        x"4c", x"4c", x"5a", x"5f", x"59", x"55", x"5a", x"34", x"1d", x"1d", x"1f", x"21", x"1c", x"18", x"22", 
        x"3b", x"68", x"4e", x"3a", x"49", x"63", x"7e", x"5d", x"5b", x"59", x"39", x"44", x"5e", x"39", x"2e", 
        x"37", x"36", x"2c", x"2d", x"43", x"44", x"33", x"28", x"3f", x"46", x"75", x"76", x"5c", x"33", x"4f", 
        x"84", x"3d", x"21", x"38", x"38", x"58", x"56", x"41", x"4b", x"54", x"54", x"3d", x"37", x"59", x"58", 
        x"3e", x"3f", x"62", x"77", x"5d", x"4d", x"5a", x"42", x"2f", x"1c", x"31", x"47", x"5c", x"66", x"6f", 
        x"79", x"4d", x"66", x"82", x"65", x"4f", x"6f", x"81", x"86", x"66", x"60", x"72", x"53", x"5e", x"46", 
        x"35", x"3f", x"55", x"68", x"68", x"89", x"63", x"5c", x"63", x"57", x"58", x"65", x"8f", x"96", x"82", 
        x"78", x"86", x"84", x"75", x"88", x"94", x"97", x"9a", x"a2", x"c4", x"a5", x"79", x"62", x"99", x"9c", 
        x"52", x"4d", x"6c", x"69", x"4d", x"77", x"92", x"89", x"8b", x"8e", x"91", x"93", x"9b", x"9c", x"87", 
        x"a3", x"be", x"c3", x"c0", x"d0", x"b4", x"a4", x"9f", x"47", x"38", x"69", x"67", x"6a", x"bb", x"d5", 
        x"bb", x"b2", x"c6", x"d6", x"cc", x"b6", x"c2", x"b1", x"a4", x"72", x"57", x"60", x"4f", x"9a", x"89", 
        x"80", x"7d", x"72", x"97", x"dc", x"d7", x"d4", x"da", x"d3", x"d4", x"dc", x"cf", x"d0", x"ce", x"d0", 
        x"d1", x"d2", x"d3", x"d2", x"d0", x"cf", x"d1", x"d2", x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d2", 
        x"d2", x"d1", x"d0", x"d2", x"d3", x"d3", x"d3", x"d4", x"d3", x"d3", x"d3", x"d2", x"d2", x"d1", x"d0", 
        x"d1", x"d2", x"d4", x"d4", x"d4", x"d4", x"d2", x"d3", x"d1", x"d3", x"d1", x"dc", x"e2", x"b2", x"95", 
        x"84", x"87", x"7a", x"71", x"70", x"91", x"9b", x"74", x"6c", x"9b", x"be", x"b8", x"8b", x"67", x"68", 
        x"6e", x"75", x"7c", x"7e", x"7d", x"7b", x"76", x"72", x"71", x"77", x"80", x"87", x"91", x"91", x"86", 
        x"7b", x"76", x"7d", x"86", x"87", x"87", x"8b", x"8e", x"8a", x"7f", x"71", x"6b", x"69", x"68", x"68", 
        x"6b", x"6f", x"71", x"70", x"8e", x"dc", x"c4", x"7c", x"75", x"7d", x"82", x"83", x"81", x"7b", x"74", 
        x"76", x"82", x"8f", x"95", x"95", x"96", x"95", x"8e", x"88", x"89", x"8f", x"92", x"95", x"97", x"99", 
        x"97", x"94", x"90", x"90", x"97", x"9e", x"a3", x"a4", x"a1", x"9a", x"91", x"87", x"7f", x"83", x"8c", 
        x"ab", x"e1", x"b2", x"8e", x"94", x"8d", x"84", x"85", x"88", x"85", x"85", x"85", x"86", x"84", x"7e", 
        x"7a", x"7a", x"80", x"86", x"89", x"88", x"87", x"87", x"88", x"8b", x"8f", x"94", x"98", x"99", x"98", 
        x"96", x"94", x"94", x"94", x"96", x"96", x"96", x"98", x"a4", x"d4", x"ba", x"81", x"84", x"7c", x"77", 
        x"77", x"78", x"7b", x"7f", x"81", x"81", x"7e", x"77", x"70", x"6d", x"6e", x"6e", x"70", x"73", x"79", 
        x"78", x"74", x"6c", x"66", x"66", x"71", x"71", x"6d", x"6d", x"6e", x"6f", x"6e", x"67", x"7c", x"bf", 
        x"d3", x"bb", x"be", x"c3", x"c2", x"bf", x"bb", x"ba", x"b9", x"b4", x"b9", x"c5", x"c9", x"c9", x"c3", 
        x"c4", x"c9", x"c8", x"c7", x"cb", x"ca", x"c3", x"bd", x"be", x"c0", x"c1", x"c0", x"c0", x"bf", x"bc", 
        x"b6", x"b5", x"cf", x"a3", x"7d", x"7d", x"7b", x"7f", x"80", x"81", x"81", x"83", x"88", x"88", x"8c", 
        x"93", x"94", x"8f", x"8a", x"8a", x"8b", x"90", x"96", x"9c", x"9d", x"93", x"8a", x"82", x"81", x"81", 
        x"82", x"af", x"d3", x"8e", x"79", x"7d", x"7c", x"7b", x"7c", x"7c", x"7d", x"7b", x"7b", x"78", x"78", 
        x"85", x"8e", x"8e", x"8e", x"8d", x"8a", x"88", x"8c", x"87", x"8b", x"8b", x"8d", x"8e", x"94", x"ca", 
        x"c1", x"85", x"8a", x"8d", x"8d", x"90", x"92", x"93", x"8f", x"92", x"8d", x"92", x"8c", x"94", x"9b", 
        x"98", x"7b", x"76", x"70", x"69", x"6a", x"6d", x"6f", x"70", x"82", x"c5", x"b8", x"78", x"75", x"77", 
        x"7a", x"7f", x"7d", x"7b", x"79", x"78", x"7b", x"7b", x"7f", x"7f", x"7f", x"7e", x"80", x"7e", x"79", 
        x"7a", x"7b", x"7e", x"86", x"bc", x"d1", x"9f", x"92", x"8d", x"86", x"87", x"92", x"9b", x"9a", x"94", 
        x"92", x"8e", x"90", x"9a", x"9a", x"8e", x"83", x"7c", x"81", x"85", x"8a", x"a0", x"db", x"f5", x"f2", 
        x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", 
        x"f2", x"f0", x"e7", x"d4", x"c1", x"ba", x"b9", x"b8", x"b9", x"ba", x"ba", x"bd", x"be", x"bb", x"ba", 
        x"b6", x"bb", x"ab", x"81", x"66", x"68", x"63", x"46", x"14", x"0a", x"17", x"28", x"35", x"49", x"4a", 
        x"47", x"47", x"4b", x"46", x"45", x"42", x"40", x"3f", x"41", x"41", x"38", x"54", x"62", x"73", x"74", 
        x"72", x"71", x"6f", x"71", x"71", x"6e", x"6e", x"70", x"70", x"70", x"6e", x"70", x"43", x"13", x"0e", 
        x"32", x"3f", x"3a", x"39", x"36", x"34", x"35", x"3b", x"35", x"1e", x"1b", x"15", x"11", x"08", x"0e", 
        x"0c", x"07", x"08", x"10", x"1b", x"1e", x"21", x"1e", x"1b", x"19", x"19", x"19", x"1c", x"19", x"0e", 
        x"07", x"09", x"0f", x"12", x"0f", x"0c", x"09", x"06", x"09", x"0d", x"0c", x"0d", x"0f", x"0e", x"0e", 
        x"0e", x"1f", x"25", x"13", x"13", x"0a", x"08", x"08", x"0d", x"0b", x"06", x"04", x"05", x"07", x"08", 
        x"04", x"0c", x"1a", x"10", x"11", x"10", x"16", x"26", x"76", x"98", x"91", x"93", x"99", x"94", x"91", 
        x"8a", x"85", x"80", x"5e", x"30", x"25", x"12", x"04", x"02", x"02", x"02", x"03", x"21", x"4f", x"50", 
        x"4e", x"4c", x"58", x"5d", x"56", x"53", x"5e", x"3c", x"23", x"23", x"23", x"23", x"1c", x"17", x"1d", 
        x"5c", x"59", x"2f", x"5d", x"81", x"89", x"6e", x"5e", x"5d", x"43", x"42", x"50", x"40", x"43", x"5b", 
        x"41", x"2f", x"34", x"41", x"55", x"41", x"3c", x"3f", x"48", x"5c", x"7b", x"87", x"65", x"5c", x"72", 
        x"88", x"75", x"50", x"4c", x"45", x"63", x"69", x"59", x"5d", x"63", x"71", x"53", x"46", x"51", x"62", 
        x"49", x"46", x"6f", x"8b", x"76", x"6b", x"5f", x"42", x"44", x"34", x"42", x"59", x"6e", x"89", x"8b", 
        x"7e", x"45", x"5a", x"7b", x"72", x"52", x"6c", x"5c", x"73", x"52", x"38", x"5a", x"3a", x"48", x"4a", 
        x"42", x"3e", x"5c", x"41", x"3a", x"5a", x"51", x"72", x"78", x"7b", x"65", x"59", x"76", x"50", x"42", 
        x"6d", x"77", x"78", x"89", x"76", x"7b", x"ab", x"8d", x"84", x"af", x"aa", x"9a", x"6d", x"7d", x"9a", 
        x"53", x"4c", x"74", x"52", x"48", x"79", x"8c", x"7f", x"85", x"98", x"9b", x"a7", x"9d", x"8b", x"98", 
        x"b4", x"a4", x"ad", x"a4", x"8c", x"8b", x"99", x"a2", x"49", x"3a", x"6d", x"72", x"6f", x"ad", x"c3", 
        x"b8", x"bb", x"c2", x"cb", x"cd", x"cd", x"d2", x"b9", x"c2", x"8b", x"5b", x"60", x"49", x"97", x"8a", 
        x"80", x"80", x"6f", x"95", x"db", x"d5", x"d4", x"d7", x"d3", x"d5", x"dd", x"ce", x"d0", x"d0", x"d0", 
        x"d0", x"d1", x"d3", x"d3", x"d0", x"d0", x"d2", x"d3", x"d3", x"d4", x"d4", x"d4", x"d4", x"d3", x"d2", 
        x"d2", x"d1", x"d1", x"d2", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d3", x"d2", x"d1", x"d0", 
        x"d1", x"d2", x"d2", x"d3", x"d3", x"d4", x"d3", x"d6", x"d3", x"d4", x"d2", x"da", x"e2", x"ac", x"7f", 
        x"67", x"68", x"6b", x"74", x"80", x"ab", x"b4", x"90", x"78", x"87", x"95", x"93", x"84", x"7d", x"7d", 
        x"7c", x"79", x"76", x"72", x"6d", x"6a", x"67", x"64", x"65", x"69", x"6a", x"67", x"6e", x"6b", x"62", 
        x"5a", x"5b", x"67", x"76", x"79", x"79", x"7e", x"85", x"83", x"7b", x"6a", x"65", x"65", x"67", x"6c", 
        x"72", x"76", x"77", x"73", x"87", x"d3", x"ce", x"9a", x"a0", x"a2", x"a4", x"a1", x"9f", x"99", x"8f", 
        x"8a", x"8c", x"90", x"90", x"8e", x"8e", x"8a", x"84", x"81", x"83", x"87", x"8c", x"91", x"92", x"8f", 
        x"8a", x"86", x"7d", x"78", x"7d", x"81", x"85", x"85", x"82", x"83", x"83", x"7c", x"7b", x"83", x"89", 
        x"a7", x"e1", x"b3", x"8e", x"94", x"93", x"91", x"91", x"92", x"99", x"99", x"99", x"9b", x"9d", x"9b", 
        x"98", x"95", x"9a", x"a0", x"a2", x"a2", x"a1", x"a1", x"9c", x"98", x"94", x"90", x"8e", x"90", x"93", 
        x"92", x"91", x"93", x"96", x"96", x"93", x"8e", x"88", x"91", x"cb", x"bb", x"79", x"73", x"70", x"72", 
        x"6a", x"65", x"64", x"68", x"6c", x"71", x"74", x"74", x"73", x"70", x"6c", x"65", x"66", x"6c", x"75", 
        x"78", x"79", x"76", x"76", x"77", x"80", x"7d", x"74", x"70", x"73", x"7b", x"7e", x"7a", x"82", x"ba", 
        x"d7", x"bd", x"ba", x"ba", x"ba", x"b9", x"bb", x"be", x"bf", x"ba", x"bb", x"bf", x"bf", x"bf", x"bb", 
        x"bd", x"bf", x"ba", x"b5", x"b8", x"ba", x"bb", x"ba", x"ba", x"bb", x"bc", x"bb", x"b8", x"b8", x"bb", 
        x"b8", x"b6", x"d4", x"ad", x"89", x"8e", x"8c", x"8a", x"86", x"89", x"8e", x"92", x"9a", x"9c", x"9a", 
        x"90", x"87", x"86", x"89", x"8b", x"91", x"92", x"8d", x"88", x"82", x"7c", x"7b", x"7a", x"7f", x"82", 
        x"82", x"aa", x"cf", x"8e", x"78", x"7c", x"7c", x"7c", x"7d", x"7e", x"82", x"82", x"82", x"7f", x"7d", 
        x"89", x"92", x"91", x"93", x"90", x"8d", x"88", x"8b", x"88", x"8c", x"8a", x"8b", x"8d", x"90", x"c6", 
        x"cb", x"8a", x"8e", x"8e", x"8e", x"8f", x"91", x"95", x"90", x"8e", x"89", x"8d", x"88", x"8e", x"96", 
        x"96", x"77", x"73", x"6f", x"6a", x"6c", x"6e", x"71", x"74", x"83", x"c1", x"bb", x"77", x"74", x"79", 
        x"78", x"78", x"77", x"76", x"76", x"76", x"7b", x"7d", x"81", x"7e", x"7b", x"79", x"7b", x"7c", x"79", 
        x"75", x"71", x"75", x"7e", x"b5", x"d2", x"97", x"8f", x"95", x"91", x"8a", x"88", x"8c", x"92", x"95", 
        x"96", x"8d", x"86", x"88", x"8d", x"90", x"91", x"8a", x"82", x"7b", x"7d", x"95", x"d4", x"f5", x"f2", 
        x"f3", x"f4", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f1", x"f1", x"f3", x"f1", 
        x"f2", x"f1", x"e8", x"d3", x"c1", x"b8", x"b9", x"bb", x"be", x"be", x"bc", x"bc", x"bc", x"ba", x"b8", 
        x"b7", x"bc", x"c2", x"a7", x"6e", x"70", x"6b", x"4f", x"17", x"0a", x"17", x"2d", x"41", x"4f", x"4c", 
        x"49", x"44", x"49", x"47", x"49", x"47", x"46", x"45", x"46", x"45", x"39", x"51", x"60", x"73", x"74", 
        x"74", x"74", x"71", x"71", x"6f", x"6d", x"6d", x"6e", x"6e", x"6d", x"6b", x"6f", x"45", x"13", x"0e", 
        x"30", x"3d", x"36", x"33", x"32", x"34", x"38", x"3e", x"37", x"21", x"18", x"11", x"11", x"09", x"11", 
        x"0e", x"06", x"09", x"10", x"19", x"1b", x"1c", x"1a", x"17", x"15", x"16", x"19", x"1f", x"1e", x"11", 
        x"07", x"09", x"12", x"16", x"10", x"0b", x"08", x"08", x"0b", x"0e", x"0d", x"0d", x"0f", x"0e", x"0e", 
        x"0d", x"1b", x"20", x"0b", x"0e", x"0b", x"09", x"07", x"0f", x"10", x"09", x"06", x"07", x"08", x"09", 
        x"06", x"0d", x"1f", x"14", x"13", x"11", x"1a", x"27", x"70", x"94", x"8f", x"92", x"98", x"95", x"92", 
        x"8d", x"86", x"7f", x"63", x"32", x"23", x"0f", x"04", x"04", x"03", x"03", x"04", x"1c", x"4d", x"4f", 
        x"4f", x"4b", x"56", x"5b", x"54", x"54", x"5f", x"3f", x"25", x"24", x"24", x"22", x"1a", x"13", x"17", 
        x"54", x"2d", x"17", x"32", x"4c", x"60", x"45", x"41", x"42", x"28", x"2a", x"51", x"40", x"43", x"42", 
        x"37", x"2e", x"3d", x"3e", x"45", x"5c", x"6f", x"92", x"a7", x"bd", x"d2", x"eb", x"ea", x"e3", x"e0", 
        x"dc", x"dd", x"e0", x"dd", x"d9", x"d7", x"d3", x"d5", x"da", x"d6", x"d1", x"cc", x"cc", x"ce", x"cb", 
        x"c9", x"c0", x"c2", x"c5", x"c9", x"d2", x"c4", x"be", x"c3", x"ab", x"9f", x"ac", x"a9", x"9d", x"a3", 
        x"ac", x"9a", x"94", x"a2", x"ad", x"ab", x"a6", x"9a", x"96", x"77", x"71", x"75", x"74", x"73", x"68", 
        x"70", x"77", x"84", x"82", x"74", x"64", x"71", x"81", x"75", x"77", x"70", x"6f", x"73", x"59", x"53", 
        x"58", x"55", x"69", x"6b", x"4b", x"49", x"8e", x"7e", x"58", x"77", x"84", x"78", x"6c", x"5e", x"7d", 
        x"57", x"53", x"7a", x"4c", x"43", x"68", x"7d", x"82", x"75", x"91", x"8b", x"7e", x"93", x"86", x"8d", 
        x"b5", x"d2", x"b3", x"93", x"a2", x"b0", x"c1", x"c0", x"45", x"2b", x"61", x"65", x"61", x"85", x"a0", 
        x"af", x"af", x"ab", x"a7", x"a6", x"b5", x"b5", x"ac", x"ab", x"81", x"53", x"4e", x"3c", x"94", x"8b", 
        x"7d", x"80", x"6c", x"93", x"da", x"d3", x"d2", x"d2", x"d3", x"d7", x"de", x"ce", x"d0", x"d2", x"d0", 
        x"cf", x"d0", x"d3", x"d3", x"d2", x"d1", x"d3", x"d3", x"d3", x"d3", x"d4", x"d4", x"d3", x"d3", x"d2", 
        x"d1", x"d2", x"d2", x"d2", x"d2", x"d2", x"d4", x"d5", x"d3", x"d2", x"d3", x"d3", x"d2", x"d1", x"d2", 
        x"d1", x"d0", x"d1", x"d3", x"d3", x"d2", x"d0", x"d5", x"d2", x"d3", x"d0", x"d8", x"e2", x"b4", x"98", 
        x"82", x"7b", x"72", x"65", x"60", x"8e", x"9d", x"80", x"65", x"5d", x"5f", x"64", x"6a", x"70", x"76", 
        x"76", x"71", x"6e", x"6e", x"6f", x"72", x"72", x"73", x"77", x"7f", x"81", x"7d", x"78", x"76", x"76", 
        x"74", x"73", x"73", x"75", x"7f", x"81", x"81", x"7b", x"73", x"72", x"73", x"6e", x"6b", x"6d", x"72", 
        x"77", x"79", x"77", x"71", x"8a", x"d9", x"cd", x"88", x"7f", x"80", x"7e", x"7e", x"76", x"71", x"72", 
        x"7b", x"85", x"8b", x"8a", x"88", x"84", x"7f", x"7d", x"81", x"88", x"90", x"92", x"94", x"94", x"93", 
        x"8e", x"89", x"8a", x"8d", x"93", x"9b", x"a0", x"a1", x"9f", x"9d", x"99", x"8e", x"85", x"89", x"90", 
        x"ab", x"e4", x"b9", x"90", x"96", x"91", x"8c", x"8e", x"8f", x"91", x"93", x"94", x"94", x"93", x"93", 
        x"90", x"87", x"83", x"82", x"82", x"83", x"83", x"82", x"84", x"8b", x"90", x"8f", x"8c", x"8c", x"90", 
        x"91", x"90", x"92", x"94", x"95", x"94", x"91", x"89", x"92", x"ce", x"c2", x"7f", x"7b", x"7b", x"82", 
        x"83", x"7e", x"7a", x"77", x"76", x"7a", x"80", x"83", x"83", x"83", x"81", x"7b", x"77", x"76", x"72", 
        x"6f", x"6e", x"6e", x"74", x"79", x"7e", x"78", x"6e", x"68", x"66", x"67", x"65", x"63", x"76", x"b7", 
        x"d4", x"bb", x"bb", x"bf", x"bd", x"b7", x"b2", x"ba", x"c1", x"c2", x"c4", x"c4", x"c0", x"bb", x"b3", 
        x"b5", x"bf", x"bf", x"bc", x"bd", x"be", x"bd", x"b9", x"b7", x"bd", x"c6", x"c8", x"c2", x"be", x"bd", 
        x"b9", x"ba", x"da", x"b1", x"82", x"82", x"83", x"84", x"85", x"8f", x"97", x"98", x"94", x"8c", x"86", 
        x"81", x"7e", x"80", x"85", x"8c", x"93", x"90", x"89", x"85", x"83", x"82", x"86", x"8b", x"93", x"91", 
        x"8c", x"ad", x"d5", x"9c", x"83", x"82", x"87", x"8a", x"89", x"88", x"83", x"83", x"88", x"82", x"7a", 
        x"88", x"92", x"8e", x"93", x"8e", x"8c", x"84", x"84", x"84", x"88", x"86", x"86", x"89", x"8a", x"bb", 
        x"c6", x"80", x"85", x"85", x"87", x"8a", x"8d", x"91", x"8b", x"8e", x"8b", x"8f", x"8a", x"8f", x"96", 
        x"98", x"7f", x"7c", x"77", x"6f", x"6d", x"6d", x"6d", x"6f", x"7c", x"bd", x"bf", x"79", x"76", x"7a", 
        x"7b", x"7b", x"7a", x"7c", x"7e", x"7c", x"7b", x"79", x"78", x"7a", x"7b", x"7d", x"80", x"81", x"80", 
        x"7d", x"75", x"77", x"7a", x"ac", x"d0", x"94", x"82", x"8b", x"94", x"93", x"8b", x"84", x"83", x"8a", 
        x"96", x"98", x"8e", x"85", x"7e", x"81", x"85", x"89", x"8d", x"87", x"7c", x"8a", x"cc", x"f5", x"f2", 
        x"f3", x"f4", x"f2", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f0", x"ef", x"f0", x"f1", x"f0", x"ee", 
        x"f0", x"f0", x"e8", x"d6", x"c6", x"be", x"bf", x"c0", x"c0", x"bc", x"b8", x"ba", x"be", x"bd", x"ba", 
        x"bf", x"be", x"bc", x"b1", x"79", x"63", x"66", x"54", x"19", x"08", x"15", x"31", x"4b", x"4f", x"4f", 
        x"4e", x"4a", x"4b", x"4a", x"4b", x"48", x"48", x"47", x"49", x"48", x"3a", x"52", x"62", x"74", x"73", 
        x"73", x"73", x"71", x"6f", x"70", x"6f", x"6b", x"6c", x"6e", x"6c", x"6c", x"74", x"4b", x"15", x"0e", 
        x"2f", x"3b", x"33", x"33", x"37", x"3b", x"3c", x"38", x"30", x"1e", x"16", x"11", x"14", x"0b", x"11", 
        x"0d", x"04", x"03", x"08", x"12", x"14", x"16", x"17", x"14", x"13", x"15", x"17", x"1d", x"1d", x"11", 
        x"09", x"09", x"11", x"14", x"0b", x"07", x"07", x"08", x"0a", x"0d", x"0c", x"0d", x"10", x"0f", x"0e", 
        x"0c", x"18", x"1e", x"06", x"09", x"06", x"06", x"07", x"12", x"14", x"0a", x"04", x"04", x"04", x"05", 
        x"07", x"0a", x"1b", x"11", x"14", x"12", x"19", x"25", x"6c", x"92", x"8e", x"91", x"97", x"95", x"92", 
        x"8d", x"88", x"82", x"69", x"36", x"29", x"14", x"05", x"04", x"05", x"04", x"05", x"18", x"4a", x"4c", 
        x"4e", x"4b", x"55", x"59", x"55", x"58", x"5c", x"3f", x"24", x"24", x"23", x"22", x"1b", x"16", x"1a", 
        x"46", x"1d", x"21", x"2b", x"3d", x"6d", x"6d", x"69", x"54", x"35", x"39", x"30", x"3c", x"4c", x"3e", 
        x"55", x"49", x"32", x"33", x"9b", x"c2", x"cc", x"d5", x"d3", x"c8", x"d5", x"ea", x"e7", x"e6", x"e8", 
        x"ea", x"ec", x"ed", x"ea", x"ed", x"eb", x"ea", x"eb", x"ed", x"eb", x"ec", x"ee", x"ec", x"ea", x"ec", 
        x"ee", x"ee", x"ec", x"ed", x"ed", x"ec", x"ef", x"f0", x"ec", x"ec", x"eb", x"eb", x"e9", x"e6", x"e8", 
        x"ec", x"ea", x"ea", x"e8", x"e8", x"ea", x"e9", x"e5", x"e7", x"e4", x"e0", x"da", x"e0", x"e0", x"dd", 
        x"df", x"da", x"d7", x"d9", x"db", x"d2", x"cd", x"cc", x"ce", x"d5", x"d2", x"ce", x"cc", x"c8", x"c9", 
        x"c2", x"c4", x"c3", x"b8", x"b5", x"b1", x"c4", x"ca", x"ae", x"ad", x"b1", x"a9", x"ad", x"a8", x"a4", 
        x"9c", x"a6", x"a7", x"8f", x"8c", x"96", x"9d", x"a2", x"98", x"ac", x"a7", x"99", x"9f", x"95", x"9e", 
        x"b8", x"c8", x"9e", x"96", x"ba", x"be", x"c4", x"bf", x"78", x"5a", x"6d", x"6e", x"71", x"9b", x"b3", 
        x"b7", x"b6", x"b2", x"bb", x"ac", x"a7", x"98", x"90", x"93", x"75", x"52", x"50", x"4a", x"88", x"82", 
        x"71", x"6e", x"62", x"90", x"d7", x"d3", x"d2", x"d1", x"cc", x"d3", x"db", x"ca", x"cb", x"cb", x"c9", 
        x"cd", x"cd", x"ce", x"ce", x"cd", x"cd", x"cf", x"d0", x"ce", x"ce", x"cd", x"ce", x"cf", x"cd", x"ce", 
        x"cf", x"d0", x"cf", x"cf", x"d0", x"d0", x"d2", x"d2", x"d1", x"d1", x"d2", x"d2", x"d2", x"d2", x"d3", 
        x"d1", x"d0", x"d1", x"d4", x"d3", x"d1", x"d0", x"d3", x"d2", x"d4", x"d1", x"d9", x"e4", x"b4", x"86", 
        x"6f", x"71", x"72", x"7e", x"86", x"9f", x"b1", x"ac", x"a5", x"a4", x"a4", x"a0", x"99", x"96", x"98", 
        x"97", x"92", x"8b", x"88", x"86", x"82", x"7f", x"7e", x"80", x"86", x"86", x"82", x"78", x"73", x"72", 
        x"72", x"72", x"72", x"73", x"77", x"78", x"76", x"70", x"69", x"66", x"62", x"63", x"66", x"6a", x"70", 
        x"78", x"7b", x"75", x"6c", x"7e", x"d0", x"d2", x"93", x"8d", x"8d", x"8a", x"86", x"7f", x"82", x"8c", 
        x"92", x"94", x"95", x"92", x"8c", x"84", x"81", x"82", x"86", x"8a", x"8c", x"8c", x"8d", x"8d", x"8a", 
        x"82", x"79", x"7d", x"82", x"85", x"87", x"87", x"86", x"84", x"81", x"7b", x"75", x"75", x"81", x"89", 
        x"a4", x"dd", x"bb", x"93", x"98", x"98", x"97", x"97", x"97", x"96", x"99", x"9a", x"99", x"98", x"99", 
        x"98", x"96", x"93", x"92", x"95", x"99", x"9a", x"99", x"9a", x"a0", x"a3", x"a0", x"98", x"95", x"98", 
        x"99", x"98", x"96", x"95", x"94", x"94", x"94", x"8f", x"97", x"d0", x"c2", x"75", x"6a", x"69", x"6f", 
        x"73", x"72", x"71", x"6d", x"68", x"66", x"68", x"69", x"66", x"67", x"6e", x"72", x"70", x"6e", x"67", 
        x"64", x"62", x"62", x"67", x"6d", x"76", x"7c", x"77", x"73", x"75", x"78", x"76", x"6f", x"79", x"b2", 
        x"d8", x"c5", x"c8", x"cd", x"cc", x"c9", x"c9", x"ca", x"c7", x"c2", x"c3", x"c6", x"c5", x"c2", x"b9", 
        x"b7", x"bb", x"ba", x"bc", x"c3", x"c6", x"c6", x"c2", x"bb", x"bb", x"be", x"c0", x"bf", x"c0", x"c5", 
        x"c7", x"be", x"d3", x"ac", x"7e", x"81", x"88", x"8f", x"92", x"95", x"94", x"90", x"8d", x"88", x"87", 
        x"8b", x"8d", x"8c", x"8c", x"8e", x"93", x"8f", x"89", x"8b", x"8e", x"91", x"97", x"94", x"90", x"89", 
        x"82", x"a5", x"d5", x"9f", x"7d", x"7c", x"81", x"84", x"83", x"81", x"81", x"83", x"86", x"80", x"76", 
        x"84", x"91", x"8e", x"91", x"8e", x"8c", x"85", x"87", x"86", x"87", x"85", x"88", x"89", x"8c", x"b9", 
        x"c7", x"81", x"85", x"86", x"8a", x"8e", x"8f", x"91", x"8b", x"8d", x"88", x"8e", x"89", x"8d", x"95", 
        x"98", x"7c", x"78", x"75", x"6d", x"6b", x"6d", x"6e", x"70", x"7d", x"bb", x"c1", x"79", x"73", x"76", 
        x"76", x"77", x"79", x"7c", x"79", x"71", x"72", x"78", x"7d", x"7e", x"7b", x"78", x"78", x"78", x"77", 
        x"7a", x"7a", x"7a", x"74", x"a4", x"d1", x"96", x"81", x"87", x"8e", x"96", x"97", x"8f", x"84", x"83", 
        x"8a", x"90", x"93", x"92", x"89", x"80", x"7b", x"7d", x"87", x"8b", x"8b", x"95", x"ce", x"f4", x"f2", 
        x"f2", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"f3", x"f2", x"f1", x"f1", x"f2", x"f2", x"f1", x"ef", 
        x"f1", x"f1", x"e9", x"d7", x"c4", x"ba", x"bd", x"bf", x"be", x"bb", x"b9", x"bb", x"be", x"bd", x"bb", 
        x"bc", x"b9", x"b7", x"c0", x"a8", x"76", x"6e", x"5d", x"1d", x"08", x"21", x"47", x"51", x"4c", x"4b", 
        x"4b", x"49", x"4a", x"49", x"47", x"46", x"48", x"46", x"47", x"49", x"3b", x"51", x"61", x"71", x"74", 
        x"72", x"75", x"74", x"72", x"72", x"71", x"6d", x"6e", x"70", x"6d", x"6d", x"74", x"50", x"19", x"11", 
        x"2e", x"3f", x"38", x"3a", x"3b", x"3c", x"39", x"37", x"32", x"23", x"1d", x"17", x"17", x"0b", x"0f", 
        x"0d", x"05", x"05", x"0a", x"14", x"17", x"18", x"1a", x"1a", x"1a", x"19", x"18", x"1c", x"1d", x"16", 
        x"15", x"20", x"1b", x"0a", x"06", x"07", x"0a", x"09", x"0a", x"0e", x"0f", x"0f", x"0f", x"0d", x"0e", 
        x"0c", x"11", x"1c", x"06", x"07", x"06", x"06", x"09", x"14", x"19", x"0d", x"03", x"03", x"03", x"05", 
        x"05", x"0a", x"1f", x"15", x"12", x"11", x"1c", x"28", x"6a", x"94", x"90", x"94", x"9a", x"97", x"92", 
        x"8c", x"88", x"86", x"6a", x"2f", x"22", x"0f", x"04", x"02", x"03", x"03", x"05", x"14", x"4a", x"4d", 
        x"4e", x"49", x"51", x"59", x"56", x"59", x"5b", x"44", x"24", x"24", x"22", x"21", x"1d", x"18", x"19", 
        x"3d", x"22", x"3f", x"62", x"66", x"82", x"5d", x"4c", x"60", x"35", x"3e", x"49", x"46", x"37", x"35", 
        x"57", x"75", x"47", x"33", x"c0", x"d3", x"cb", x"ca", x"c9", x"c1", x"d3", x"e8", x"e6", x"e7", x"e8", 
        x"e8", x"ea", x"ec", x"e9", x"e6", x"e7", x"e7", x"e8", x"e8", x"e6", x"e5", x"e5", x"e5", x"e5", x"e6", 
        x"e9", x"e9", x"e7", x"e7", x"e8", x"e8", x"e8", x"e7", x"e8", x"e9", x"e9", x"ea", x"e8", x"e8", x"e9", 
        x"e8", x"ea", x"ea", x"eb", x"ea", x"ea", x"ea", x"e4", x"e8", x"ed", x"ec", x"ed", x"ed", x"ee", x"ee", 
        x"ee", x"ed", x"ed", x"ef", x"f1", x"e7", x"ee", x"f2", x"ed", x"f0", x"f3", x"f0", x"f0", x"f2", x"f3", 
        x"f3", x"f2", x"f0", x"f2", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", 
        x"f1", x"ef", x"ed", x"ec", x"ee", x"ed", x"ea", x"e9", x"e8", x"e5", x"e4", x"e4", x"e0", x"dd", x"de", 
        x"e1", x"e4", x"de", x"e3", x"e9", x"e9", x"e5", x"de", x"d5", x"d0", x"cf", x"c9", x"c4", x"d8", x"dc", 
        x"d2", x"d2", x"d0", x"d7", x"d8", x"d1", x"c6", x"c4", x"cb", x"b6", x"a1", x"a2", x"a1", x"b9", x"b8", 
        x"a9", x"a7", x"9f", x"bb", x"e2", x"dd", x"de", x"da", x"d4", x"d9", x"e1", x"d4", x"d4", x"d3", x"d2", 
        x"d7", x"d6", x"d5", x"d6", x"d5", x"d2", x"d3", x"d6", x"d4", x"d3", x"cf", x"d1", x"d4", x"cf", x"cf", 
        x"d1", x"d0", x"cf", x"d0", x"d1", x"d2", x"d2", x"d0", x"d0", x"d0", x"d1", x"d2", x"d2", x"d3", x"d1", 
        x"cf", x"ce", x"cf", x"d0", x"d0", x"cf", x"d1", x"d0", x"cf", x"ce", x"cc", x"d7", x"e4", x"b4", x"94", 
        x"95", x"9b", x"95", x"98", x"9d", x"ba", x"d1", x"d3", x"da", x"e1", x"e2", x"dd", x"d4", x"cc", x"ca", 
        x"cb", x"cd", x"cd", x"cb", x"ca", x"c6", x"bf", x"ba", x"ba", x"be", x"bf", x"bf", x"bd", x"b8", x"b5", 
        x"b3", x"ae", x"ab", x"ab", x"ad", x"af", x"af", x"ab", x"a8", x"a3", x"9d", x"98", x"97", x"96", x"97", 
        x"9b", x"9d", x"97", x"90", x"9a", x"d4", x"d4", x"a1", x"9c", x"a1", x"9c", x"91", x"86", x"83", x"84", 
        x"81", x"81", x"87", x"87", x"7e", x"75", x"75", x"7a", x"80", x"84", x"88", x"8d", x"92", x"93", x"8c", 
        x"83", x"7c", x"7c", x"80", x"85", x"87", x"88", x"8b", x"90", x"91", x"8d", x"89", x"82", x"88", x"8d", 
        x"a9", x"dd", x"bd", x"95", x"98", x"96", x"93", x"8d", x"88", x"88", x"8d", x"8f", x"8e", x"8e", x"8d", 
        x"8a", x"8c", x"87", x"83", x"83", x"87", x"8b", x"8b", x"8b", x"8f", x"94", x"92", x"8b", x"85", x"82", 
        x"86", x"8b", x"8f", x"92", x"94", x"95", x"96", x"96", x"9b", x"ce", x"c7", x"7b", x"6c", x"6b", x"6e", 
        x"71", x"79", x"80", x"84", x"84", x"82", x"7f", x"78", x"72", x"70", x"73", x"78", x"7d", x"83", x"83", 
        x"81", x"82", x"80", x"79", x"79", x"84", x"83", x"7a", x"72", x"76", x"7e", x"80", x"79", x"82", x"b5", 
        x"d8", x"c2", x"c0", x"c1", x"c1", x"c2", x"c8", x"c8", x"c3", x"bc", x"b9", x"b9", x"b9", x"b9", x"b9", 
        x"c0", x"c9", x"c9", x"c8", x"cb", x"cb", x"c9", x"c9", x"c9", x"ca", x"cd", x"ce", x"ca", x"c8", x"ca", 
        x"ce", x"c6", x"d8", x"b5", x"8e", x"93", x"95", x"96", x"95", x"91", x"8c", x"89", x"89", x"8b", x"8e", 
        x"8f", x"8d", x"89", x"85", x"80", x"82", x"84", x"84", x"8b", x"95", x"95", x"91", x"87", x"7d", x"7a", 
        x"77", x"9e", x"d4", x"9f", x"76", x"7b", x"81", x"84", x"86", x"86", x"8a", x"88", x"86", x"82", x"7c", 
        x"88", x"95", x"91", x"92", x"92", x"8f", x"89", x"8f", x"8a", x"8b", x"8d", x"8f", x"8e", x"91", x"bb", 
        x"ce", x"85", x"88", x"88", x"8c", x"8e", x"8e", x"8f", x"8b", x"8d", x"86", x"8c", x"87", x"8a", x"91", 
        x"95", x"7a", x"76", x"73", x"6b", x"69", x"6d", x"6e", x"6c", x"79", x"b8", x"c5", x"7b", x"74", x"7a", 
        x"7b", x"7e", x"7d", x"79", x"6d", x"62", x"66", x"70", x"76", x"79", x"78", x"76", x"75", x"73", x"71", 
        x"71", x"75", x"74", x"6e", x"a1", x"d3", x"a0", x"89", x"87", x"85", x"8b", x"95", x"98", x"8f", x"87", 
        x"87", x"87", x"8d", x"90", x"8e", x"8a", x"81", x"7b", x"7c", x"82", x"8b", x"99", x"cf", x"f4", x"f3", 
        x"f3", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f0", x"ef", 
        x"ef", x"f2", x"eb", x"db", x"c6", x"b8", x"bb", x"bd", x"bd", x"ba", x"ba", x"bb", x"bd", x"bc", x"bd", 
        x"bf", x"c0", x"c1", x"c5", x"ba", x"88", x"6b", x"60", x"21", x"08", x"2b", x"52", x"4f", x"48", x"4a", 
        x"4a", x"47", x"4a", x"49", x"4a", x"4a", x"4d", x"4a", x"49", x"4d", x"3d", x"51", x"62", x"70", x"7a", 
        x"73", x"77", x"75", x"72", x"6e", x"6c", x"6c", x"70", x"70", x"6d", x"6b", x"71", x"54", x"1a", x"0f", 
        x"25", x"3a", x"38", x"3b", x"38", x"36", x"35", x"39", x"38", x"28", x"1e", x"19", x"15", x"0c", x"16", 
        x"18", x"0b", x"06", x"0a", x"16", x"19", x"19", x"1d", x"1f", x"1d", x"1d", x"20", x"25", x"25", x"1d", 
        x"20", x"3a", x"2d", x"08", x"07", x"0b", x"0d", x"0c", x"0d", x"10", x"11", x"10", x"0d", x"0b", x"0c", 
        x"0b", x"0f", x"1c", x"09", x"09", x"0a", x"08", x"09", x"13", x"1c", x"10", x"03", x"03", x"03", x"05", 
        x"07", x"0a", x"20", x"17", x"0f", x"0d", x"16", x"1f", x"64", x"97", x"94", x"94", x"9a", x"97", x"92", 
        x"8b", x"88", x"89", x"72", x"36", x"28", x"14", x"08", x"05", x"05", x"05", x"07", x"12", x"4a", x"4f", 
        x"4e", x"47", x"4f", x"5b", x"56", x"56", x"5c", x"4b", x"24", x"24", x"21", x"1d", x"1a", x"16", x"17", 
        x"37", x"23", x"35", x"40", x"3d", x"6c", x"5d", x"30", x"43", x"30", x"30", x"47", x"4c", x"57", x"3d", 
        x"41", x"57", x"39", x"33", x"b6", x"cf", x"c9", x"c7", x"c8", x"c4", x"d3", x"e5", x"e8", x"ed", x"eb", 
        x"ea", x"ec", x"ed", x"ec", x"e9", x"e8", x"e9", x"e9", x"e9", x"e8", x"e8", x"e7", x"e7", x"e7", x"e9", 
        x"eb", x"eb", x"e9", x"e9", x"ea", x"ea", x"e8", x"e7", x"ea", x"ed", x"ed", x"eb", x"e9", x"ec", x"ec", 
        x"e9", x"eb", x"ea", x"e9", x"e9", x"e8", x"e8", x"e6", x"e9", x"eb", x"eb", x"ea", x"ea", x"eb", x"ec", 
        x"eb", x"e9", x"ea", x"ea", x"e7", x"dc", x"e3", x"ea", x"e8", x"e9", x"ea", x"e9", x"e9", x"ea", x"eb", 
        x"eb", x"ea", x"ea", x"e9", x"e9", x"e9", x"eb", x"ed", x"ee", x"ee", x"ed", x"eb", x"eb", x"ea", x"ea", 
        x"eb", x"ec", x"ec", x"ec", x"eb", x"e9", x"e9", x"ec", x"ee", x"ee", x"ef", x"ed", x"ee", x"ed", x"ed", 
        x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", x"ef", x"ed", x"ee", x"f0", x"f1", x"f2", x"ed", x"ed", x"ef", 
        x"f0", x"f2", x"f0", x"ef", x"ef", x"f3", x"f2", x"f0", x"f0", x"ed", x"f0", x"f2", x"ee", x"f1", x"ec", 
        x"ec", x"f2", x"ed", x"ec", x"ed", x"eb", x"f2", x"ef", x"ec", x"ed", x"f1", x"eb", x"ef", x"ef", x"ec", 
        x"eb", x"eb", x"ed", x"ef", x"ec", x"eb", x"ee", x"ed", x"ea", x"ea", x"e8", x"eb", x"ed", x"e9", x"e8", 
        x"ea", x"ea", x"ea", x"ea", x"ea", x"ea", x"eb", x"ea", x"e9", x"e8", x"e8", x"e9", x"e9", x"e9", x"e6", 
        x"e5", x"e4", x"e4", x"e4", x"e3", x"e2", x"e2", x"e3", x"e3", x"e4", x"e0", x"e5", x"ee", x"e3", x"dc", 
        x"d6", x"cd", x"c6", x"c7", x"c6", x"d7", x"e3", x"dd", x"dc", x"e1", x"e6", x"e9", x"ea", x"eb", x"ed", 
        x"ef", x"ee", x"ed", x"ec", x"ec", x"ee", x"ec", x"ec", x"ee", x"f0", x"f0", x"ee", x"ec", x"e8", x"e6", 
        x"e6", x"e5", x"e3", x"e2", x"e3", x"e5", x"e7", x"e5", x"e6", x"e6", x"e2", x"dc", x"d9", x"d8", x"d5", 
        x"d4", x"d8", x"db", x"d8", x"d6", x"e3", x"de", x"cf", x"d3", x"d0", x"cf", x"d3", x"d3", x"d4", x"cf", 
        x"c6", x"c3", x"c8", x"c7", x"c4", x"c1", x"c0", x"c0", x"be", x"ba", x"b3", x"b5", x"bc", x"c0", x"be", 
        x"b9", x"b5", x"b4", x"b3", x"b0", x"ac", x"a9", x"ac", x"b1", x"b2", x"af", x"ad", x"a4", x"9c", x"99", 
        x"af", x"da", x"be", x"96", x"9c", x"9c", x"9b", x"97", x"93", x"94", x"95", x"93", x"95", x"9b", x"a3", 
        x"a5", x"a2", x"9c", x"94", x"90", x"8f", x"8f", x"8e", x"91", x"98", x"9f", x"a3", x"a1", x"9d", x"9a", 
        x"94", x"90", x"8e", x"8d", x"8d", x"8d", x"8d", x"8c", x"92", x"c7", x"c8", x"82", x"70", x"6a", x"66", 
        x"64", x"68", x"6e", x"74", x"77", x"78", x"77", x"71", x"6e", x"6c", x"67", x"61", x"64", x"6b", x"73", 
        x"75", x"78", x"7b", x"77", x"76", x"7d", x"77", x"6e", x"68", x"68", x"6a", x"6b", x"67", x"73", x"ab", 
        x"da", x"cb", x"c9", x"c7", x"c2", x"c1", x"c2", x"c5", x"c4", x"c4", x"c9", x"ce", x"ce", x"c6", x"c4", 
        x"c6", x"c8", x"c9", x"c8", x"c7", x"c9", x"c9", x"c7", x"c3", x"c1", x"c0", x"c2", x"c0", x"c1", x"bc", 
        x"bb", x"bb", x"d2", x"b0", x"85", x"8a", x"84", x"80", x"7f", x"7f", x"80", x"83", x"89", x"8c", x"8c", 
        x"86", x"80", x"80", x"82", x"83", x"88", x"92", x"96", x"9a", x"9b", x"94", x"8a", x"87", x"83", x"82", 
        x"7f", x"a2", x"d8", x"af", x"85", x"88", x"8f", x"8e", x"8e", x"8d", x"8d", x"8c", x"8c", x"87", x"7d", 
        x"83", x"89", x"88", x"8e", x"8f", x"8d", x"88", x"8b", x"87", x"8b", x"8b", x"8c", x"86", x"88", x"b5", 
        x"d2", x"89", x"8a", x"88", x"8b", x"8b", x"8c", x"8e", x"8b", x"90", x"8a", x"8e", x"89", x"8b", x"92", 
        x"95", x"7c", x"78", x"74", x"6d", x"6d", x"71", x"71", x"72", x"7b", x"b4", x"cb", x"84", x"7d", x"80", 
        x"7b", x"79", x"79", x"78", x"75", x"71", x"6f", x"71", x"73", x"78", x"7a", x"7a", x"7a", x"7a", x"77", 
        x"75", x"74", x"73", x"79", x"a9", x"d3", x"a3", x"96", x"95", x"8b", x"85", x"88", x"8e", x"90", x"8f", 
        x"8d", x"87", x"83", x"7e", x"83", x"8d", x"8e", x"8f", x"8d", x"86", x"80", x"89", x"c6", x"f3", x"f2", 
        x"f2", x"f2", x"f3", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ee", 
        x"ee", x"f0", x"e8", x"d9", x"c7", x"bb", x"be", x"c0", x"c0", x"bd", x"bc", x"bd", x"bf", x"bd", x"b9", 
        x"b8", x"ba", x"ba", x"bb", x"bf", x"ad", x"7a", x"60", x"24", x"0a", x"2d", x"50", x"4c", x"4a", x"4c", 
        x"4a", x"45", x"45", x"45", x"48", x"45", x"45", x"43", x"47", x"49", x"39", x"4e", x"61", x"70", x"7c", 
        x"75", x"76", x"73", x"72", x"71", x"6f", x"6e", x"6f", x"70", x"6d", x"6b", x"71", x"59", x"1f", x"14", 
        x"28", x"37", x"37", x"32", x"33", x"34", x"35", x"38", x"36", x"24", x"17", x"14", x"14", x"13", x"26", 
        x"2a", x"13", x"06", x"0a", x"1a", x"1e", x"1f", x"21", x"24", x"20", x"21", x"24", x"26", x"22", x"1b", 
        x"1e", x"3b", x"35", x"0c", x"08", x"0b", x"0c", x"0a", x"0d", x"0e", x"0b", x"0a", x"0b", x"0b", x"09", 
        x"06", x"0d", x"1b", x"0a", x"08", x"08", x"08", x"0a", x"0b", x"14", x"0f", x"05", x"05", x"05", x"07", 
        x"09", x"08", x"1d", x"18", x"10", x"0c", x"14", x"1f", x"62", x"9b", x"99", x"98", x"9c", x"98", x"94", 
        x"90", x"8b", x"84", x"70", x"3a", x"2c", x"18", x"07", x"04", x"05", x"05", x"05", x"0c", x"42", x"4d", 
        x"4b", x"47", x"51", x"5c", x"54", x"50", x"57", x"47", x"20", x"22", x"22", x"1e", x"19", x"13", x"17", 
        x"33", x"29", x"29", x"2e", x"3d", x"62", x"4f", x"5e", x"4f", x"45", x"56", x"2f", x"32", x"59", x"48", 
        x"29", x"30", x"31", x"35", x"b7", x"ce", x"c5", x"c4", x"c6", x"c7", x"d5", x"e4", x"e5", x"ea", x"e9", 
        x"e9", x"e9", x"ea", x"ec", x"ec", x"ea", x"ec", x"eb", x"e9", x"e9", x"e8", x"e7", x"e5", x"e6", x"e8", 
        x"ea", x"eb", x"ea", x"ea", x"eb", x"ed", x"ec", x"e9", x"eb", x"ed", x"ed", x"ec", x"ea", x"eb", x"eb", 
        x"e7", x"ed", x"e9", x"e9", x"eb", x"e9", x"e9", x"e8", x"e9", x"ea", x"e8", x"e8", x"e9", x"ea", x"ea", 
        x"ea", x"ea", x"ec", x"ed", x"e6", x"dd", x"e3", x"ea", x"e9", x"e9", x"e9", x"e9", x"ea", x"ea", x"eb", 
        x"eb", x"ec", x"ed", x"eb", x"ea", x"eb", x"ec", x"ed", x"ed", x"ec", x"ec", x"ec", x"ec", x"ec", x"ed", 
        x"ed", x"ed", x"ec", x"ea", x"eb", x"eb", x"ea", x"eb", x"eb", x"ec", x"ec", x"ec", x"ee", x"ec", x"e8", 
        x"ea", x"ed", x"ed", x"e9", x"e9", x"ed", x"ec", x"ea", x"eb", x"ed", x"ec", x"ee", x"ed", x"ea", x"eb", 
        x"ef", x"ef", x"f0", x"f0", x"ed", x"eb", x"ed", x"ed", x"ed", x"ee", x"ee", x"eb", x"ee", x"ee", x"ea", 
        x"eb", x"e7", x"e9", x"ee", x"f0", x"ed", x"ec", x"ef", x"ef", x"ee", x"f0", x"ed", x"f1", x"f0", x"ee", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"f0", x"ec", x"ec", x"f0", x"f1", x"f1", x"f2", x"f0", x"ef", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"ee", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"f1", x"f0", x"ee", x"ee", x"ee", x"f2", 
        x"ef", x"e8", x"e7", x"e7", x"e1", x"e9", x"ee", x"e8", x"e6", x"e8", x"ea", x"ec", x"ed", x"eb", x"ea", 
        x"ed", x"ee", x"ec", x"ea", x"ec", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", x"ed", x"f1", x"ef", x"ee", 
        x"f0", x"f1", x"f0", x"ee", x"ef", x"f1", x"f1", x"f0", x"f1", x"f3", x"f0", x"f0", x"f1", x"f2", x"ef", 
        x"ee", x"ee", x"ef", x"ee", x"ea", x"e6", x"e3", x"e3", x"e6", x"e5", x"e6", x"e9", x"eb", x"ec", x"eb", 
        x"e7", x"e6", x"e7", x"e6", x"e6", x"e7", x"e9", x"e9", x"e9", x"e7", x"e3", x"e3", x"e5", x"e5", x"e3", 
        x"e2", x"e2", x"e3", x"e4", x"e3", x"e0", x"de", x"dd", x"df", x"e0", x"de", x"df", x"dc", x"de", x"dd", 
        x"de", x"e9", x"da", x"ca", x"ce", x"cb", x"ca", x"cb", x"cb", x"cb", x"c8", x"c2", x"c2", x"c5", x"c9", 
        x"cb", x"ca", x"c7", x"c4", x"c2", x"c0", x"bd", x"ba", x"b4", x"b4", x"b7", x"ba", x"ba", x"ba", x"b9", 
        x"b4", x"b0", x"af", x"af", x"ae", x"ac", x"a9", x"a7", x"aa", x"cd", x"c9", x"90", x"80", x"80", x"83", 
        x"86", x"87", x"89", x"8c", x"8d", x"8c", x"8a", x"86", x"82", x"7f", x"7c", x"78", x"77", x"79", x"7c", 
        x"7d", x"81", x"84", x"82", x"80", x"83", x"80", x"7c", x"79", x"76", x"74", x"71", x"6d", x"77", x"ad", 
        x"d8", x"c3", x"bd", x"c0", x"c0", x"c2", x"c0", x"c0", x"bc", x"b9", x"be", x"c3", x"c5", x"c5", x"c2", 
        x"c0", x"bf", x"c0", x"bc", x"b8", x"b9", x"bc", x"be", x"bc", x"ba", x"b7", x"b8", x"b7", x"bd", x"ba", 
        x"bc", x"bf", x"d0", x"af", x"7d", x"81", x"81", x"86", x"8c", x"93", x"98", x"99", x"96", x"90", x"8b", 
        x"89", x"89", x"87", x"89", x"93", x"99", x"a1", x"9d", x"95", x"8f", x"88", x"83", x"81", x"7d", x"7e", 
        x"7e", x"9e", x"d6", x"ad", x"7d", x"7e", x"88", x"8a", x"8c", x"8d", x"8c", x"8c", x"8e", x"8a", x"7f", 
        x"83", x"8c", x"8c", x"90", x"92", x"90", x"8b", x"8e", x"8c", x"8f", x"8e", x"8f", x"8a", x"8c", x"b3", 
        x"d4", x"91", x"8d", x"8b", x"8e", x"8f", x"8f", x"92", x"8f", x"90", x"8b", x"8f", x"8a", x"8c", x"91", 
        x"93", x"7d", x"77", x"73", x"6f", x"6f", x"70", x"6e", x"6c", x"74", x"af", x"cd", x"8c", x"7f", x"82", 
        x"7f", x"7b", x"79", x"7a", x"77", x"7a", x"8b", x"92", x"76", x"78", x"79", x"78", x"78", x"77", x"76", 
        x"7e", x"7b", x"75", x"78", x"a4", x"cf", x"9d", x"90", x"96", x"92", x"88", x"81", x"81", x"84", x"8c", 
        x"90", x"91", x"8f", x"83", x"80", x"84", x"84", x"8e", x"93", x"90", x"8e", x"95", x"c8", x"f1", x"f0", 
        x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f0", x"ef", x"eb", 
        x"ec", x"f0", x"e8", x"d9", x"c9", x"bc", x"c0", x"c3", x"c3", x"c0", x"be", x"be", x"be", x"bb", x"b9", 
        x"bb", x"c0", x"c2", x"c2", x"c5", x"ba", x"90", x"67", x"2a", x"13", x"36", x"58", x"51", x"4f", x"4e", 
        x"49", x"44", x"46", x"49", x"47", x"46", x"47", x"47", x"4b", x"4c", x"3e", x"50", x"63", x"70", x"7b", 
        x"76", x"78", x"76", x"75", x"74", x"72", x"72", x"73", x"72", x"71", x"6e", x"74", x"5d", x"27", x"25", 
        x"3a", x"38", x"36", x"34", x"36", x"37", x"36", x"39", x"36", x"24", x"17", x"1a", x"19", x"17", x"29", 
        x"2f", x"14", x"0b", x"11", x"1f", x"21", x"1e", x"1e", x"1f", x"1c", x"1e", x"1f", x"20", x"1e", x"1a", 
        x"1d", x"3b", x"3b", x"10", x"09", x"0b", x"0b", x"0a", x"0b", x"0d", x"0a", x"08", x"0a", x"0a", x"07", 
        x"03", x"0c", x"1b", x"0c", x"07", x"07", x"08", x"0a", x"0b", x"16", x"14", x"0b", x"07", x"05", x"07", 
        x"0a", x"08", x"1c", x"1a", x"12", x"0d", x"13", x"22", x"5e", x"94", x"93", x"94", x"9c", x"9a", x"97", 
        x"92", x"8c", x"85", x"76", x"3f", x"2b", x"1b", x"07", x"02", x"06", x"06", x"06", x"0b", x"40", x"4e", 
        x"4c", x"49", x"4e", x"57", x"52", x"50", x"57", x"4b", x"25", x"26", x"26", x"22", x"1d", x"15", x"16", 
        x"49", x"3b", x"37", x"2a", x"37", x"5e", x"63", x"73", x"6f", x"4c", x"43", x"41", x"71", x"7c", x"42", 
        x"2d", x"29", x"30", x"35", x"b4", x"cf", x"c7", x"c9", x"cb", x"ce", x"db", x"eb", x"e9", x"ea", x"eb", 
        x"ed", x"ef", x"ed", x"ef", x"f0", x"ea", x"ee", x"ee", x"ed", x"ed", x"ee", x"ed", x"eb", x"e9", x"ea", 
        x"ec", x"ed", x"ed", x"ee", x"ee", x"ea", x"eb", x"eb", x"ed", x"eb", x"ea", x"ea", x"ea", x"eb", x"eb", 
        x"e7", x"ec", x"e6", x"e6", x"e9", x"eb", x"ea", x"ea", x"ea", x"ea", x"e9", x"e9", x"e9", x"eb", x"ed", 
        x"ec", x"ec", x"ee", x"ef", x"ed", x"e8", x"eb", x"ee", x"eb", x"ea", x"eb", x"eb", x"eb", x"ea", x"ea", 
        x"ea", x"eb", x"eb", x"eb", x"eb", x"ec", x"ed", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", 
        x"ef", x"ef", x"ed", x"ec", x"ea", x"e9", x"e8", x"ea", x"ed", x"ee", x"eb", x"ec", x"ec", x"ed", x"ed", 
        x"ed", x"ee", x"ef", x"ec", x"eb", x"ec", x"ee", x"ee", x"ee", x"ec", x"ed", x"ea", x"eb", x"ed", x"eb", 
        x"ed", x"ed", x"ed", x"ef", x"ed", x"eb", x"ee", x"ed", x"eb", x"eb", x"ed", x"eb", x"ed", x"eb", x"ed", 
        x"f1", x"ee", x"ee", x"f0", x"f1", x"ef", x"eb", x"ef", x"ec", x"ec", x"ee", x"ed", x"ed", x"ea", x"eb", 
        x"ed", x"ed", x"ed", x"ee", x"f0", x"ee", x"e9", x"e1", x"e5", x"ef", x"f1", x"ed", x"ec", x"ed", x"ed", 
        x"ed", x"ed", x"ed", x"ed", x"ed", x"ec", x"ed", x"ee", x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ec", 
        x"ec", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", x"ef", x"ee", x"ef", x"f2", x"ed", x"f0", 
        x"f1", x"f0", x"f3", x"ec", x"de", x"e7", x"f0", x"ee", x"f0", x"f3", x"f1", x"ef", x"ef", x"eb", x"e6", 
        x"ea", x"f0", x"f0", x"ee", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"ef", x"f0", x"ef", x"ed", x"ed", 
        x"ef", x"f2", x"f2", x"f0", x"ef", x"f0", x"ef", x"ed", x"ed", x"ef", x"ed", x"ef", x"f1", x"ef", x"ef", 
        x"ee", x"ed", x"ec", x"ed", x"ee", x"eb", x"ed", x"eb", x"e9", x"ed", x"ed", x"f0", x"ef", x"ee", x"ef", 
        x"f1", x"f1", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f1", x"f0", x"f0", x"f0", x"ee", x"ed", x"ec", x"ed", x"ee", x"ed", x"ef", x"f1", x"ef", x"ec", 
        x"ec", x"f2", x"ed", x"ea", x"e7", x"e6", x"ea", x"e9", x"ec", x"eb", x"ea", x"eb", x"ec", x"ed", x"ea", 
        x"e8", x"e7", x"e8", x"e8", x"ea", x"eb", x"ea", x"e8", x"e8", x"e7", x"e6", x"e6", x"e6", x"e7", x"e7", 
        x"e7", x"e5", x"e4", x"e4", x"e2", x"df", x"db", x"da", x"d5", x"dc", x"e2", x"d4", x"d6", x"d3", x"d2", 
        x"d2", x"d1", x"d1", x"d2", x"d2", x"d0", x"ce", x"cd", x"c9", x"c6", x"c5", x"c5", x"c3", x"bf", x"be", 
        x"be", x"c0", x"c3", x"c3", x"c2", x"c3", x"c4", x"c2", x"bd", x"b4", x"ac", x"a7", x"a5", x"a3", x"be", 
        x"db", x"cb", x"c5", x"ca", x"cb", x"d2", x"da", x"d9", x"d4", x"d0", x"d0", x"d0", x"ce", x"ce", x"d1", 
        x"d4", x"d8", x"da", x"d6", x"cc", x"c7", x"c7", x"c8", x"c7", x"c6", x"c7", x"cb", x"cf", x"d4", x"cc", 
        x"c9", x"c5", x"ca", x"b3", x"89", x"88", x"8b", x"8f", x"91", x"90", x"8d", x"89", x"84", x"7f", x"7c", 
        x"7c", x"80", x"83", x"87", x"8a", x"89", x"8b", x"84", x"7d", x"7c", x"7c", x"7c", x"7a", x"7a", x"7f", 
        x"81", x"9b", x"d0", x"b2", x"83", x"7b", x"7e", x"7e", x"83", x"87", x"8b", x"90", x"95", x"95", x"8c", 
        x"89", x"8a", x"88", x"8b", x"8d", x"8d", x"8e", x"92", x"95", x"9c", x"98", x"95", x"90", x"90", x"bc", 
        x"dc", x"8e", x"8a", x"89", x"8d", x"8d", x"8c", x"8d", x"8a", x"8b", x"88", x"8c", x"8a", x"8e", x"92", 
        x"92", x"7d", x"74", x"6d", x"68", x"68", x"69", x"67", x"67", x"70", x"ae", x"cd", x"87", x"75", x"7f", 
        x"7f", x"7c", x"7a", x"79", x"74", x"79", x"92", x"a0", x"81", x"82", x"81", x"7e", x"7e", x"7d", x"7a", 
        x"77", x"7b", x"7c", x"76", x"9c", x"d2", x"a1", x"87", x"8f", x"97", x"93", x"8b", x"86", x"84", x"86", 
        x"8a", x"96", x"9e", x"96", x"8e", x"87", x"7d", x"7e", x"83", x"89", x"94", x"9f", x"ca", x"ef", x"ef", 
        x"f0", x"f0", x"f1", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f3", x"f1", 
        x"f1", x"f3", x"ea", x"da", x"c7", x"bb", x"bd", x"be", x"bd", x"bd", x"bf", x"c3", x"c6", x"c5", x"bf", 
        x"b8", x"b5", x"b5", x"b5", x"b7", x"b9", x"ad", x"72", x"26", x"10", x"30", x"4e", x"48", x"4b", x"4c", 
        x"4a", x"46", x"48", x"4a", x"45", x"47", x"49", x"49", x"4b", x"4c", x"43", x"4c", x"5e", x"6a", x"76", 
        x"71", x"72", x"71", x"72", x"72", x"71", x"70", x"71", x"70", x"6f", x"6d", x"72", x"5c", x"2a", x"30", 
        x"47", x"39", x"37", x"3c", x"3b", x"38", x"33", x"33", x"30", x"1f", x"1a", x"1d", x"1b", x"18", x"27", 
        x"30", x"15", x"06", x"0b", x"18", x"1a", x"17", x"18", x"1b", x"16", x"14", x"14", x"17", x"1a", x"19", 
        x"19", x"38", x"40", x"14", x"0d", x"0f", x"0f", x"0e", x"0d", x"0d", x"0c", x"0a", x"09", x"07", x"06", 
        x"04", x"0b", x"1b", x"0e", x"07", x"06", x"07", x"0a", x"0d", x"16", x"17", x"0d", x"07", x"03", x"03", 
        x"08", x"06", x"18", x"1a", x"11", x"0d", x"11", x"21", x"5a", x"93", x"91", x"8c", x"97", x"99", x"9a", 
        x"94", x"8b", x"84", x"79", x"43", x"2a", x"1e", x"0c", x"06", x"09", x"09", x"08", x"0d", x"40", x"51", 
        x"4e", x"49", x"4b", x"53", x"50", x"51", x"53", x"4b", x"26", x"25", x"23", x"1f", x"1d", x"16", x"14", 
        x"51", x"2d", x"43", x"2e", x"47", x"83", x"5e", x"4e", x"37", x"26", x"22", x"4d", x"8b", x"96", x"57", 
        x"3b", x"2e", x"36", x"58", x"c7", x"d2", x"c4", x"c4", x"bd", x"af", x"ab", x"bc", x"bb", x"ba", x"bc", 
        x"ba", x"b8", x"b3", x"bc", x"c8", x"c5", x"c2", x"c1", x"c1", x"c2", x"c3", x"c3", x"c3", x"c4", x"c5", 
        x"c7", x"c8", x"c9", x"ca", x"c9", x"c8", x"cd", x"d2", x"d4", x"d2", x"d3", x"d7", x"dc", x"d9", x"db", 
        x"db", x"de", x"d8", x"dc", x"dd", x"de", x"da", x"dd", x"df", x"e1", x"e2", x"e0", x"e2", x"e5", x"e7", 
        x"e6", x"e5", x"e4", x"e4", x"e7", x"e6", x"e8", x"eb", x"ea", x"e9", x"eb", x"eb", x"ea", x"e9", x"e8", 
        x"e8", x"e8", x"e9", x"ea", x"ea", x"ea", x"e9", x"e8", x"e8", x"e9", x"ea", x"ea", x"ea", x"ea", x"ea", 
        x"ec", x"ed", x"ec", x"ea", x"e8", x"ea", x"ec", x"eb", x"ea", x"eb", x"ed", x"ee", x"ee", x"ec", x"ee", 
        x"ed", x"e8", x"ec", x"ed", x"ed", x"ed", x"ee", x"ee", x"ec", x"ea", x"ee", x"ec", x"ec", x"f0", x"f0", 
        x"f0", x"ee", x"ea", x"ee", x"ee", x"ed", x"f2", x"f0", x"ee", x"ef", x"ef", x"f1", x"f1", x"ee", x"f0", 
        x"f1", x"f3", x"ef", x"ed", x"ed", x"eb", x"eb", x"ef", x"ef", x"f1", x"f2", x"f1", x"ef", x"ee", x"ef", 
        x"ee", x"ed", x"ec", x"ed", x"f0", x"f2", x"ee", x"e3", x"e6", x"ef", x"f2", x"ef", x"ee", x"f1", x"f0", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", x"ee", x"ee", x"ee", x"ee", x"ed", 
        x"ef", x"ef", x"ef", x"ee", x"ed", x"ec", x"ed", x"ec", x"ea", x"ed", x"ee", x"ed", x"ed", x"ee", x"ec", 
        x"ec", x"ee", x"ef", x"ec", x"df", x"e7", x"f1", x"ec", x"ee", x"f0", x"ed", x"ed", x"ef", x"ed", x"e6", 
        x"ea", x"f0", x"f0", x"ef", x"f0", x"ef", x"f0", x"f1", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ee", 
        x"ee", x"f0", x"f0", x"ee", x"ef", x"f1", x"f1", x"ee", x"ef", x"f1", x"ef", x"ef", x"ee", x"ed", x"ef", 
        x"f0", x"ef", x"ee", x"f0", x"ee", x"eb", x"ef", x"f1", x"f0", x"f4", x"f0", x"f2", x"f2", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f1", x"ef", x"ef", x"ef", x"ee", x"ed", 
        x"ef", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", 
        x"ee", x"ec", x"ee", x"f0", x"ef", x"f2", x"f0", x"ed", x"f1", x"f1", x"ef", x"ee", x"ef", x"f0", x"f0", 
        x"f1", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"f0", x"f2", x"f1", x"f1", x"ef", x"ed", x"ea", x"eb", x"eb", x"ec", x"f0", x"f1", x"f0", x"ec", x"ee", 
        x"ed", x"ee", x"ef", x"f1", x"f2", x"f2", x"f1", x"f1", x"f1", x"f0", x"ee", x"ef", x"ee", x"ec", x"ee", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f2", x"f2", x"f1", x"f1", x"ef", x"ec", x"ec", x"ed", x"ea", x"ed", 
        x"ed", x"e8", x"e7", x"ea", x"e9", x"ee", x"ee", x"ed", x"e9", x"e5", x"e5", x"e5", x"e3", x"e5", x"e7", 
        x"e7", x"e8", x"ea", x"e9", x"e3", x"df", x"de", x"de", x"dd", x"de", x"e1", x"e5", x"e7", x"e7", x"e1", 
        x"de", x"db", x"df", x"da", x"c8", x"c8", x"c8", x"c8", x"c8", x"c8", x"c6", x"c3", x"c0", x"bf", x"bf", 
        x"bf", x"c1", x"c2", x"c3", x"c1", x"b9", x"b5", x"ae", x"a8", x"a7", x"a7", x"a9", x"aa", x"ad", x"b0", 
        x"af", x"b4", x"d1", x"bb", x"9d", x"9a", x"9b", x"9b", x"9a", x"99", x"96", x"91", x"90", x"91", x"8f", 
        x"8b", x"86", x"83", x"85", x"83", x"80", x"7f", x"7f", x"7f", x"84", x"82", x"85", x"85", x"82", x"af", 
        x"cf", x"7c", x"71", x"71", x"74", x"73", x"6f", x"6e", x"69", x"66", x"64", x"68", x"69", x"6f", x"75", 
        x"76", x"75", x"73", x"6d", x"68", x"68", x"68", x"67", x"65", x"6a", x"a8", x"d1", x"8e", x"7c", x"81", 
        x"7c", x"7a", x"77", x"75", x"74", x"75", x"7c", x"80", x"7a", x"7c", x"7b", x"78", x"79", x"79", x"78", 
        x"7b", x"81", x"85", x"79", x"9a", x"d5", x"a4", x"80", x"82", x"89", x"8d", x"8f", x"8e", x"8a", x"85", 
        x"82", x"86", x"8e", x"90", x"94", x"96", x"90", x"8e", x"89", x"81", x"83", x"8c", x"bf", x"f1", x"f1", 
        x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f1", x"f0", x"ee", 
        x"ee", x"f0", x"ea", x"dd", x"c8", x"b9", x"bd", x"c1", x"c1", x"bd", x"b8", x"b5", x"b2", x"b1", x"b2", 
        x"b1", x"b0", x"b4", x"b9", x"bc", x"be", x"c0", x"94", x"3a", x"14", x"2f", x"4e", x"50", x"55", x"53", 
        x"4f", x"4c", x"48", x"48", x"4a", x"4c", x"4b", x"47", x"46", x"48", x"42", x"4b", x"60", x"6d", x"7c", 
        x"79", x"77", x"76", x"73", x"72", x"6f", x"6e", x"6e", x"6c", x"6a", x"68", x"6d", x"5d", x"29", x"2e", 
        x"4c", x"3d", x"3b", x"39", x"38", x"36", x"32", x"34", x"33", x"24", x"1c", x"1b", x"17", x"17", x"25", 
        x"32", x"19", x"05", x"07", x"14", x"16", x"14", x"16", x"19", x"15", x"12", x"12", x"17", x"1a", x"18", 
        x"19", x"34", x"3f", x"16", x"0f", x"11", x"10", x"0f", x"0d", x"0d", x"0d", x"0c", x"09", x"05", x"06", 
        x"05", x"0b", x"1a", x"0f", x"06", x"06", x"09", x"0a", x"0a", x"12", x"14", x"0d", x"08", x"06", x"05", 
        x"07", x"06", x"18", x"1c", x"13", x"12", x"15", x"23", x"53", x"8f", x"90", x"8c", x"96", x"93", x"90", 
        x"90", x"91", x"8d", x"7c", x"43", x"27", x"1e", x"0a", x"03", x"04", x"05", x"06", x"0a", x"3d", x"51", 
        x"4b", x"47", x"4b", x"57", x"54", x"51", x"52", x"4e", x"28", x"25", x"24", x"20", x"1e", x"19", x"15", 
        x"76", x"3d", x"3c", x"37", x"6b", x"8e", x"36", x"30", x"3a", x"49", x"2a", x"46", x"85", x"7f", x"4c", 
        x"40", x"3b", x"44", x"67", x"8f", x"95", x"83", x"78", x"76", x"71", x"80", x"ab", x"b3", x"b2", x"b4", 
        x"ae", x"a6", x"9e", x"ad", x"c3", x"c0", x"a6", x"a3", x"a2", x"9f", x"9e", x"9c", x"9c", x"98", x"98", 
        x"99", x"9a", x"99", x"99", x"99", x"99", x"9c", x"9c", x"9c", x"9e", x"a7", x"b4", x"b6", x"a3", x"98", 
        x"90", x"94", x"9f", x"b8", x"ba", x"a6", x"9d", x"9c", x"9d", x"a1", x"a4", x"a5", x"ab", x"ac", x"ab", 
        x"a8", x"a5", x"a4", x"a4", x"a4", x"a4", x"a8", x"af", x"b6", x"b9", x"bc", x"be", x"be", x"bd", x"bc", 
        x"bc", x"bc", x"bd", x"be", x"bf", x"c0", x"c1", x"c3", x"c7", x"cc", x"cf", x"d0", x"d0", x"d0", x"d0", 
        x"d0", x"cf", x"cd", x"ca", x"cf", x"d3", x"d3", x"d0", x"d5", x"dd", x"dd", x"d8", x"da", x"d9", x"e0", 
        x"ea", x"e0", x"dc", x"dd", x"dd", x"dc", x"dd", x"de", x"de", x"de", x"e1", x"e4", x"e2", x"e7", x"eb", 
        x"e9", x"e8", x"e6", x"e9", x"ea", x"e7", x"ea", x"eb", x"eb", x"e9", x"ea", x"eb", x"e9", x"e6", x"ea", 
        x"ec", x"e6", x"e6", x"eb", x"ee", x"eb", x"ec", x"ee", x"ea", x"ec", x"ec", x"ec", x"ec", x"ee", x"ed", 
        x"ec", x"ed", x"ec", x"e9", x"ea", x"ee", x"ef", x"ea", x"ed", x"ef", x"ef", x"ed", x"ed", x"ef", x"ed", 
        x"ee", x"ed", x"ed", x"ee", x"ef", x"f1", x"f2", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", 
        x"f1", x"f3", x"f2", x"f1", x"ef", x"ef", x"f3", x"f1", x"ed", x"ef", x"f2", x"f0", x"ef", x"f1", x"ed", 
        x"ef", x"f1", x"f0", x"ef", x"e0", x"e4", x"ef", x"ed", x"f2", x"f3", x"ef", x"ee", x"f0", x"ef", x"ee", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"ee", 
        x"ec", x"ee", x"f0", x"ef", x"ee", x"ef", x"ef", x"ee", x"ef", x"f0", x"ee", x"f0", x"f0", x"ef", x"f0", 
        x"f0", x"ed", x"ec", x"ee", x"ef", x"ee", x"f0", x"ef", x"ec", x"f1", x"f1", x"ef", x"ef", x"f0", x"f1", 
        x"f0", x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", 
        x"f0", x"f2", x"f0", x"ee", x"f0", x"f1", x"f2", x"f1", x"f0", x"ef", x"f2", x"f1", x"ee", x"f0", x"f4", 
        x"f3", x"f0", x"f0", x"f1", x"f2", x"f1", x"ee", x"f1", x"f3", x"f1", x"f0", x"f1", x"f2", x"f0", x"f0", 
        x"f2", x"f0", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f0", x"f0", x"f3", x"f3", x"f3", x"f1", x"f0", 
        x"f1", x"f3", x"f2", x"f1", x"f0", x"f0", x"f1", x"f2", x"f3", x"f1", x"f0", x"f0", x"ef", x"f0", x"f3", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", x"f0", 
        x"f0", x"f0", x"f0", x"f2", x"f3", x"f4", x"f2", x"f1", x"f3", x"f2", x"f2", x"f0", x"ef", x"f0", x"ec", 
        x"e7", x"f0", x"f2", x"f3", x"f2", x"f2", x"f3", x"f3", x"f0", x"ef", x"f2", x"f3", x"f1", x"ef", x"f1", 
        x"f2", x"f3", x"f5", x"f5", x"f3", x"f3", x"f4", x"f5", x"f5", x"f5", x"f5", x"f6", x"f5", x"f5", x"f5", 
        x"f3", x"f2", x"f5", x"f5", x"f4", x"f5", x"f5", x"f3", x"f2", x"f0", x"ec", x"ec", x"f0", x"ef", x"f0", 
        x"f2", x"f2", x"ef", x"ec", x"e7", x"e4", x"e6", x"e4", x"e2", x"e3", x"e3", x"e4", x"e5", x"e6", x"e3", 
        x"e0", x"dc", x"e3", x"e0", x"d6", x"d5", x"d6", x"db", x"db", x"dc", x"dd", x"dc", x"dc", x"dd", x"dc", 
        x"d3", x"ca", x"c7", x"c9", x"c7", x"c6", x"c8", x"c8", x"c7", x"c9", x"c9", x"cd", x"cb", x"c3", x"cd", 
        x"d7", x"a5", x"9b", x"9a", x"9c", x"9a", x"97", x"96", x"93", x"8b", x"87", x"87", x"86", x"8a", x"8f", 
        x"8f", x"91", x"92", x"92", x"94", x"94", x"91", x"8d", x"8a", x"8c", x"b3", x"d2", x"9e", x"8b", x"87", 
        x"85", x"82", x"7f", x"81", x"85", x"85", x"82", x"81", x"81", x"80", x"7b", x"77", x"7a", x"7e", x"81", 
        x"80", x"7e", x"7a", x"73", x"93", x"d1", x"aa", x"88", x"87", x"88", x"88", x"8c", x"94", x"98", x"93", 
        x"8c", x"86", x"83", x"82", x"85", x"8a", x"8d", x"96", x"97", x"8f", x"88", x"87", x"b9", x"f1", x"f1", 
        x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f3", x"f2", x"f3", x"f2", 
        x"ef", x"ee", x"eb", x"e0", x"c8", x"b4", x"b4", x"b5", x"b5", x"b4", x"b5", x"b9", x"be", x"c2", x"c2", 
        x"bd", x"b8", x"b7", x"b5", x"b4", x"b4", x"b7", x"b6", x"5c", x"2c", x"3f", x"4d", x"4e", x"4f", x"49", 
        x"47", x"49", x"47", x"47", x"48", x"48", x"46", x"45", x"47", x"49", x"43", x"48", x"5d", x"69", x"7a", 
        x"78", x"76", x"75", x"73", x"71", x"6e", x"6f", x"6f", x"6f", x"6d", x"6b", x"71", x"64", x"2b", x"28", 
        x"49", x"3c", x"39", x"35", x"37", x"38", x"36", x"38", x"36", x"25", x"18", x"15", x"15", x"18", x"20", 
        x"33", x"23", x"0c", x"0c", x"19", x"1c", x"1b", x"1e", x"20", x"1d", x"1c", x"1d", x"21", x"1e", x"17", 
        x"19", x"33", x"3e", x"16", x"10", x"12", x"0e", x"0d", x"0c", x"0d", x"0c", x"0b", x"08", x"06", x"05", 
        x"05", x"0c", x"1a", x"12", x"0a", x"0c", x"0f", x"10", x"12", x"16", x"17", x"11", x"0b", x"08", x"07", 
        x"08", x"08", x"19", x"1c", x"0f", x"0f", x"10", x"21", x"51", x"92", x"9f", x"a9", x"bb", x"b9", x"a7", 
        x"8e", x"8b", x"8c", x"7f", x"48", x"28", x"1c", x"0b", x"04", x"04", x"06", x"07", x"0a", x"3c", x"4f", 
        x"48", x"47", x"4c", x"59", x"58", x"56", x"58", x"50", x"27", x"23", x"22", x"1a", x"15", x"1b", x"15", 
        x"59", x"3d", x"33", x"2a", x"5a", x"62", x"32", x"2e", x"57", x"5d", x"3f", x"55", x"7c", x"40", x"2a", 
        x"2d", x"28", x"29", x"36", x"40", x"81", x"93", x"99", x"a0", x"9d", x"ad", x"dc", x"e1", x"de", x"e1", 
        x"e2", x"de", x"d4", x"d8", x"da", x"d8", x"da", x"d6", x"d9", x"da", x"da", x"da", x"dc", x"d9", x"d7", 
        x"d8", x"d8", x"d7", x"d6", x"d6", x"d8", x"db", x"da", x"d9", x"d9", x"db", x"de", x"dc", x"cf", x"cd", 
        x"ca", x"d0", x"d3", x"dd", x"dc", x"d6", x"d1", x"d1", x"d0", x"ce", x"cc", x"c9", x"cb", x"ca", x"c5", 
        x"c2", x"bf", x"bd", x"be", x"bd", x"bc", x"ba", x"ba", x"bc", x"bb", x"ba", x"bb", x"bc", x"b7", x"b8", 
        x"b5", x"b3", x"b3", x"b4", x"b4", x"b1", x"b4", x"b2", x"b2", x"b6", x"b7", x"b5", x"b4", x"b1", x"ae", 
        x"a9", x"a5", x"a2", x"a2", x"a0", x"9f", x"9d", x"a5", x"bc", x"cc", x"b5", x"a5", x"a9", x"ad", x"bd", 
        x"cd", x"c2", x"a7", x"a2", x"a4", x"a2", x"a3", x"a4", x"a6", x"a8", x"a7", x"ac", x"af", x"b3", x"bd", 
        x"ba", x"b9", x"b8", x"b8", x"b7", x"b3", x"b5", x"b7", x"b7", x"b7", x"b8", x"b8", x"ba", x"ba", x"ba", 
        x"be", x"c0", x"c3", x"c6", x"c4", x"c2", x"c5", x"c2", x"c3", x"c2", x"c0", x"c1", x"c3", x"c7", x"c6", 
        x"c9", x"d0", x"d5", x"d5", x"d2", x"d8", x"e4", x"e9", x"d9", x"d0", x"d1", x"d2", x"e1", x"e5", x"d4", 
        x"d0", x"cf", x"d0", x"d2", x"d4", x"d8", x"dc", x"dd", x"de", x"e0", x"de", x"de", x"df", x"dc", x"da", 
        x"dd", x"df", x"e0", x"df", x"e2", x"e1", x"e0", x"e0", x"de", x"df", x"e2", x"e1", x"e2", x"e4", x"e2", 
        x"e6", x"e7", x"e5", x"e7", x"dd", x"df", x"e7", x"e4", x"e5", x"e4", x"e2", x"e5", x"ea", x"eb", x"ec", 
        x"ea", x"e9", x"eb", x"f0", x"ec", x"eb", x"eb", x"ea", x"eb", x"ec", x"eb", x"ed", x"ef", x"f0", x"ef", 
        x"ed", x"ef", x"f0", x"f0", x"ee", x"f0", x"f1", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"ef", x"f1", 
        x"f0", x"ef", x"f1", x"f3", x"f3", x"ef", x"f0", x"f3", x"f1", x"f2", x"f2", x"f2", x"f0", x"f1", x"f4", 
        x"f4", x"f2", x"f2", x"f1", x"f0", x"f0", x"f0", x"f2", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", 
        x"f0", x"f1", x"f0", x"f1", x"f0", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f1", x"f2", x"f1", 
        x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"f0", x"f3", x"ee", x"ee", x"ed", x"f0", x"f1", x"f0", x"ed", 
        x"f1", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"ef", x"f0", x"f1", x"f2", x"f0", x"ef", x"f0", 
        x"f1", x"f3", x"f3", x"f3", x"f2", x"f0", x"f0", x"f1", x"f2", x"f0", x"f0", x"f3", x"f3", x"f2", x"f1", 
        x"f1", x"f1", x"f1", x"f0", x"f2", x"f2", x"f2", x"f1", x"f3", x"f3", x"f3", x"f4", x"f3", x"f1", x"f2", 
        x"f2", x"f3", x"f1", x"f2", x"f2", x"f3", x"f3", x"f2", x"f2", x"f2", x"f2", x"f1", x"f1", x"f3", x"ed", 
        x"e7", x"f1", x"ef", x"f0", x"f3", x"f1", x"f2", x"f3", x"f4", x"f2", x"f4", x"f2", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f2", x"f1", x"f2", x"f2", x"f2", x"f3", x"f3", x"f2", x"f1", x"f0", x"f1", x"f3", 
        x"f1", x"f1", x"f3", x"f1", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f2", x"f2", x"f2", x"f3", x"f4", 
        x"f3", x"f2", x"f2", x"f2", x"f2", x"f3", x"f4", x"f2", x"f1", x"f3", x"f4", x"f3", x"f3", x"f3", x"f2", 
        x"f3", x"f0", x"ef", x"f2", x"f0", x"f2", x"f1", x"f6", x"f7", x"f7", x"f6", x"f5", x"f4", x"f4", x"f3", 
        x"f1", x"f1", x"f3", x"f3", x"f1", x"f1", x"f4", x"f1", x"ef", x"f0", x"f1", x"ee", x"ea", x"eb", x"e5", 
        x"e8", x"e3", x"e0", x"e0", x"e2", x"e3", x"e0", x"e0", x"df", x"e0", x"dd", x"d8", x"d4", x"d4", x"d5", 
        x"d5", x"d8", x"d7", x"d8", x"d9", x"da", x"db", x"da", x"dc", x"da", x"e0", x"ea", x"da", x"d5", x"ce", 
        x"d1", x"cd", x"cf", x"d6", x"d9", x"d1", x"c9", x"c6", x"c1", x"bf", x"bb", x"b9", x"bf", x"c8", x"cc", 
        x"c6", x"c0", x"b7", x"ad", x"ba", x"da", x"c0", x"b4", x"b6", x"b1", x"a7", x"a0", x"9f", x"a0", x"a2", 
        x"a4", x"a5", x"a5", x"a3", x"9c", x"98", x"97", x"9c", x"9e", x"9b", x"9a", x"97", x"bc", x"ed", x"f0", 
        x"ee", x"ed", x"ee", x"ee", x"ef", x"f1", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f2", x"f1", 
        x"ef", x"ef", x"ec", x"e1", x"ce", x"c1", x"c3", x"c5", x"c3", x"be", x"ba", x"b8", x"b9", x"ba", x"bb", 
        x"b9", x"bb", x"bf", x"c0", x"bf", x"bf", x"bf", x"cd", x"73", x"41", x"53", x"49", x"4e", x"51", x"4e", 
        x"4e", x"4f", x"4d", x"4c", x"4d", x"4e", x"4b", x"49", x"4b", x"49", x"41", x"47", x"5f", x"6a", x"7a", 
        x"78", x"77", x"78", x"78", x"76", x"74", x"73", x"73", x"72", x"6e", x"6d", x"71", x"66", x"2b", x"24", 
        x"47", x"3d", x"3c", x"3c", x"3f", x"3e", x"37", x"35", x"32", x"20", x"12", x"11", x"14", x"1a", x"21", 
        x"35", x"2d", x"12", x"10", x"1d", x"20", x"1e", x"20", x"21", x"1f", x"1e", x"1d", x"1c", x"15", x"12", 
        x"18", x"32", x"41", x"19", x"12", x"12", x"0e", x"0f", x"0d", x"0d", x"0a", x"09", x"08", x"06", x"04", 
        x"02", x"09", x"18", x"11", x"08", x"0b", x"12", x"0f", x"0e", x"10", x"11", x"0d", x"08", x"06", x"07", 
        x"06", x"07", x"18", x"1d", x"0e", x"11", x"11", x"20", x"50", x"9c", x"ac", x"b9", x"d2", x"d9", x"d5", 
        x"bc", x"9b", x"80", x"7d", x"53", x"32", x"23", x"0d", x"06", x"07", x"08", x"06", x"09", x"37", x"4c", 
        x"48", x"4a", x"4c", x"58", x"59", x"58", x"5a", x"54", x"27", x"22", x"25", x"1d", x"14", x"18", x"15", 
        x"51", x"49", x"58", x"2f", x"5a", x"75", x"37", x"42", x"88", x"6c", x"43", x"33", x"4e", x"41", x"31", 
        x"20", x"28", x"27", x"2b", x"4e", x"a7", x"a8", x"a4", x"a4", x"9b", x"ab", x"de", x"de", x"de", x"de", 
        x"de", x"da", x"d5", x"d5", x"d0", x"d1", x"b8", x"a4", x"d2", x"d7", x"d8", x"da", x"da", x"db", x"d6", 
        x"d9", x"d9", x"d7", x"d7", x"d8", x"d9", x"de", x"de", x"db", x"da", x"d5", x"d0", x"d0", x"d9", x"db", 
        x"d4", x"e0", x"de", x"d4", x"d1", x"db", x"df", x"df", x"dd", x"dd", x"de", x"e0", x"e3", x"e4", x"e1", 
        x"e3", x"e5", x"e2", x"e2", x"e2", x"d6", x"de", x"e4", x"e3", x"e5", x"e6", x"e6", x"e5", x"e1", x"e8", 
        x"ea", x"e8", x"e9", x"e9", x"e8", x"e7", x"eb", x"ea", x"e8", x"e7", x"e9", x"e8", x"e7", x"e6", x"e5", 
        x"e4", x"e4", x"e5", x"e7", x"e2", x"e1", x"e1", x"df", x"e1", x"e3", x"de", x"dd", x"dd", x"db", x"de", 
        x"e0", x"df", x"d4", x"d6", x"d6", x"cf", x"d0", x"ce", x"ca", x"cd", x"cd", x"cb", x"cd", x"c7", x"ca", 
        x"c4", x"c3", x"c2", x"c1", x"c1", x"bf", x"bc", x"bc", x"bb", x"bc", x"bc", x"ba", x"b9", x"bb", x"b9", 
        x"bb", x"ba", x"b9", x"bb", x"b4", x"b4", x"b6", x"b5", x"b2", x"ad", x"ab", x"ab", x"ad", x"ae", x"af", 
        x"af", x"b2", x"b4", x"b7", x"b2", x"b4", x"cf", x"e0", x"b5", x"a3", x"a8", x"ab", x"cb", x"d1", x"ae", 
        x"a3", x"a4", x"a5", x"a8", x"ac", x"b0", x"b3", x"b8", x"b8", x"b8", x"b4", x"b4", x"b2", x"ae", x"ad", 
        x"b0", x"b2", x"b5", x"b5", x"bb", x"ba", x"b9", x"b3", x"af", x"ad", x"af", x"b5", x"b6", x"b8", x"bc", 
        x"be", x"bf", x"bd", x"c2", x"cd", x"c8", x"bd", x"bb", x"b9", x"b7", x"b4", x"bc", x"d2", x"e2", x"d1", 
        x"c8", x"ca", x"d5", x"e8", x"da", x"cd", x"cc", x"c9", x"ca", x"cb", x"c9", x"cd", x"d0", x"d4", x"d5", 
        x"d8", x"d7", x"d6", x"d7", x"d6", x"d6", x"d9", x"d6", x"d6", x"d7", x"d9", x"d9", x"db", x"dc", x"e1", 
        x"e3", x"e3", x"e4", x"e2", x"e2", x"e0", x"e3", x"e4", x"e3", x"e5", x"e3", x"e4", x"e0", x"e5", x"e6", 
        x"e6", x"e4", x"eb", x"ed", x"e7", x"e8", x"e9", x"f0", x"eb", x"e7", x"e9", x"e9", x"ea", x"ed", x"ef", 
        x"f0", x"f0", x"ef", x"f1", x"ef", x"f1", x"ee", x"ef", x"ef", x"f1", x"ee", x"f1", x"f3", x"f3", x"f3", 
        x"f1", x"f1", x"f1", x"f2", x"f3", x"f4", x"f2", x"f4", x"f2", x"f2", x"f1", x"f4", x"f3", x"f4", x"ef", 
        x"f2", x"f4", x"f3", x"ef", x"f3", x"f4", x"f2", x"f1", x"f2", x"f3", x"f4", x"f4", x"f2", x"f2", x"f3", 
        x"f3", x"f3", x"f3", x"f3", x"f3", x"f3", x"f2", x"f3", x"f3", x"f0", x"ef", x"f0", x"f4", x"ef", x"f1", 
        x"f0", x"f0", x"f1", x"f2", x"f4", x"f3", x"f0", x"f1", x"f2", x"f1", x"f4", x"f4", x"f2", x"ef", x"f1", 
        x"f1", x"f4", x"f1", x"f2", x"f2", x"f2", x"f4", x"f1", x"f0", x"f2", x"f2", x"f1", x"f0", x"f4", x"f1", 
        x"e1", x"f0", x"f1", x"ef", x"f5", x"f3", x"f2", x"f2", x"f3", x"ef", x"f1", x"ef", x"f0", x"f2", x"f3", 
        x"f5", x"f2", x"f1", x"f2", x"f1", x"f3", x"f2", x"f1", x"f4", x"f4", x"f3", x"f2", x"f3", x"f0", x"f1", 
        x"f2", x"f3", x"f4", x"f2", x"f2", x"f3", x"f4", x"f4", x"f2", x"f2", x"f2", x"f2", x"f1", x"f3", x"f3", 
        x"f1", x"f2", x"f3", x"f3", x"f4", x"f5", x"f5", x"f3", x"f3", x"f1", x"f2", x"f1", x"ef", x"f4", x"f4", 
        x"f5", x"f1", x"f2", x"f2", x"f1", x"f0", x"f2", x"f4", x"f7", x"f9", x"f9", x"f6", x"f3", x"f1", x"f2", 
        x"f3", x"f3", x"f4", x"f3", x"f2", x"f4", x"f2", x"f1", x"f2", x"f1", x"f0", x"f2", x"f2", x"f2", x"f2", 
        x"f1", x"f1", x"f3", x"f5", x"f4", x"f7", x"f4", x"f5", x"f4", x"f6", x"f5", x"f4", x"f4", x"f5", x"f5", 
        x"f3", x"f4", x"f4", x"f4", x"f3", x"f6", x"f8", x"f9", x"f8", x"f6", x"f4", x"ef", x"f4", x"fa", x"f8", 
        x"f9", x"f8", x"f7", x"f5", x"f3", x"f1", x"f0", x"f0", x"f0", x"f0", x"f2", x"f3", x"f4", x"f5", x"f5", 
        x"f1", x"ed", x"e9", x"e5", x"e5", x"e7", x"ea", x"f0", x"f0", x"ec", x"e7", x"e4", x"e1", x"df", x"e1", 
        x"e4", x"ea", x"ef", x"f0", x"e9", x"e0", x"d9", x"d4", x"cd", x"cb", x"cd", x"cd", x"d7", x"ee", x"f3", 
        x"f0", x"f0", x"f1", x"f0", x"f2", x"f4", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"ef", 
        x"f5", x"f2", x"ee", x"dd", x"d5", x"c7", x"c2", x"c1", x"c0", x"bf", x"c0", x"c3", x"c8", x"cc", x"cd", 
        x"cd", x"cc", x"c9", x"c8", x"c4", x"be", x"be", x"c9", x"76", x"3c", x"5e", x"57", x"58", x"57", x"58", 
        x"54", x"4e", x"4b", x"47", x"47", x"4a", x"49", x"45", x"45", x"45", x"41", x"48", x"66", x"71", x"7c", 
        x"78", x"77", x"77", x"73", x"73", x"74", x"72", x"71", x"71", x"6f", x"6d", x"6f", x"69", x"2f", x"22", 
        x"42", x"3c", x"37", x"36", x"3a", x"37", x"2d", x"2b", x"2f", x"1f", x"11", x"10", x"11", x"19", x"24", 
        x"36", x"2a", x"0d", x"0b", x"15", x"19", x"15", x"18", x"19", x"17", x"16", x"12", x"10", x"0c", x"14", 
        x"18", x"30", x"47", x"1b", x"11", x"10", x"0e", x"13", x"10", x"0d", x"0c", x"08", x"07", x"07", x"04", 
        x"02", x"08", x"16", x"11", x"05", x"08", x"0f", x"0b", x"0a", x"0b", x"0a", x"0d", x"08", x"07", x"09", 
        x"08", x"0a", x"19", x"21", x"11", x"14", x"13", x"23", x"54", x"a3", x"ad", x"b5", x"ce", x"d6", x"de", 
        x"e7", x"cf", x"92", x"76", x"51", x"2d", x"20", x"0a", x"03", x"05", x"02", x"02", x"07", x"30", x"4d", 
        x"48", x"4a", x"4a", x"56", x"54", x"4e", x"53", x"53", x"25", x"1a", x"1c", x"19", x"15", x"14", x"16", 
        x"4f", x"3c", x"5d", x"45", x"73", x"93", x"4b", x"63", x"60", x"2c", x"31", x"32", x"31", x"30", x"2e", 
        x"32", x"28", x"32", x"3c", x"53", x"a6", x"a5", x"a6", x"a6", x"a0", x"b0", x"e1", x"e0", x"e1", x"e0", 
        x"df", x"db", x"d4", x"d3", x"d9", x"cf", x"80", x"95", x"e0", x"dd", x"da", x"d9", x"dd", x"df", x"d7", 
        x"dc", x"db", x"dd", x"dc", x"d9", x"dc", x"dc", x"dd", x"db", x"dd", x"d8", x"dd", x"dd", x"e0", x"dd", 
        x"d4", x"df", x"df", x"dd", x"dc", x"d8", x"da", x"db", x"da", x"db", x"da", x"dc", x"dd", x"df", x"db", 
        x"db", x"de", x"dc", x"dc", x"d6", x"94", x"be", x"e0", x"db", x"e0", x"df", x"e0", x"da", x"dc", x"df", 
        x"e2", x"e3", x"e2", x"de", x"db", x"e3", x"de", x"e1", x"e0", x"dc", x"e1", x"e0", x"df", x"df", x"df", 
        x"de", x"df", x"df", x"df", x"df", x"e1", x"e0", x"da", x"d5", x"d5", x"dc", x"e0", x"dd", x"db", x"d7", 
        x"d5", x"d5", x"db", x"dd", x"dd", x"dc", x"dd", x"df", x"de", x"df", x"dd", x"e2", x"e1", x"e3", x"e0", 
        x"dd", x"de", x"de", x"de", x"e2", x"df", x"e4", x"e3", x"e0", x"df", x"de", x"df", x"e3", x"e4", x"e1", 
        x"df", x"e0", x"df", x"e1", x"e1", x"e0", x"e3", x"ce", x"dd", x"e1", x"e3", x"e2", x"e2", x"e1", x"e1", 
        x"e0", x"e1", x"e0", x"dd", x"e3", x"de", x"d9", x"d9", x"dc", x"da", x"dd", x"de", x"dc", x"da", x"de", 
        x"db", x"dd", x"df", x"e0", x"e1", x"e3", x"de", x"dc", x"dd", x"df", x"df", x"dd", x"d9", x"dd", x"d9", 
        x"d9", x"da", x"d8", x"d9", x"d8", x"db", x"dd", x"dc", x"d3", x"d5", x"d7", x"d7", x"d8", x"d7", x"d5", 
        x"d4", x"d5", x"d6", x"d5", x"dc", x"d8", x"d3", x"d2", x"d1", x"d2", x"cc", x"ce", x"d8", x"e3", x"d8", 
        x"d0", x"cd", x"d5", x"e3", x"da", x"ce", x"d0", x"cc", x"cb", x"c7", x"c4", x"c3", x"c2", x"c4", x"c5", 
        x"c8", x"c9", x"c5", x"c5", x"c6", x"c2", x"c3", x"c5", x"c2", x"c1", x"c2", x"be", x"c2", x"c3", x"c4", 
        x"c5", x"c5", x"c6", x"c1", x"c0", x"be", x"c0", x"c2", x"c0", x"c5", x"c6", x"c4", x"c4", x"c2", x"c0", 
        x"c4", x"c1", x"dd", x"e0", x"c0", x"bc", x"ca", x"df", x"de", x"c6", x"c4", x"c2", x"c5", x"c7", x"c8", 
        x"c8", x"c8", x"cb", x"c8", x"c8", x"c8", x"c4", x"c8", x"c4", x"c1", x"c0", x"c2", x"c8", x"cd", x"cc", 
        x"ce", x"d4", x"d3", x"d3", x"d2", x"d0", x"cf", x"d0", x"cf", x"ce", x"cc", x"ce", x"cd", x"d3", x"e7", 
        x"df", x"d3", x"d6", x"e3", x"e4", x"d8", x"d8", x"d6", x"d6", x"d8", x"db", x"db", x"dd", x"e1", x"e6", 
        x"e7", x"e6", x"e7", x"e7", x"e7", x"e8", x"e8", x"e9", x"e9", x"ea", x"ed", x"e9", x"ec", x"e7", x"ee", 
        x"ec", x"ee", x"ef", x"f1", x"ef", x"ee", x"f3", x"f4", x"f5", x"ef", x"f2", x"f5", x"f3", x"f1", x"f4", 
        x"f3", x"f1", x"f2", x"f4", x"f6", x"f6", x"f4", x"f4", x"f4", x"f5", x"f7", x"f7", x"f6", x"f6", x"f6", 
        x"e4", x"ef", x"f3", x"f4", x"f5", x"f3", x"f4", x"f4", x"f3", x"f4", x"f6", x"f4", x"f4", x"f5", x"f5", 
        x"f3", x"f6", x"f4", x"f4", x"f6", x"f5", x"f2", x"f3", x"f3", x"f3", x"f3", x"f5", x"f5", x"f2", x"f3", 
        x"f4", x"f3", x"f4", x"f4", x"f3", x"f4", x"f4", x"f4", x"f3", x"f3", x"f3", x"f3", x"f4", x"f4", x"f2", 
        x"f2", x"f4", x"f4", x"f3", x"f4", x"f8", x"f6", x"f2", x"f3", x"f3", x"f0", x"ef", x"f0", x"f4", x"f2", 
        x"f2", x"f1", x"f2", x"f2", x"f1", x"f1", x"f3", x"f6", x"f8", x"f9", x"f8", x"f6", x"f3", x"f2", x"f3", 
        x"f4", x"f4", x"f4", x"f1", x"f0", x"f3", x"f0", x"f1", x"f4", x"f2", x"f3", x"f4", x"f3", x"f2", x"f2", 
        x"f2", x"f0", x"f2", x"f5", x"f1", x"f0", x"f1", x"f4", x"f2", x"f4", x"f4", x"f3", x"f4", x"f4", x"f3", 
        x"f3", x"ef", x"f1", x"f1", x"f2", x"f6", x"f4", x"f2", x"f4", x"f4", x"f3", x"ee", x"f1", x"f9", x"f7", 
        x"f4", x"f4", x"f3", x"f1", x"f1", x"f2", x"f3", x"f3", x"f0", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", 
        x"f1", x"ef", x"f0", x"f2", x"f1", x"f1", x"f1", x"f1", x"f1", x"f2", x"f3", x"f3", x"f3", x"f2", x"f1", 
        x"f1", x"f0", x"f2", x"f2", x"f2", x"f0", x"f1", x"f0", x"ed", x"f1", x"ee", x"ed", x"f1", x"f0", x"f0", 
        x"f0", x"f1", x"f3", x"f0", x"ee", x"ef", x"ee", x"ee", x"ef", x"f0", x"f0", x"f1", x"f1", x"f2", x"f0", 
        x"f0", x"ef", x"f1", x"eb", x"eb", x"e2", x"df", x"df", x"df", x"e0", x"e2", x"e6", x"e8", x"ea", x"ea", 
        x"e8", x"e2", x"de", x"d9", x"d8", x"d8", x"da", x"e0", x"89", x"39", x"5d", x"6e", x"6b", x"67", x"68", 
        x"6a", x"6b", x"69", x"66", x"64", x"64", x"63", x"61", x"5f", x"5d", x"5c", x"59", x"68", x"73", x"79", 
        x"76", x"72", x"6e", x"6c", x"6c", x"6e", x"6c", x"6b", x"6a", x"68", x"67", x"66", x"64", x"30", x"21", 
        x"48", x"4d", x"45", x"43", x"42", x"40", x"38", x"36", x"36", x"27", x"19", x"1a", x"1b", x"20", x"24", 
        x"3a", x"3d", x"2b", x"28", x"2e", x"2f", x"2a", x"29", x"23", x"24", x"23", x"1b", x"1a", x"20", x"22", 
        x"18", x"2f", x"47", x"1b", x"0a", x"0c", x"0b", x"0d", x"0a", x"08", x"08", x"06", x"04", x"06", x"07", 
        x"05", x"07", x"14", x"11", x"0a", x"09", x"05", x"09", x"0a", x"0b", x"09", x"09", x"07", x"06", x"06", 
        x"05", x"06", x"10", x"16", x"08", x"09", x"09", x"1f", x"4f", x"9d", x"aa", x"b4", x"ce", x"d6", x"d9", 
        x"e1", x"e7", x"d3", x"93", x"58", x"33", x"29", x"0f", x"05", x"04", x"02", x"04", x"0a", x"30", x"4e", 
        x"46", x"47", x"47", x"54", x"54", x"4d", x"4f", x"50", x"25", x"16", x"17", x"26", x"30", x"1f", x"17", 
        x"4e", x"38", x"42", x"46", x"88", x"88", x"42", x"56", x"45", x"2e", x"3e", x"3e", x"32", x"36", x"2d", 
        x"33", x"33", x"4a", x"4a", x"56", x"a6", x"a6", x"a4", x"a5", x"a0", x"b1", x"e0", x"e0", x"e0", x"e1", 
        x"e2", x"d8", x"d2", x"d8", x"d8", x"c7", x"9d", x"ca", x"e1", x"db", x"d6", x"d9", x"dd", x"da", x"db", 
        x"dc", x"d8", x"db", x"d8", x"d8", x"dd", x"e0", x"da", x"db", x"df", x"db", x"db", x"dc", x"de", x"d9", 
        x"d0", x"dc", x"dc", x"dd", x"de", x"db", x"de", x"df", x"df", x"e0", x"dd", x"dd", x"dc", x"df", x"dc", 
        x"db", x"dd", x"dc", x"dd", x"d7", x"7f", x"b5", x"e2", x"dc", x"de", x"dd", x"df", x"e0", x"de", x"e1", 
        x"df", x"e2", x"e5", x"e3", x"e2", x"db", x"df", x"e2", x"df", x"df", x"e1", x"df", x"df", x"df", x"df", 
        x"df", x"e0", x"e0", x"de", x"de", x"df", x"e0", x"df", x"df", x"df", x"de", x"de", x"d8", x"db", x"db", 
        x"da", x"db", x"de", x"dc", x"dc", x"dc", x"db", x"e0", x"e0", x"df", x"dc", x"dd", x"dc", x"df", x"dc", 
        x"dd", x"dc", x"db", x"dc", x"dc", x"dc", x"dc", x"dd", x"dd", x"dc", x"dc", x"e1", x"c2", x"cd", x"dd", 
        x"dd", x"de", x"de", x"de", x"dc", x"dd", x"de", x"a7", x"d2", x"e0", x"df", x"de", x"de", x"dd", x"dd", 
        x"de", x"de", x"e1", x"dd", x"e0", x"df", x"d9", x"d5", x"de", x"dd", x"df", x"de", x"dc", x"d9", x"e3", 
        x"e2", x"e2", x"e4", x"e4", x"e1", x"e5", x"e6", x"e4", x"e4", x"e6", x"e7", x"e6", x"e0", x"e6", x"e6", 
        x"e5", x"e6", x"e5", x"e6", x"e5", x"e7", x"e8", x"e7", x"c5", x"cf", x"ec", x"e7", x"e8", x"e8", x"e6", 
        x"e8", x"e8", x"e9", x"e6", x"e5", x"e4", x"ea", x"ea", x"e8", x"eb", x"ea", x"e9", x"e1", x"df", x"e7", 
        x"ea", x"e2", x"de", x"e1", x"df", x"e3", x"e8", x"e6", x"e5", x"e6", x"e3", x"e3", x"e2", x"e2", x"e5", 
        x"e3", x"e0", x"e1", x"e2", x"e5", x"e1", x"e0", x"e1", x"e4", x"e0", x"e0", x"dd", x"dd", x"df", x"dc", 
        x"d9", x"d9", x"d9", x"d7", x"d6", x"d8", x"d8", x"d5", x"d7", x"d9", x"d5", x"d7", x"d7", x"d1", x"d7", 
        x"d1", x"d0", x"de", x"e0", x"cd", x"cb", x"d5", x"de", x"dc", x"d2", x"d0", x"cb", x"c9", x"c8", x"c9", 
        x"c9", x"c9", x"ca", x"c5", x"c8", x"c6", x"c2", x"c7", x"c1", x"bd", x"bb", x"bb", x"c3", x"c3", x"c1", 
        x"c5", x"c5", x"c6", x"c7", x"c3", x"c4", x"c6", x"c0", x"bd", x"bb", x"b6", x"b4", x"b2", x"bf", x"dc", 
        x"ce", x"b9", x"bf", x"d6", x"d4", x"c0", x"bf", x"bd", x"bb", x"bd", x"be", x"bd", x"bc", x"c1", x"c7", 
        x"c9", x"c9", x"c9", x"c9", x"ca", x"cb", x"cb", x"cd", x"ca", x"c7", x"ca", x"c8", x"c7", x"c0", x"c2", 
        x"c2", x"c9", x"cb", x"ce", x"ce", x"cd", x"d1", x"d3", x"d1", x"d5", x"e4", x"e1", x"d1", x"cc", x"e2", 
        x"e1", x"d5", x"d4", x"d9", x"dd", x"dd", x"dc", x"e0", x"e1", x"e1", x"de", x"db", x"da", x"da", x"dc", 
        x"e0", x"e1", x"e6", x"e1", x"de", x"dc", x"dc", x"d7", x"d5", x"da", x"d8", x"d7", x"db", x"e0", x"e0", 
        x"df", x"df", x"e3", x"ed", x"e8", x"e1", x"e6", x"eb", x"e2", x"e3", x"e6", x"e5", x"e6", x"e7", x"ec", 
        x"ed", x"ea", x"ee", x"ee", x"ed", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ef", x"f2", x"f3", x"f2", x"f3", x"f2", x"f3", x"f4", x"f3", x"f3", x"f1", x"f1", x"f2", x"f4", x"f2", 
        x"f2", x"f2", x"f4", x"f4", x"f3", x"f4", x"f5", x"f8", x"f8", x"f8", x"f7", x"f6", x"f4", x"f4", x"f5", 
        x"f5", x"f4", x"f5", x"f3", x"f2", x"f5", x"f5", x"f3", x"f4", x"f6", x"f3", x"f3", x"f2", x"f2", x"f3", 
        x"f4", x"f2", x"f2", x"f4", x"f3", x"f3", x"f4", x"f5", x"f4", x"f2", x"f3", x"f3", x"f4", x"f3", x"f4", 
        x"f5", x"f1", x"f2", x"f4", x"f4", x"f5", x"f5", x"f3", x"f4", x"f5", x"f5", x"f1", x"ef", x"f7", x"f9", 
        x"f5", x"f3", x"f2", x"f1", x"f1", x"f2", x"f4", x"f3", x"f1", x"f1", x"f1", x"f1", x"f2", x"f2", x"f2", 
        x"f0", x"f2", x"f1", x"f1", x"f3", x"f2", x"f2", x"ef", x"ee", x"f0", x"f1", x"f1", x"f0", x"ee", x"ef", 
        x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f3", x"f4", x"ef", x"f1", x"f2", x"f0", x"f1", x"ef", x"ef", 
        x"f0", x"f0", x"f2", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", 
        x"ec", x"ec", x"f0", x"ef", x"f1", x"f0", x"f0", x"f1", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"ee", x"ed", x"ed", x"ef", x"ec", x"ec", x"f2", x"a0", x"3f", x"63", x"88", x"86", x"86", x"87", 
        x"87", x"86", x"85", x"86", x"85", x"83", x"82", x"81", x"7e", x"7b", x"7b", x"75", x"76", x"79", x"7a", 
        x"77", x"76", x"73", x"74", x"74", x"74", x"71", x"6f", x"6e", x"6d", x"6b", x"6a", x"6a", x"37", x"21", 
        x"51", x"6f", x"6c", x"69", x"66", x"65", x"63", x"61", x"60", x"51", x"3d", x"39", x"39", x"35", x"28", 
        x"3b", x"54", x"4d", x"4c", x"55", x"5a", x"55", x"56", x"52", x"50", x"49", x"45", x"48", x"51", x"46", 
        x"21", x"2a", x"50", x"3f", x"34", x"34", x"30", x"30", x"2e", x"2a", x"27", x"27", x"1c", x"0d", x"0b", 
        x"0a", x"0e", x"22", x"29", x"23", x"22", x"23", x"21", x"23", x"25", x"23", x"24", x"23", x"23", x"27", 
        x"25", x"23", x"26", x"2b", x"25", x"25", x"25", x"2e", x"50", x"99", x"a8", x"b2", x"cb", x"d4", x"d8", 
        x"dd", x"e4", x"ec", x"bb", x"5d", x"36", x"25", x"0d", x"04", x"03", x"03", x"06", x"07", x"28", x"4c", 
        x"47", x"49", x"4a", x"55", x"54", x"4f", x"53", x"55", x"2e", x"19", x"18", x"31", x"42", x"27", x"16", 
        x"3c", x"3e", x"35", x"52", x"99", x"70", x"3e", x"4d", x"44", x"3c", x"42", x"4b", x"41", x"40", x"2c", 
        x"2f", x"3f", x"48", x"3f", x"5e", x"a6", x"a3", x"a1", x"a2", x"9e", x"b0", x"df", x"de", x"df", x"e0", 
        x"e0", x"dd", x"d8", x"d8", x"a9", x"7e", x"75", x"86", x"bc", x"dc", x"d8", x"d9", x"d8", x"d9", x"de", 
        x"dc", x"da", x"d6", x"da", x"de", x"c9", x"8f", x"7d", x"8f", x"c7", x"e6", x"dc", x"dc", x"dd", x"d7", 
        x"ce", x"dd", x"de", x"db", x"dc", x"e3", x"cc", x"9a", x"93", x"af", x"e0", x"df", x"db", x"dc", x"dd", 
        x"dd", x"de", x"de", x"dd", x"d9", x"89", x"b6", x"e2", x"dc", x"dd", x"de", x"e0", x"de", x"dc", x"e0", 
        x"e5", x"d5", x"b8", x"bc", x"dd", x"e8", x"e1", x"dc", x"df", x"e1", x"de", x"dd", x"dd", x"dd", x"de", 
        x"de", x"df", x"e0", x"e0", x"e1", x"e0", x"e1", x"e0", x"df", x"de", x"de", x"de", x"d9", x"d9", x"de", 
        x"e0", x"e8", x"d8", x"d4", x"da", x"e7", x"da", x"da", x"d9", x"df", x"de", x"de", x"df", x"d9", x"e0", 
        x"e2", x"e2", x"e0", x"e5", x"dc", x"da", x"db", x"de", x"de", x"df", x"de", x"e8", x"9e", x"b4", x"e2", 
        x"dd", x"db", x"de", x"dd", x"dc", x"dc", x"e5", x"d2", x"dd", x"e3", x"de", x"de", x"e0", x"e0", x"de", 
        x"dd", x"e0", x"e5", x"e9", x"e6", x"e1", x"df", x"df", x"de", x"d5", x"dc", x"e0", x"e2", x"e5", x"e6", 
        x"eb", x"e9", x"e9", x"e2", x"e6", x"e1", x"e6", x"e6", x"e7", x"e7", x"e3", x"e4", x"e9", x"eb", x"e8", 
        x"e5", x"e1", x"e6", x"e5", x"e2", x"e1", x"e5", x"e1", x"a3", x"b3", x"eb", x"e3", x"e3", x"e5", x"e8", 
        x"e5", x"e0", x"e7", x"ea", x"e7", x"e2", x"e2", x"e4", x"e4", x"e2", x"e3", x"e4", x"e3", x"e4", x"e2", 
        x"e1", x"de", x"e2", x"e2", x"de", x"df", x"e2", x"e2", x"e2", x"e1", x"df", x"e1", x"e5", x"e0", x"e0", 
        x"e0", x"e1", x"df", x"dc", x"e0", x"e2", x"e6", x"de", x"e5", x"e3", x"e5", x"e3", x"e6", x"e7", x"e3", 
        x"e4", x"e3", x"e2", x"e3", x"df", x"e2", x"e7", x"e4", x"e1", x"e4", x"e4", x"e3", x"e1", x"e9", x"ce", 
        x"b4", x"da", x"de", x"dd", x"e0", x"e0", x"e6", x"e1", x"e0", x"e6", x"e4", x"e5", x"e4", x"e2", x"e6", 
        x"dd", x"c2", x"d6", x"e7", x"e9", x"e7", x"e5", x"e4", x"e3", x"e7", x"e5", x"e4", x"e8", x"e6", x"e4", 
        x"e5", x"e1", x"e2", x"e2", x"e3", x"e2", x"df", x"df", x"e2", x"e0", x"dd", x"dd", x"db", x"da", x"de", 
        x"dc", x"db", x"da", x"d9", x"d9", x"dd", x"de", x"db", x"db", x"dc", x"dc", x"d9", x"d6", x"d7", x"d9", 
        x"d9", x"d9", x"d9", x"d9", x"da", x"db", x"db", x"d9", x"da", x"db", x"d4", x"d5", x"d5", x"d5", x"cd", 
        x"cd", x"d1", x"d3", x"d3", x"d2", x"d2", x"d0", x"d1", x"d2", x"d2", x"de", x"dd", x"d0", x"cd", x"de", 
        x"dc", x"d1", x"d1", x"d3", x"d4", x"d2", x"d3", x"d2", x"d0", x"d1", x"cc", x"cc", x"cc", x"cc", x"cd", 
        x"d7", x"d8", x"d9", x"d3", x"cb", x"c9", x"c8", x"c4", x"c5", x"c4", x"c1", x"be", x"c1", x"c6", x"c6", 
        x"ca", x"c8", x"ce", x"e0", x"d4", x"c7", x"d3", x"dc", x"c8", x"c5", x"c7", x"c6", x"c5", x"c4", x"c5", 
        x"c5", x"c0", x"c1", x"c3", x"c8", x"cf", x"cb", x"c6", x"c3", x"c3", x"c3", x"c2", x"c1", x"c3", x"c7", 
        x"cc", x"d2", x"d3", x"d1", x"cc", x"cb", x"db", x"dc", x"ca", x"cf", x"e1", x"d1", x"cb", x"cc", x"d0", 
        x"d0", x"cf", x"d1", x"d1", x"d1", x"d2", x"d4", x"d7", x"d7", x"d6", x"d3", x"d2", x"d3", x"d4", x"d7", 
        x"d9", x"d9", x"d9", x"dd", x"de", x"e2", x"eb", x"e8", x"e6", x"ee", x"e9", x"e5", x"e5", x"e6", x"e5", 
        x"e4", x"e6", x"e7", x"e5", x"e8", x"eb", x"ec", x"ee", x"f2", x"f0", x"f0", x"f0", x"f0", x"ef", x"f0", 
        x"f2", x"f3", x"f3", x"f3", x"f2", x"f5", x"f4", x"f4", x"fa", x"f6", x"f5", x"f5", x"f4", x"f8", x"f9", 
        x"f8", x"f7", x"f8", x"f7", x"f7", x"f8", x"f8", x"f7", x"f5", x"f6", x"f7", x"f8", x"f7", x"f6", x"f5", 
        x"f7", x"f7", x"f4", x"f3", x"f4", x"f5", x"f6", x"f4", x"f3", x"f4", x"f4", x"f5", x"f5", x"f5", x"f4", 
        x"f4", x"f4", x"f3", x"f2", x"f2", x"f2", x"f5", x"f6", x"f3", x"f4", x"f3", x"f0", x"f1", x"f1", x"f1", 
        x"f1", x"ef", x"ef", x"f0", x"f2", x"f2", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f0", x"f0", x"ee", x"ed", x"ee", x"ee", x"ef", x"ee", 
        x"ec", x"eb", x"ec", x"ee", x"f0", x"ec", x"ed", x"f5", x"b2", x"3d", x"64", x"a5", x"8b", x"8a", x"8e", 
        x"89", x"85", x"82", x"83", x"82", x"81", x"7f", x"7d", x"7b", x"7a", x"79", x"7a", x"77", x"74", x"73", 
        x"70", x"6f", x"6d", x"6e", x"70", x"6e", x"6a", x"68", x"69", x"69", x"66", x"63", x"67", x"3a", x"20", 
        x"4e", x"6e", x"69", x"67", x"63", x"62", x"64", x"63", x"63", x"56", x"40", x"41", x"44", x"3f", x"2c", 
        x"39", x"52", x"41", x"42", x"50", x"59", x"57", x"5b", x"5d", x"54", x"4a", x"50", x"52", x"58", x"52", 
        x"26", x"27", x"59", x"66", x"63", x"5f", x"5a", x"5a", x"5a", x"52", x"52", x"4e", x"3b", x"46", x"6c", 
        x"76", x"42", x"33", x"4c", x"48", x"48", x"4e", x"4d", x"51", x"53", x"53", x"54", x"52", x"52", x"5f", 
        x"60", x"56", x"4d", x"4e", x"4d", x"4a", x"46", x"46", x"5a", x"9c", x"ac", x"b4", x"ca", x"d6", x"da", 
        x"dd", x"df", x"e6", x"cd", x"63", x"30", x"29", x"21", x"1c", x"19", x"17", x"18", x"16", x"2c", x"47", 
        x"43", x"43", x"42", x"4a", x"4e", x"4f", x"52", x"52", x"30", x"17", x"10", x"29", x"3c", x"27", x"19", 
        x"45", x"46", x"36", x"50", x"a0", x"65", x"3f", x"4a", x"52", x"65", x"4f", x"4c", x"5f", x"67", x"3c", 
        x"22", x"2d", x"3e", x"4a", x"6a", x"a4", x"a3", x"a3", x"a3", x"9f", x"b0", x"e0", x"df", x"e1", x"dd", 
        x"de", x"dc", x"da", x"a6", x"7c", x"a7", x"b7", x"9f", x"7b", x"bc", x"df", x"d9", x"d9", x"d9", x"d9", 
        x"da", x"db", x"d8", x"e3", x"bb", x"7a", x"92", x"a7", x"93", x"7a", x"c0", x"dd", x"dd", x"de", x"d9", 
        x"ce", x"dd", x"df", x"dd", x"de", x"b3", x"81", x"95", x"9e", x"84", x"94", x"dc", x"dd", x"db", x"dd", 
        x"de", x"de", x"dd", x"dd", x"db", x"8d", x"b4", x"e2", x"db", x"e0", x"de", x"dc", x"dc", x"dc", x"e1", 
        x"bf", x"8b", x"8e", x"92", x"8e", x"c4", x"e4", x"e1", x"e0", x"dd", x"de", x"de", x"de", x"de", x"de", 
        x"df", x"df", x"df", x"df", x"e0", x"df", x"df", x"e0", x"df", x"df", x"de", x"dc", x"db", x"dc", x"db", 
        x"ab", x"9d", x"8e", x"82", x"94", x"cd", x"dd", x"dd", x"dd", x"db", x"df", x"de", x"db", x"e0", x"cb", 
        x"96", x"8b", x"90", x"be", x"df", x"dd", x"de", x"df", x"db", x"e0", x"dd", x"cb", x"70", x"78", x"bb", 
        x"db", x"dc", x"dd", x"dc", x"dd", x"dd", x"e2", x"c6", x"d6", x"e2", x"dd", x"de", x"e0", x"df", x"dd", 
        x"de", x"de", x"bc", x"a6", x"b5", x"da", x"df", x"dc", x"e1", x"da", x"e0", x"e2", x"e2", x"dc", x"cf", 
        x"c3", x"ad", x"bf", x"de", x"e6", x"e4", x"e4", x"e5", x"e6", x"e6", x"e6", x"e2", x"c7", x"b7", x"c8", 
        x"e2", x"e7", x"e3", x"e4", x"e4", x"e3", x"e4", x"e0", x"a4", x"b6", x"ea", x"e3", x"e5", x"e6", x"e5", 
        x"e3", x"e4", x"d9", x"c8", x"ce", x"e3", x"e4", x"e2", x"e6", x"e5", x"e3", x"e4", x"e6", x"e5", x"e5", 
        x"e4", x"e2", x"e3", x"e2", x"e2", x"e3", x"e1", x"de", x"e2", x"e2", x"e3", x"dc", x"d7", x"e0", x"e4", 
        x"e0", x"e7", x"e5", x"e0", x"e1", x"e3", x"e4", x"e4", x"e3", x"e4", x"e6", x"e7", x"e7", x"e4", x"e3", 
        x"e3", x"e6", x"e7", x"e2", x"e1", x"e2", x"e2", x"e4", x"e3", x"e1", x"e3", x"e3", x"e2", x"e7", x"b7", 
        x"b0", x"e1", x"e5", x"e5", x"e0", x"da", x"e3", x"e0", x"e6", x"e5", x"e1", x"e6", x"e3", x"e2", x"e4", 
        x"de", x"c7", x"d8", x"e3", x"e1", x"e5", x"e7", x"e2", x"e4", x"e4", x"e5", x"e6", x"e2", x"e4", x"e4", 
        x"e3", x"e9", x"e7", x"e5", x"e2", x"e6", x"e3", x"e3", x"e5", x"e4", x"e5", x"e5", x"e6", x"e5", x"e0", 
        x"e3", x"e3", x"e3", x"e1", x"df", x"e1", x"e7", x"e8", x"e7", x"e8", x"e8", x"e6", x"e4", x"e3", x"e4", 
        x"e4", x"e3", x"e4", x"e4", x"e5", x"e5", x"e5", x"e5", x"e6", x"e8", x"ea", x"e9", x"c4", x"d2", x"e3", 
        x"e5", x"e9", x"e6", x"e2", x"e6", x"e8", x"e3", x"e2", x"e7", x"e1", x"e0", x"e1", x"e1", x"e3", x"df", 
        x"e1", x"e1", x"e3", x"e1", x"e3", x"e6", x"c9", x"d2", x"df", x"e2", x"e1", x"d3", x"c7", x"df", x"e2", 
        x"e2", x"e6", x"df", x"ca", x"df", x"e0", x"dd", x"df", x"e0", x"c8", x"dc", x"e1", x"df", x"dd", x"de", 
        x"df", x"df", x"e0", x"e1", x"dd", x"dc", x"de", x"e1", x"dd", x"e0", x"e1", x"de", x"de", x"da", x"da", 
        x"d9", x"d8", x"d6", x"d8", x"dd", x"de", x"dc", x"d9", x"d6", x"d6", x"d9", x"d7", x"d3", x"d5", x"d5", 
        x"d8", x"d9", x"d9", x"d6", x"d4", x"d2", x"de", x"df", x"cf", x"d5", x"e0", x"d4", x"d0", x"d1", x"d6", 
        x"d4", x"d1", x"cf", x"ce", x"cf", x"d1", x"d5", x"d7", x"d6", x"d5", x"d1", x"ce", x"cd", x"cd", x"ce", 
        x"ce", x"cd", x"ca", x"c9", x"c8", x"d1", x"de", x"d6", x"d4", x"e1", x"d5", x"cf", x"ce", x"ce", x"c9", 
        x"c6", x"c6", x"c3", x"be", x"c2", x"c5", x"c4", x"c4", x"c9", x"c8", x"c8", x"c9", x"cb", x"cc", x"ce", 
        x"cf", x"cd", x"cd", x"d0", x"d3", x"df", x"d9", x"d9", x"e5", x"db", x"d7", x"dd", x"e1", x"de", x"d6", 
        x"d4", x"d4", x"d4", x"d3", x"d1", x"cd", x"ca", x"c9", x"c8", x"c8", x"c9", x"cc", x"d1", x"d5", x"db", 
        x"e8", x"dc", x"e3", x"e4", x"d9", x"db", x"dc", x"dc", x"db", x"db", x"dc", x"df", x"e2", x"e5", x"e5", 
        x"e4", x"e4", x"e5", x"e5", x"e6", x"e8", x"e7", x"ea", x"ef", x"e9", x"eb", x"ee", x"e9", x"eb", x"ee", 
        x"ef", x"ed", x"ed", x"ed", x"ed", x"ec", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"f0", x"f1", x"ed", x"f1", x"ee", x"ec", x"ed", x"ed", x"ec", x"ec", x"ee", x"f0", x"ef", x"ee", x"ef", 
        x"ef", x"ee", x"ee", x"ef", x"f0", x"ee", x"ee", x"f5", x"bd", x"3b", x"5e", x"c1", x"9a", x"87", x"8c", 
        x"8a", x"87", x"83", x"81", x"7f", x"80", x"7e", x"7c", x"7b", x"7a", x"79", x"78", x"77", x"73", x"70", 
        x"73", x"71", x"72", x"72", x"74", x"73", x"6e", x"6c", x"6c", x"6c", x"69", x"66", x"68", x"3a", x"1f", 
        x"49", x"6b", x"68", x"66", x"62", x"5e", x"5e", x"5d", x"5f", x"55", x"3d", x"3e", x"40", x"3d", x"2d", 
        x"38", x"53", x"41", x"40", x"4f", x"58", x"57", x"59", x"58", x"53", x"4d", x"54", x"50", x"51", x"4e", 
        x"24", x"22", x"54", x"63", x"5d", x"58", x"53", x"4f", x"4c", x"46", x"44", x"3e", x"41", x"89", x"c2", 
        x"c1", x"81", x"47", x"43", x"48", x"44", x"41", x"45", x"47", x"47", x"47", x"46", x"42", x"3f", x"51", 
        x"5c", x"4f", x"40", x"40", x"44", x"44", x"40", x"48", x"61", x"a0", x"b1", x"b8", x"cc", x"d9", x"dc", 
        x"e1", x"e2", x"ea", x"d5", x"77", x"44", x"4a", x"47", x"4a", x"4b", x"4a", x"4b", x"48", x"58", x"73", 
        x"70", x"6f", x"6b", x"6b", x"6d", x"71", x"73", x"74", x"58", x"41", x"3b", x"50", x"60", x"39", x"1a", 
        x"49", x"43", x"26", x"3d", x"79", x"4f", x"4e", x"4f", x"36", x"43", x"69", x"89", x"82", x"65", x"59", 
        x"5f", x"31", x"50", x"83", x"7a", x"a6", x"a3", x"a4", x"a4", x"9e", x"af", x"e1", x"e1", x"e1", x"dc", 
        x"dc", x"de", x"ca", x"7c", x"af", x"e0", x"e2", x"db", x"94", x"95", x"d7", x"dc", x"db", x"d9", x"db", 
        x"dd", x"dd", x"de", x"d9", x"88", x"92", x"d8", x"d9", x"d8", x"9b", x"9d", x"dd", x"d8", x"dd", x"da", 
        x"d0", x"da", x"db", x"df", x"ce", x"85", x"9a", x"dc", x"de", x"ce", x"7f", x"b4", x"de", x"dc", x"dd", 
        x"df", x"de", x"de", x"df", x"dc", x"8b", x"b2", x"e3", x"db", x"df", x"dd", x"e0", x"dd", x"e0", x"d4", 
        x"89", x"a7", x"db", x"d8", x"9e", x"8f", x"db", x"e2", x"e0", x"dd", x"e0", x"de", x"de", x"de", x"de", 
        x"df", x"df", x"de", x"de", x"df", x"de", x"dd", x"de", x"df", x"de", x"e0", x"db", x"d9", x"de", x"dc", 
        x"80", x"72", x"bd", x"c6", x"97", x"93", x"dc", x"dc", x"de", x"e3", x"dc", x"d8", x"e3", x"d1", x"8c", 
        x"9a", x"be", x"a8", x"8d", x"cb", x"de", x"db", x"db", x"dd", x"df", x"de", x"d5", x"7b", x"81", x"c8", 
        x"df", x"dd", x"dd", x"dd", x"df", x"e6", x"e6", x"8f", x"c3", x"df", x"dc", x"de", x"df", x"de", x"df", 
        x"e0", x"ac", x"7c", x"93", x"89", x"98", x"d9", x"de", x"de", x"dd", x"e1", x"e0", x"e4", x"c5", x"79", 
        x"8a", x"9b", x"7e", x"b5", x"e7", x"e5", x"e5", x"e6", x"e1", x"e2", x"e4", x"b2", x"88", x"94", x"8c", 
        x"ad", x"e7", x"e5", x"e2", x"e0", x"e1", x"e3", x"e1", x"a9", x"b9", x"e9", x"e1", x"e2", x"e3", x"e5", 
        x"ea", x"cd", x"92", x"7f", x"81", x"b7", x"e5", x"e8", x"e5", x"e4", x"e4", x"e4", x"e6", x"e4", x"e5", 
        x"e5", x"e4", x"e2", x"e0", x"e2", x"e5", x"e2", x"e3", x"e2", x"e5", x"cd", x"9c", x"89", x"a4", x"d7", 
        x"ea", x"e1", x"e0", x"e3", x"e3", x"db", x"c2", x"e8", x"e3", x"cf", x"d0", x"e7", x"e3", x"e3", x"e4", 
        x"e4", x"d5", x"c3", x"ac", x"9b", x"cc", x"e8", x"e4", x"e1", x"e0", x"df", x"e2", x"e3", x"d7", x"a4", 
        x"ac", x"db", x"e6", x"e3", x"dd", x"da", x"e8", x"e7", x"dd", x"cc", x"d0", x"e3", x"e5", x"e4", x"e1", 
        x"e5", x"e0", x"e2", x"e2", x"e2", x"e5", x"e4", x"e7", x"e4", x"cf", x"ca", x"df", x"ea", x"e6", x"e3", 
        x"e2", x"ea", x"e4", x"e0", x"e4", x"e7", x"df", x"e4", x"e3", x"e5", x"e5", x"e6", x"e5", x"e0", x"e6", 
        x"e5", x"e3", x"df", x"e3", x"e6", x"e4", x"e1", x"e2", x"e6", x"e6", x"e4", x"e4", x"e3", x"e3", x"e2", 
        x"e3", x"e4", x"e4", x"e4", x"e5", x"e5", x"e5", x"e5", x"e4", x"e6", x"e7", x"e5", x"ac", x"c7", x"e8", 
        x"e1", x"e7", x"e4", x"e4", x"e4", x"e4", x"ea", x"e6", x"e8", x"e6", x"e6", x"e3", x"e3", x"e7", x"e1", 
        x"e1", x"e4", x"e2", x"e1", x"e3", x"e9", x"aa", x"c3", x"e4", x"e6", x"e7", x"cc", x"b1", x"de", x"e2", 
        x"e7", x"e6", x"d1", x"aa", x"e1", x"e6", x"e5", x"e3", x"db", x"a6", x"d3", x"e6", x"e6", x"e2", x"e4", 
        x"e7", x"e7", x"e7", x"e0", x"e1", x"e2", x"e1", x"e4", x"e6", x"e5", x"e2", x"e3", x"e4", x"e6", x"e4", 
        x"d7", x"dd", x"e5", x"e2", x"e3", x"e4", x"e6", x"e4", x"e1", x"df", x"e2", x"e3", x"e1", x"e3", x"e2", 
        x"e2", x"e3", x"e4", x"e4", x"e6", x"e2", x"e0", x"e0", x"e0", x"e4", x"d4", x"cf", x"db", x"e3", x"e9", 
        x"e9", x"e8", x"e5", x"e4", x"e6", x"e9", x"ed", x"ef", x"ed", x"ec", x"ea", x"e8", x"e7", x"e7", x"e7", 
        x"e7", x"e6", x"e4", x"e5", x"e3", x"e3", x"e7", x"e2", x"df", x"e5", x"e4", x"e1", x"e1", x"e2", x"e3", 
        x"e0", x"de", x"de", x"dc", x"de", x"dd", x"dd", x"db", x"dc", x"dd", x"dd", x"dd", x"de", x"df", x"df", 
        x"de", x"de", x"df", x"e3", x"d7", x"e1", x"e4", x"df", x"e9", x"e2", x"dd", x"e3", x"e9", x"e4", x"d8", 
        x"d9", x"db", x"da", x"d9", x"d6", x"d2", x"cf", x"cd", x"cf", x"cc", x"c9", x"c8", x"cb", x"d0", x"d5", 
        x"de", x"d2", x"d9", x"dc", x"d0", x"d2", x"d2", x"d5", x"d4", x"cf", x"c9", x"c6", x"c4", x"c4", x"c4", 
        x"c5", x"c7", x"c9", x"c9", x"cc", x"ce", x"cd", x"d3", x"da", x"cd", x"d1", x"d5", x"c7", x"c7", x"c3", 
        x"c5", x"c6", x"c7", x"c9", x"c9", x"c6", x"c8", x"c9", x"ca", x"cb", x"cd", x"cd", x"cd", x"c9", x"cb", 
        x"d7", x"db", x"d4", x"d7", x"ce", x"c8", x"c8", x"ca", x"cb", x"cd", x"d0", x"d4", x"d8", x"dc", x"dd", 
        x"dd", x"dc", x"db", x"db", x"dc", x"de", x"e4", x"f0", x"bc", x"3e", x"5d", x"c4", x"ae", x"85", x"88", 
        x"89", x"86", x"82", x"80", x"80", x"7f", x"7f", x"7f", x"7d", x"7b", x"7b", x"77", x"77", x"78", x"70", 
        x"77", x"72", x"71", x"70", x"71", x"72", x"6e", x"6d", x"6c", x"6a", x"69", x"6c", x"6d", x"3d", x"21", 
        x"44", x"65", x"68", x"67", x"65", x"5f", x"5c", x"5d", x"61", x"5a", x"41", x"3f", x"3f", x"3c", x"2d", 
        x"33", x"4f", x"3f", x"3f", x"50", x"59", x"59", x"5b", x"5a", x"56", x"52", x"56", x"51", x"53", x"4f", 
        x"27", x"22", x"51", x"66", x"62", x"5b", x"55", x"4b", x"47", x"46", x"44", x"3a", x"2b", x"5f", x"8b", 
        x"99", x"b6", x"7b", x"46", x"43", x"40", x"41", x"45", x"42", x"41", x"42", x"44", x"45", x"42", x"54", 
        x"65", x"57", x"46", x"44", x"47", x"4b", x"48", x"4a", x"5e", x"9d", x"b3", x"b9", x"cc", x"dc", x"e1", 
        x"da", x"be", x"c3", x"d2", x"85", x"48", x"42", x"39", x"41", x"46", x"43", x"41", x"38", x"49", x"76", 
        x"78", x"7a", x"77", x"75", x"76", x"77", x"78", x"7a", x"62", x"4c", x"47", x"59", x"6c", x"43", x"19", 
        x"45", x"39", x"2e", x"49", x"97", x"64", x"46", x"3f", x"25", x"20", x"3c", x"4b", x"41", x"78", x"81", 
        x"76", x"49", x"39", x"4b", x"61", x"a4", x"a4", x"a3", x"a4", x"9c", x"ac", x"e0", x"e1", x"e0", x"e1", 
        x"dd", x"e1", x"b8", x"67", x"a2", x"b7", x"b7", x"b8", x"88", x"7f", x"d0", x"de", x"da", x"dc", x"de", 
        x"db", x"db", x"e0", x"cc", x"82", x"ba", x"e2", x"de", x"dd", x"d5", x"d0", x"df", x"db", x"dd", x"dc", 
        x"d5", x"db", x"d9", x"e2", x"bd", x"84", x"c0", x"e0", x"db", x"e1", x"a0", x"8d", x"dc", x"db", x"dc", 
        x"dd", x"dc", x"dc", x"dd", x"dd", x"8e", x"b3", x"e5", x"df", x"de", x"de", x"dd", x"e1", x"e2", x"be", 
        x"78", x"c2", x"d9", x"dd", x"ba", x"6d", x"d0", x"e0", x"e0", x"e0", x"df", x"dd", x"de", x"dd", x"dd", 
        x"de", x"df", x"df", x"e1", x"e1", x"df", x"dc", x"de", x"de", x"dc", x"dc", x"df", x"db", x"db", x"df", 
        x"8b", x"ab", x"dd", x"e6", x"b6", x"76", x"d9", x"e2", x"de", x"dd", x"df", x"df", x"dd", x"d2", x"ab", 
        x"d3", x"e3", x"cd", x"7f", x"c8", x"e2", x"da", x"de", x"e0", x"de", x"dd", x"e3", x"99", x"a9", x"de", 
        x"df", x"df", x"dd", x"de", x"dd", x"df", x"e8", x"8b", x"be", x"df", x"de", x"de", x"de", x"df", x"e2", 
        x"ce", x"82", x"c6", x"dd", x"c9", x"8f", x"b9", x"e7", x"df", x"db", x"dd", x"e1", x"e7", x"bd", x"76", 
        x"c2", x"e3", x"ad", x"9e", x"e3", x"e4", x"e3", x"e6", x"e3", x"e6", x"db", x"9e", x"bb", x"dd", x"bb", 
        x"93", x"dd", x"e4", x"e4", x"e4", x"e4", x"e4", x"e3", x"a5", x"b5", x"ee", x"e3", x"e4", x"e6", x"e3", 
        x"e4", x"ac", x"9d", x"d3", x"bd", x"93", x"c7", x"ea", x"e3", x"e2", x"e2", x"e4", x"e6", x"e7", x"e6", 
        x"e3", x"e2", x"df", x"e0", x"e1", x"e0", x"e3", x"e1", x"e1", x"e0", x"a6", x"9c", x"bb", x"95", x"b7", 
        x"e4", x"df", x"e4", x"e2", x"e2", x"d0", x"98", x"e4", x"e3", x"b5", x"b3", x"e5", x"e2", x"e6", x"e1", 
        x"e7", x"af", x"76", x"a2", x"a2", x"98", x"cf", x"e8", x"df", x"e1", x"e2", x"e4", x"d7", x"a0", x"8f", 
        x"90", x"a0", x"de", x"e3", x"e2", x"de", x"e8", x"da", x"9b", x"7f", x"bb", x"e1", x"e2", x"e5", x"e6", 
        x"de", x"b2", x"c9", x"e4", x"e3", x"e4", x"e5", x"e4", x"b6", x"88", x"88", x"af", x"e4", x"e6", x"e6", 
        x"e6", x"e6", x"c9", x"bf", x"e8", x"d4", x"ba", x"de", x"e3", x"e3", x"e4", x"e1", x"bb", x"9c", x"c4", 
        x"e1", x"e0", x"e1", x"e4", x"d7", x"a7", x"8a", x"af", x"e0", x"ea", x"e6", x"e4", x"e5", x"e4", x"e2", 
        x"e3", x"e4", x"e5", x"e5", x"e4", x"e4", x"e4", x"e4", x"e7", x"e0", x"b0", x"a9", x"92", x"cb", x"e9", 
        x"e6", x"e4", x"e6", x"e3", x"c4", x"b8", x"d0", x"e5", x"e4", x"e1", x"e5", x"e4", x"e4", x"e4", x"e6", 
        x"e3", x"e4", x"e2", x"e4", x"e5", x"e7", x"aa", x"c0", x"e3", x"e4", x"e5", x"d6", x"bb", x"e3", x"e6", 
        x"e4", x"e3", x"c7", x"b1", x"e3", x"e5", x"e1", x"e4", x"e4", x"a4", x"d4", x"e5", x"e3", x"e2", x"e2", 
        x"dd", x"ce", x"da", x"e4", x"e3", x"e0", x"e0", x"e2", x"dc", x"d6", x"de", x"e6", x"e2", x"e8", x"dd", 
        x"b6", x"c3", x"e8", x"e3", x"e4", x"e5", x"e2", x"de", x"e4", x"e2", x"e4", x"e6", x"e0", x"dc", x"e4", 
        x"e4", x"e2", x"e2", x"e4", x"e5", x"e1", x"e4", x"e5", x"e4", x"ea", x"dc", x"db", x"ea", x"ea", x"e7", 
        x"e8", x"e8", x"e8", x"e8", x"e9", x"ec", x"f0", x"f2", x"f1", x"f0", x"ea", x"e8", x"e9", x"ea", x"ec", 
        x"e8", x"e8", x"ec", x"ea", x"e7", x"e9", x"e8", x"e6", x"e6", x"e8", x"e6", x"e6", x"e5", x"e6", x"e7", 
        x"e6", x"e4", x"e4", x"e5", x"e0", x"d4", x"df", x"e5", x"e3", x"e5", x"e4", x"e4", x"e5", x"e6", x"e6", 
        x"e5", x"e8", x"e3", x"e4", x"c7", x"cd", x"ec", x"ea", x"eb", x"e9", x"e8", x"eb", x"ee", x"eb", x"e6", 
        x"e9", x"e7", x"e7", x"e7", x"e6", x"e6", x"e7", x"e7", x"e6", x"e5", x"e5", x"e5", x"e4", x"e4", x"e4", 
        x"e5", x"e4", x"e4", x"e8", x"e9", x"e8", x"e9", x"eb", x"ea", x"e7", x"e4", x"e4", x"e4", x"e5", x"e5", 
        x"e7", x"e5", x"e3", x"e2", x"e5", x"e8", x"ea", x"e7", x"e6", x"db", x"d9", x"df", x"d6", x"d6", x"d5", 
        x"d8", x"d3", x"d0", x"d6", x"d4", x"ce", x"d6", x"d6", x"d6", x"d7", x"d7", x"d6", x"d5", x"d1", x"d0", 
        x"d7", x"d9", x"d2", x"da", x"d5", x"d0", x"cf", x"cc", x"cc", x"cc", x"c8", x"c6", x"c6", x"c7", x"c7", 
        x"c6", x"c4", x"c3", x"c3", x"c6", x"c9", x"d5", x"e6", x"a6", x"33", x"55", x"aa", x"a5", x"6e", x"66", 
        x"68", x"61", x"5e", x"5f", x"5e", x"5a", x"5b", x"5e", x"59", x"55", x"58", x"56", x"58", x"60", x"5a", 
        x"63", x"5c", x"55", x"54", x"55", x"58", x"57", x"56", x"54", x"50", x"4c", x"4b", x"55", x"34", x"21", 
        x"3e", x"53", x"51", x"4c", x"4a", x"44", x"40", x"42", x"46", x"40", x"25", x"24", x"25", x"26", x"29", 
        x"34", x"49", x"2a", x"29", x"39", x"41", x"3b", x"3b", x"3c", x"39", x"3a", x"39", x"34", x"3b", x"3b", 
        x"22", x"21", x"4d", x"66", x"62", x"55", x"4f", x"49", x"45", x"3f", x"3c", x"40", x"32", x"4f", x"92", 
        x"bf", x"bf", x"67", x"2f", x"3f", x"3c", x"3a", x"40", x"42", x"41", x"42", x"43", x"47", x"44", x"4f", 
        x"61", x"56", x"45", x"3f", x"3e", x"3f", x"3d", x"42", x"58", x"99", x"b3", x"bd", x"d0", x"d2", x"ab", 
        x"5e", x"2e", x"32", x"8a", x"8a", x"4a", x"42", x"37", x"41", x"46", x"45", x"44", x"3f", x"4f", x"78", 
        x"77", x"76", x"75", x"75", x"76", x"78", x"77", x"7c", x"64", x"4b", x"44", x"54", x"6a", x"45", x"20", 
        x"4b", x"3f", x"28", x"4b", x"a0", x"55", x"2c", x"3a", x"23", x"1e", x"25", x"24", x"21", x"47", x"60", 
        x"56", x"44", x"3f", x"31", x"61", x"a5", x"a7", x"a4", x"a1", x"9d", x"ae", x"e1", x"e2", x"df", x"e1", 
        x"de", x"e0", x"b3", x"5a", x"79", x"86", x"87", x"83", x"84", x"aa", x"d6", x"dd", x"db", x"dc", x"db", 
        x"dc", x"da", x"e1", x"c0", x"84", x"c3", x"df", x"db", x"d9", x"de", x"dd", x"dc", x"db", x"de", x"da", 
        x"d4", x"da", x"da", x"e0", x"b4", x"87", x"cb", x"de", x"d8", x"df", x"b0", x"77", x"d7", x"dc", x"de", 
        x"e0", x"dd", x"dd", x"df", x"dd", x"91", x"b1", x"e5", x"dd", x"de", x"dd", x"dc", x"e0", x"e1", x"b1", 
        x"4f", x"72", x"79", x"7c", x"72", x"6d", x"d0", x"df", x"e0", x"df", x"dc", x"dc", x"de", x"dc", x"dc", 
        x"df", x"e0", x"de", x"df", x"e0", x"de", x"dc", x"de", x"e0", x"de", x"e0", x"e1", x"de", x"dc", x"dd", 
        x"92", x"ba", x"e0", x"df", x"bd", x"77", x"d6", x"df", x"dd", x"de", x"dc", x"dc", x"db", x"e1", x"d5", 
        x"af", x"97", x"83", x"66", x"c4", x"e0", x"db", x"db", x"db", x"dc", x"dc", x"e1", x"9e", x"a6", x"de", 
        x"dd", x"dc", x"de", x"de", x"dc", x"de", x"eb", x"8c", x"bd", x"df", x"de", x"dd", x"de", x"dd", x"df", 
        x"b6", x"8f", x"dd", x"de", x"e0", x"a4", x"a4", x"e4", x"de", x"db", x"df", x"e3", x"e6", x"c1", x"90", 
        x"da", x"ea", x"c6", x"97", x"df", x"e5", x"e6", x"e5", x"e3", x"e5", x"e5", x"df", x"cf", x"ba", x"97", 
        x"7d", x"de", x"e3", x"e2", x"e4", x"e2", x"e3", x"e2", x"aa", x"b3", x"f0", x"e5", x"e4", x"e3", x"e3", 
        x"e4", x"8f", x"a7", x"bf", x"b9", x"83", x"af", x"e9", x"e2", x"e1", x"e3", x"e4", x"e5", x"e7", x"e9", 
        x"e5", x"e2", x"e2", x"e2", x"e1", x"e0", x"df", x"e3", x"e4", x"e4", x"a4", x"a2", x"d3", x"d5", x"d3", 
        x"e4", x"e1", x"e6", x"e3", x"e3", x"d2", x"98", x"e3", x"e0", x"b5", x"b0", x"e6", x"e4", x"e3", x"e6", 
        x"e6", x"b0", x"91", x"e1", x"e9", x"99", x"af", x"e1", x"e4", x"e2", x"e1", x"e4", x"b6", x"97", x"d5", 
        x"d6", x"88", x"c5", x"e8", x"e4", x"dd", x"e8", x"dd", x"85", x"b8", x"e7", x"e6", x"e4", x"e4", x"e4", 
        x"e2", x"a7", x"c2", x"e5", x"e4", x"e3", x"e4", x"d6", x"9c", x"bd", x"d4", x"9e", x"ce", x"e9", x"e3", 
        x"e4", x"ea", x"bf", x"aa", x"e7", x"cd", x"a3", x"dc", x"e4", x"e3", x"e5", x"df", x"8e", x"8f", x"da", 
        x"e5", x"e2", x"e3", x"e3", x"b7", x"9c", x"c9", x"9e", x"c2", x"e9", x"e3", x"e2", x"e7", x"e4", x"e3", 
        x"e2", x"e4", x"e6", x"e6", x"e5", x"e4", x"e6", x"e7", x"e3", x"ab", x"9f", x"a6", x"6f", x"c6", x"ea", 
        x"e5", x"e5", x"eb", x"c2", x"95", x"9f", x"92", x"d4", x"eb", x"e4", x"e7", x"e5", x"e4", x"e6", x"e6", 
        x"e5", x"e4", x"e5", x"e5", x"e3", x"ea", x"b7", x"c2", x"e5", x"e8", x"e6", x"e1", x"e0", x"e3", x"e4", 
        x"eb", x"c6", x"90", x"8e", x"ac", x"e3", x"e5", x"e3", x"e5", x"ac", x"ce", x"e8", x"e2", x"e3", x"d9", 
        x"a4", x"85", x"a4", x"dc", x"e5", x"e2", x"e3", x"db", x"9d", x"86", x"ad", x"df", x"e1", x"e4", x"da", 
        x"95", x"9d", x"e9", x"e2", x"e4", x"de", x"a8", x"a8", x"de", x"e5", x"e6", x"df", x"a9", x"99", x"c9", 
        x"e9", x"e2", x"e3", x"e2", x"b8", x"9a", x"b5", x"e1", x"e6", x"e5", x"dd", x"d3", x"eb", x"e7", x"e7", 
        x"e1", x"b2", x"ab", x"c5", x"e8", x"e9", x"ec", x"e8", x"e6", x"e6", x"d8", x"e3", x"e6", x"e8", x"df", 
        x"ba", x"c2", x"e5", x"e9", x"e5", x"e7", x"e8", x"e7", x"e5", x"e8", x"e5", x"e2", x"e9", x"e6", x"ca", 
        x"c5", x"e1", x"e7", x"e8", x"d7", x"ad", x"ce", x"ea", x"e6", x"e5", x"e5", x"e5", x"e5", x"e5", x"e5", 
        x"e5", x"e7", x"de", x"c4", x"b7", x"cc", x"ef", x"ec", x"ed", x"da", x"d2", x"ea", x"ec", x"e7", x"e8", 
        x"e9", x"e8", x"e5", x"e5", x"e5", x"e6", x"ea", x"e0", x"de", x"e8", x"e5", x"e5", x"e6", x"df", x"e3", 
        x"e5", x"e6", x"e6", x"e8", x"e1", x"e6", x"e8", x"e8", x"ea", x"e8", x"e4", x"e6", x"e9", x"e8", x"ea", 
        x"ec", x"df", x"e9", x"e7", x"ec", x"eb", x"ea", x"e6", x"e7", x"e4", x"df", x"df", x"de", x"df", x"e2", 
        x"e5", x"cd", x"c5", x"df", x"dc", x"c6", x"df", x"e1", x"e0", x"e1", x"e2", x"e2", x"e0", x"e3", x"e1", 
        x"da", x"df", x"e2", x"d5", x"d6", x"e5", x"e6", x"d1", x"d9", x"e7", x"e5", x"e4", x"e5", x"e6", x"e5", 
        x"e5", x"e4", x"e5", x"e2", x"e6", x"e8", x"e8", x"ef", x"ad", x"36", x"4f", x"b3", x"d1", x"a8", x"81", 
        x"7f", x"7c", x"7c", x"7b", x"7b", x"79", x"74", x"75", x"6d", x"69", x"6f", x"6e", x"62", x"61", x"62", 
        x"6b", x"69", x"69", x"66", x"63", x"63", x"5e", x"5e", x"57", x"52", x"5b", x"54", x"58", x"3b", x"20", 
        x"3b", x"56", x"59", x"5f", x"53", x"51", x"52", x"51", x"4e", x"44", x"27", x"24", x"29", x"28", x"2c", 
        x"32", x"4d", x"30", x"29", x"34", x"48", x"45", x"45", x"43", x"44", x"44", x"40", x"3a", x"40", x"3c", 
        x"21", x"20", x"48", x"4d", x"3f", x"32", x"30", x"27", x"26", x"23", x"25", x"27", x"1d", x"25", x"65", 
        x"b5", x"a2", x"48", x"1c", x"20", x"21", x"24", x"23", x"28", x"23", x"21", x"20", x"21", x"24", x"20", 
        x"20", x"26", x"1f", x"20", x"1f", x"1d", x"1b", x"2a", x"4c", x"8c", x"a7", x"b9", x"c9", x"81", x"20", 
        x"0a", x"08", x"09", x"24", x"6e", x"49", x"3c", x"38", x"3c", x"3e", x"40", x"40", x"3c", x"49", x"71", 
        x"74", x"70", x"71", x"71", x"71", x"71", x"6e", x"77", x"63", x"43", x"3f", x"4e", x"65", x"45", x"23", 
        x"3b", x"34", x"2f", x"32", x"7a", x"50", x"2b", x"35", x"23", x"1e", x"26", x"1d", x"16", x"2f", x"5c", 
        x"6f", x"75", x"6e", x"74", x"7b", x"a2", x"a1", x"a4", x"a2", x"9e", x"ad", x"df", x"e0", x"de", x"de", 
        x"de", x"df", x"ba", x"77", x"c4", x"e2", x"db", x"e0", x"d1", x"c8", x"d9", x"df", x"d7", x"d7", x"db", 
        x"dd", x"d9", x"de", x"cd", x"82", x"b6", x"e1", x"dc", x"df", x"cd", x"b8", x"d6", x"dd", x"dd", x"da", 
        x"d6", x"dd", x"dd", x"e1", x"b9", x"82", x"c4", x"e2", x"da", x"e6", x"a4", x"80", x"d8", x"db", x"dc", 
        x"de", x"dd", x"dd", x"df", x"db", x"94", x"b0", x"e3", x"df", x"dd", x"dd", x"dd", x"dd", x"de", x"ba", 
        x"73", x"bc", x"cd", x"cc", x"ca", x"c1", x"df", x"df", x"de", x"de", x"de", x"de", x"dd", x"dc", x"dd", 
        x"e0", x"e0", x"de", x"de", x"df", x"dd", x"db", x"de", x"df", x"de", x"de", x"de", x"dd", x"db", x"dc", 
        x"94", x"b9", x"de", x"dd", x"bc", x"76", x"d5", x"de", x"db", x"dc", x"dc", x"e1", x"dc", x"ce", x"8b", 
        x"8f", x"ab", x"b6", x"83", x"c2", x"e2", x"dc", x"da", x"dd", x"dd", x"de", x"e2", x"a4", x"a2", x"dc", 
        x"dc", x"dd", x"e0", x"df", x"df", x"de", x"e6", x"8f", x"c0", x"e2", x"de", x"dc", x"dd", x"dd", x"e1", 
        x"b5", x"8f", x"df", x"df", x"e2", x"a5", x"a1", x"e1", x"e1", x"da", x"de", x"e4", x"e3", x"c2", x"97", 
        x"dc", x"e9", x"cb", x"94", x"e1", x"e7", x"e5", x"e4", x"e5", x"e5", x"e0", x"ae", x"93", x"94", x"90", 
        x"80", x"dc", x"e8", x"e4", x"e1", x"e4", x"e6", x"e1", x"ac", x"b2", x"ef", x"e6", x"e3", x"e1", x"e5", 
        x"e1", x"7f", x"8b", x"99", x"9b", x"97", x"c9", x"e6", x"e4", x"e4", x"e4", x"e5", x"e5", x"e5", x"e7", 
        x"e5", x"e2", x"e3", x"e3", x"e3", x"e2", x"e2", x"e5", x"e2", x"e7", x"d4", x"98", x"93", x"a6", x"d0", 
        x"e3", x"e6", x"e2", x"e5", x"e4", x"d4", x"92", x"e4", x"e6", x"b1", x"b0", x"e4", x"e5", x"e5", x"e5", 
        x"e2", x"b9", x"a4", x"e3", x"ea", x"aa", x"ab", x"e0", x"e6", x"e3", x"e1", x"e6", x"a9", x"7a", x"a5", 
        x"a7", x"7e", x"c1", x"e8", x"e3", x"e0", x"e4", x"db", x"98", x"ca", x"e6", x"e2", x"e4", x"e5", x"e4", 
        x"e5", x"a6", x"bd", x"e8", x"e5", x"e5", x"e7", x"ca", x"8a", x"a9", x"b3", x"8d", x"c8", x"e4", x"e3", 
        x"e5", x"eb", x"c2", x"af", x"e2", x"d2", x"a1", x"de", x"e5", x"e6", x"e9", x"dc", x"a5", x"bf", x"ec", 
        x"e2", x"e1", x"df", x"de", x"a5", x"95", x"c6", x"9d", x"b6", x"e3", x"e6", x"e4", x"e4", x"e2", x"e4", 
        x"e4", x"e5", x"e4", x"e5", x"e7", x"e7", x"e6", x"e8", x"d8", x"a0", x"ce", x"e5", x"9f", x"c4", x"e7", 
        x"e5", x"e6", x"e7", x"ab", x"ac", x"bd", x"90", x"c0", x"e6", x"e5", x"e4", x"e4", x"e4", x"e3", x"e5", 
        x"e5", x"e4", x"e4", x"e3", x"e2", x"eb", x"b7", x"c0", x"e5", x"e6", x"e4", x"e3", x"e3", x"e7", x"e4", 
        x"e8", x"ab", x"b6", x"bf", x"93", x"d3", x"e7", x"e2", x"e4", x"ab", x"cb", x"e6", x"e5", x"e5", x"c5", 
        x"a0", x"c5", x"9f", x"c3", x"e4", x"e2", x"e3", x"c3", x"a2", x"c6", x"b5", x"d7", x"e5", x"e2", x"e3", 
        x"ae", x"b4", x"ec", x"e1", x"e1", x"d2", x"8b", x"c1", x"e3", x"df", x"e3", x"c3", x"a7", x"b7", x"a5", 
        x"db", x"e6", x"e4", x"da", x"9d", x"a8", x"a8", x"d0", x"e8", x"e5", x"d2", x"b6", x"e6", x"ea", x"e9", 
        x"c4", x"a8", x"a5", x"8e", x"e1", x"f0", x"ed", x"d5", x"d4", x"cf", x"ba", x"df", x"ea", x"ea", x"c2", 
        x"9d", x"a6", x"cb", x"e9", x"e6", x"e7", x"e8", x"e8", x"e7", x"e7", x"e3", x"e2", x"ed", x"d0", x"a4", 
        x"9f", x"c4", x"e7", x"e6", x"d7", x"a9", x"c7", x"e8", x"e9", x"e6", x"e6", x"e6", x"e6", x"e5", x"e5", 
        x"e5", x"e6", x"be", x"9d", x"92", x"c0", x"ed", x"ed", x"da", x"b1", x"a2", x"cf", x"ec", x"e8", x"e5", 
        x"e9", x"e9", x"e3", x"e4", x"e8", x"e7", x"d8", x"b1", x"b7", x"e0", x"e4", x"e6", x"d4", x"af", x"b2", 
        x"de", x"e8", x"ea", x"c6", x"ac", x"d0", x"e8", x"e7", x"e9", x"e8", x"e6", x"e7", x"e9", x"e8", x"e9", 
        x"c8", x"ad", x"d5", x"e8", x"ed", x"e3", x"be", x"b3", x"d9", x"e2", x"df", x"cb", x"af", x"bf", x"e1", 
        x"e6", x"ce", x"c8", x"de", x"e3", x"cc", x"db", x"e3", x"dc", x"bb", x"ba", x"dd", x"e0", x"e1", x"c6", 
        x"b9", x"da", x"e5", x"c2", x"b6", x"db", x"e4", x"d7", x"dc", x"e2", x"e0", x"ca", x"cb", x"e1", x"e2", 
        x"e0", x"c8", x"ce", x"e5", x"e8", x"e1", x"d2", x"e6", x"b8", x"3b", x"46", x"aa", x"d5", x"c1", x"8d", 
        x"75", x"7d", x"7d", x"78", x"73", x"6e", x"74", x"72", x"6c", x"6b", x"6d", x"69", x"5a", x"60", x"68", 
        x"6d", x"67", x"67", x"64", x"64", x"5e", x"5c", x"62", x"5c", x"59", x"5e", x"54", x"57", x"3b", x"20", 
        x"3d", x"5c", x"50", x"50", x"56", x"54", x"48", x"4a", x"51", x"48", x"27", x"25", x"27", x"23", x"29", 
        x"31", x"47", x"2c", x"26", x"34", x"42", x"3f", x"45", x"43", x"42", x"41", x"41", x"3e", x"41", x"3e", 
        x"25", x"1f", x"49", x"53", x"46", x"31", x"24", x"28", x"2c", x"2a", x"2a", x"2a", x"25", x"18", x"3f", 
        x"64", x"3f", x"25", x"34", x"39", x"26", x"21", x"26", x"29", x"2d", x"2a", x"30", x"2d", x"25", x"1b", 
        x"14", x"1e", x"2a", x"2d", x"32", x"32", x"29", x"30", x"48", x"88", x"a5", x"b5", x"bf", x"79", x"1d", 
        x"17", x"15", x"11", x"1f", x"54", x"33", x"1f", x"24", x"1d", x"1a", x"1a", x"1b", x"1b", x"2d", x"60", 
        x"69", x"65", x"63", x"60", x"63", x"63", x"5f", x"64", x"51", x"2b", x"23", x"2f", x"4a", x"3e", x"1f", 
        x"33", x"36", x"34", x"4b", x"97", x"64", x"32", x"37", x"28", x"39", x"26", x"2a", x"37", x"34", x"59", 
        x"92", x"81", x"7c", x"72", x"64", x"a1", x"a4", x"a2", x"a2", x"9e", x"ad", x"df", x"e1", x"df", x"df", 
        x"de", x"d9", x"d1", x"7e", x"97", x"d8", x"dc", x"d1", x"95", x"9f", x"d9", x"db", x"db", x"db", x"db", 
        x"da", x"d9", x"dc", x"db", x"90", x"93", x"d1", x"e0", x"d7", x"95", x"8d", x"d6", x"dc", x"de", x"db", 
        x"d6", x"df", x"dd", x"e0", x"d0", x"86", x"9b", x"dc", x"dc", x"d2", x"7e", x"a6", x"dd", x"da", x"da", 
        x"dd", x"dc", x"dd", x"de", x"da", x"90", x"ae", x"e2", x"de", x"de", x"dd", x"de", x"db", x"e1", x"c7", 
        x"7b", x"b4", x"e7", x"e8", x"c5", x"98", x"d3", x"e2", x"e0", x"d8", x"df", x"de", x"dc", x"db", x"dc", 
        x"de", x"de", x"dc", x"de", x"de", x"dc", x"db", x"dd", x"de", x"de", x"de", x"dd", x"dd", x"dd", x"de", 
        x"90", x"b7", x"de", x"df", x"bc", x"74", x"d3", x"e1", x"da", x"dc", x"df", x"dc", x"de", x"b4", x"77", 
        x"dd", x"ed", x"d2", x"7b", x"c2", x"dd", x"db", x"dc", x"d8", x"da", x"e2", x"e0", x"a7", x"a2", x"e1", 
        x"db", x"db", x"dd", x"de", x"df", x"df", x"ea", x"8f", x"bc", x"e0", x"dd", x"db", x"dd", x"dc", x"e1", 
        x"c7", x"83", x"d8", x"e6", x"e0", x"9e", x"a5", x"e6", x"e1", x"da", x"dd", x"e1", x"e5", x"c4", x"95", 
        x"d9", x"e7", x"cd", x"8e", x"df", x"e4", x"e2", x"e3", x"e3", x"ea", x"d0", x"7e", x"bf", x"e4", x"c7", 
        x"84", x"d9", x"e6", x"e3", x"e2", x"e2", x"e1", x"e2", x"ad", x"af", x"ed", x"e2", x"e3", x"e7", x"e6", 
        x"df", x"9b", x"b7", x"e5", x"e5", x"ca", x"d6", x"e3", x"e2", x"e5", x"e2", x"e2", x"e4", x"e4", x"e6", 
        x"e4", x"e2", x"e3", x"e4", x"e3", x"e2", x"e4", x"e0", x"e1", x"e4", x"d8", x"d9", x"be", x"91", x"a3", 
        x"eb", x"e5", x"e5", x"e5", x"e4", x"d5", x"93", x"e0", x"e7", x"b4", x"ae", x"e7", x"e6", x"e4", x"e4", 
        x"e1", x"b7", x"a1", x"e6", x"eb", x"a9", x"ae", x"e3", x"e2", x"e0", x"e6", x"e6", x"ab", x"86", x"ac", 
        x"b1", x"a5", x"d9", x"e8", x"e2", x"e1", x"e6", x"dc", x"9c", x"cd", x"e4", x"e3", x"e6", x"e4", x"e0", 
        x"e5", x"a5", x"bc", x"e6", x"e4", x"e8", x"e6", x"c9", x"87", x"9c", x"a5", x"a4", x"d3", x"e4", x"e7", 
        x"e4", x"e6", x"c2", x"ae", x"e6", x"d5", x"9b", x"d8", x"e6", x"e4", x"e9", x"e0", x"ad", x"c9", x"e9", 
        x"e3", x"e2", x"e6", x"dd", x"9b", x"79", x"9c", x"95", x"c3", x"e4", x"e4", x"e4", x"e4", x"e1", x"e5", 
        x"e6", x"e5", x"e3", x"e5", x"e8", x"e8", x"e6", x"e9", x"cf", x"a1", x"d7", x"ed", x"ba", x"bf", x"ec", 
        x"e7", x"e6", x"e5", x"a3", x"87", x"94", x"89", x"c1", x"e5", x"e3", x"e3", x"e4", x"e3", x"e5", x"e6", 
        x"e6", x"e4", x"e4", x"e2", x"e3", x"ec", x"b5", x"be", x"e6", x"e5", x"e3", x"e4", x"e5", x"e3", x"e4", 
        x"e5", x"9c", x"97", x"a6", x"98", x"d0", x"e6", x"e0", x"e3", x"a9", x"c7", x"e6", x"e8", x"e9", x"bf", 
        x"87", x"a2", x"90", x"c1", x"e6", x"e3", x"de", x"bb", x"b9", x"eb", x"e3", x"e5", x"e5", x"e3", x"e2", 
        x"b7", x"ba", x"e9", x"e4", x"e9", x"d4", x"a5", x"dd", x"e9", x"e4", x"df", x"b4", x"be", x"e1", x"a2", 
        x"d2", x"e6", x"e8", x"db", x"b6", x"d7", x"b3", x"c9", x"ea", x"e7", x"d3", x"b7", x"e7", x"e4", x"e5", 
        x"bc", x"cc", x"dc", x"a2", x"dc", x"f3", x"ee", x"d0", x"cf", x"d0", x"b5", x"e0", x"eb", x"e5", x"ac", 
        x"aa", x"aa", x"b4", x"e7", x"e6", x"e6", x"e7", x"e7", x"e6", x"e7", x"e6", x"e5", x"ea", x"bd", x"a1", 
        x"ae", x"a7", x"e2", x"e3", x"e0", x"c1", x"d8", x"ea", x"e5", x"e6", x"e6", x"e5", x"e5", x"e6", x"e6", 
        x"e6", x"e6", x"ad", x"cc", x"c3", x"c2", x"ee", x"f1", x"c6", x"a9", x"a9", x"b8", x"eb", x"e9", x"e4", 
        x"e6", x"e6", x"e7", x"e5", x"e3", x"e9", x"cd", x"a3", x"bc", x"da", x"e6", x"e9", x"b7", x"ab", x"9c", 
        x"d2", x"e9", x"e3", x"b6", x"a8", x"cd", x"ea", x"e8", x"e8", x"e9", x"e8", x"e9", x"ea", x"e9", x"e8", 
        x"bf", x"a8", x"b9", x"e7", x"ef", x"cd", x"a2", x"a2", x"c2", x"df", x"e4", x"ae", x"98", x"a3", x"d3", 
        x"e7", x"d2", x"c9", x"dc", x"de", x"b6", x"d7", x"e1", x"cb", x"9c", x"a2", x"d4", x"e4", x"da", x"a9", 
        x"9c", x"ca", x"e7", x"c0", x"b1", x"dc", x"e4", x"cb", x"cd", x"e3", x"d3", x"9f", x"a1", x"d2", x"e5", 
        x"d1", x"9a", x"a7", x"e1", x"ed", x"c9", x"a5", x"d5", x"bc", x"38", x"3e", x"9b", x"d3", x"d0", x"a3", 
        x"6f", x"6e", x"7c", x"79", x"6b", x"60", x"6c", x"71", x"69", x"68", x"6c", x"68", x"53", x"60", x"6a", 
        x"62", x"57", x"64", x"67", x"60", x"4d", x"51", x"62", x"5d", x"57", x"5e", x"56", x"59", x"3e", x"20", 
        x"3b", x"5e", x"41", x"3b", x"52", x"52", x"37", x"3c", x"52", x"50", x"2a", x"26", x"28", x"2a", x"2a", 
        x"2f", x"45", x"2c", x"39", x"43", x"3c", x"37", x"40", x"43", x"36", x"31", x"3c", x"41", x"41", x"3e", 
        x"23", x"1d", x"47", x"4c", x"4b", x"3a", x"19", x"25", x"2f", x"2a", x"2f", x"28", x"2e", x"30", x"12", 
        x"0b", x"10", x"30", x"63", x"6f", x"52", x"36", x"25", x"2a", x"34", x"31", x"2a", x"29", x"17", x"10", 
        x"12", x"3b", x"60", x"37", x"24", x"30", x"23", x"2e", x"42", x"81", x"a7", x"b0", x"cb", x"ba", x"55", 
        x"3f", x"4b", x"28", x"34", x"5e", x"3b", x"19", x"29", x"25", x"22", x"21", x"26", x"24", x"2c", x"63", 
        x"6a", x"68", x"6a", x"61", x"66", x"6d", x"6b", x"6a", x"5a", x"30", x"26", x"35", x"52", x"44", x"21", 
        x"48", x"57", x"5b", x"7f", x"9e", x"5e", x"40", x"38", x"20", x"31", x"2e", x"55", x"66", x"52", x"68", 
        x"6f", x"42", x"3c", x"65", x"78", x"a0", x"a5", x"a3", x"a3", x"9f", x"ad", x"de", x"df", x"df", x"de", 
        x"e0", x"da", x"d8", x"c1", x"80", x"89", x"94", x"81", x"85", x"cb", x"e0", x"da", x"db", x"db", x"d9", 
        x"da", x"db", x"d9", x"e4", x"c7", x"81", x"82", x"91", x"86", x"82", x"c7", x"e2", x"da", x"df", x"db", 
        x"d3", x"dc", x"da", x"dc", x"e4", x"b7", x"82", x"92", x"93", x"7e", x"8d", x"d8", x"df", x"d9", x"da", 
        x"dd", x"dd", x"dd", x"dc", x"d8", x"94", x"b4", x"e0", x"da", x"de", x"dd", x"db", x"da", x"da", x"de", 
        x"ad", x"7e", x"90", x"94", x"81", x"a3", x"df", x"dc", x"dc", x"dd", x"dc", x"dc", x"dd", x"dc", x"da", 
        x"da", x"db", x"dd", x"df", x"de", x"dd", x"dc", x"dd", x"de", x"de", x"dd", x"dc", x"da", x"da", x"da", 
        x"95", x"b4", x"dc", x"de", x"bb", x"7d", x"cc", x"df", x"db", x"dd", x"dc", x"dd", x"de", x"c3", x"7d", 
        x"a3", x"ae", x"95", x"62", x"9d", x"d5", x"dd", x"dc", x"d7", x"d9", x"da", x"de", x"ae", x"88", x"c2", 
        x"dd", x"db", x"db", x"e0", x"dc", x"dd", x"e6", x"8d", x"b9", x"dc", x"dc", x"dc", x"de", x"da", x"de", 
        x"dd", x"92", x"96", x"bd", x"a9", x"85", x"be", x"e5", x"db", x"d7", x"de", x"df", x"e5", x"c5", x"92", 
        x"d6", x"e9", x"cf", x"8a", x"d5", x"e3", x"e2", x"e3", x"e2", x"e6", x"d4", x"88", x"ae", x"c3", x"91", 
        x"64", x"bf", x"e3", x"df", x"e2", x"e4", x"e3", x"e2", x"ac", x"aa", x"eb", x"e0", x"e3", x"e4", x"de", 
        x"e8", x"ba", x"83", x"b9", x"b0", x"92", x"c6", x"e9", x"e4", x"e3", x"e4", x"e4", x"e5", x"e5", x"e6", 
        x"e3", x"e1", x"e2", x"e3", x"e2", x"e1", x"df", x"e2", x"e5", x"e7", x"ac", x"a7", x"d7", x"b4", x"9a", 
        x"e7", x"e1", x"e5", x"e2", x"e3", x"dc", x"91", x"bc", x"cb", x"88", x"a2", x"e6", x"e5", x"e6", x"e4", 
        x"e9", x"b5", x"79", x"c7", x"d6", x"93", x"b6", x"e6", x"e4", x"df", x"e1", x"e4", x"c1", x"9a", x"d2", 
        x"da", x"a3", x"cd", x"e5", x"e2", x"da", x"e4", x"de", x"98", x"cc", x"e5", x"e2", x"e2", x"e3", x"e4", 
        x"e8", x"a5", x"ba", x"e5", x"df", x"e1", x"e6", x"d3", x"a4", x"c5", x"e9", x"ba", x"cd", x"eb", x"e3", 
        x"e5", x"e8", x"c9", x"ab", x"dc", x"c3", x"8e", x"da", x"e3", x"e2", x"e3", x"de", x"a6", x"c0", x"e9", 
        x"e1", x"dd", x"e9", x"e2", x"b2", x"a7", x"e9", x"c8", x"c9", x"e0", x"e6", x"e7", x"e7", x"e4", x"e5", 
        x"e4", x"e4", x"e5", x"e6", x"e6", x"e6", x"e6", x"e9", x"d8", x"a5", x"cd", x"e9", x"a5", x"bd", x"e9", 
        x"e6", x"e8", x"e6", x"aa", x"b4", x"d9", x"c3", x"d1", x"e9", x"e5", x"e3", x"e4", x"e2", x"e5", x"e6", 
        x"e7", x"e6", x"e4", x"e4", x"e5", x"ed", x"b4", x"b9", x"e4", x"e5", x"e1", x"e5", x"e6", x"e5", x"e2", 
        x"e7", x"ad", x"b1", x"cd", x"c2", x"dc", x"e8", x"e3", x"e6", x"a9", x"c3", x"e7", x"e6", x"e7", x"c1", 
        x"97", x"c0", x"b7", x"d3", x"e5", x"e3", x"e3", x"bd", x"ac", x"e9", x"cf", x"d8", x"e3", x"e4", x"e2", 
        x"bc", x"b5", x"eb", x"e3", x"e8", x"d2", x"a9", x"de", x"e6", x"e2", x"e2", x"ba", x"bf", x"e7", x"9d", 
        x"cc", x"e7", x"e4", x"dd", x"b9", x"da", x"b6", x"c6", x"e9", x"e8", x"d6", x"b4", x"e8", x"e6", x"e7", 
        x"be", x"cf", x"e6", x"ac", x"df", x"e9", x"ef", x"ce", x"c7", x"d2", x"b4", x"e2", x"e7", x"e4", x"aa", 
        x"95", x"ab", x"c8", x"e7", x"e4", x"e4", x"e5", x"e4", x"e5", x"e7", x"e5", x"e6", x"ed", x"bf", x"99", 
        x"aa", x"b8", x"e4", x"e5", x"df", x"ba", x"cf", x"e9", x"e7", x"e6", x"e6", x"e6", x"e6", x"e6", x"e6", 
        x"e6", x"e1", x"b1", x"dc", x"db", x"c5", x"ec", x"ef", x"c5", x"9d", x"9f", x"c3", x"e9", x"e7", x"e8", 
        x"e6", x"e9", x"e5", x"e8", x"ea", x"e9", x"db", x"ac", x"b0", x"dc", x"e7", x"e8", x"af", x"9e", x"9f", 
        x"d6", x"ea", x"ec", x"cb", x"af", x"cc", x"ec", x"ea", x"e8", x"e8", x"e8", x"e8", x"ea", x"eb", x"ec", 
        x"c5", x"a2", x"b5", x"ec", x"eb", x"d6", x"ca", x"cc", x"bf", x"da", x"e6", x"b9", x"d2", x"c3", x"c7", 
        x"e8", x"d4", x"c7", x"df", x"e7", x"b2", x"d3", x"e1", x"c3", x"c7", x"e3", x"de", x"e4", x"e1", x"b5", 
        x"9c", x"c8", x"e9", x"cc", x"c1", x"df", x"e6", x"c8", x"c5", x"e7", x"c8", x"b2", x"b5", x"c9", x"e3", 
        x"d1", x"b9", x"bd", x"da", x"eb", x"c8", x"a8", x"da", x"bf", x"39", x"41", x"97", x"d0", x"d1", x"c7", 
        x"90", x"6b", x"7d", x"7a", x"6a", x"6c", x"68", x"74", x"6a", x"67", x"6d", x"6a", x"57", x"64", x"69", 
        x"5e", x"57", x"65", x"67", x"62", x"5c", x"52", x"5e", x"5c", x"51", x"5d", x"54", x"58", x"42", x"22", 
        x"36", x"5d", x"48", x"4f", x"5a", x"56", x"39", x"41", x"52", x"4f", x"51", x"64", x"67", x"58", x"38", 
        x"2d", x"40", x"5c", x"84", x"7d", x"5c", x"3d", x"37", x"46", x"34", x"2a", x"3b", x"43", x"41", x"3f", 
        x"27", x"1f", x"45", x"41", x"3d", x"3c", x"1b", x"20", x"2a", x"31", x"2c", x"26", x"62", x"6d", x"26", 
        x"24", x"36", x"4f", x"65", x"63", x"76", x"81", x"45", x"22", x"29", x"26", x"17", x"12", x"0d", x"0a", 
        x"1d", x"92", x"be", x"63", x"15", x"25", x"1f", x"24", x"33", x"7f", x"a7", x"a7", x"c4", x"cf", x"7e", 
        x"47", x"83", x"7e", x"8f", x"7c", x"48", x"22", x"26", x"30", x"2f", x"26", x"2c", x"2f", x"30", x"61", 
        x"5c", x"5a", x"65", x"58", x"59", x"69", x"6c", x"6d", x"5e", x"2a", x"1a", x"2a", x"45", x"43", x"20", 
        x"38", x"43", x"45", x"59", x"9d", x"75", x"63", x"4e", x"25", x"39", x"4f", x"47", x"4a", x"5f", x"64", 
        x"43", x"46", x"65", x"6f", x"74", x"a4", x"a4", x"a5", x"a5", x"a0", x"ae", x"de", x"de", x"dd", x"df", 
        x"de", x"d5", x"d5", x"dc", x"ca", x"a9", x"a2", x"ac", x"ce", x"dc", x"db", x"de", x"d9", x"d9", x"da", 
        x"dc", x"da", x"d8", x"de", x"e1", x"ce", x"a9", x"9c", x"a5", x"c9", x"dc", x"dd", x"db", x"dc", x"d8", 
        x"cf", x"da", x"d9", x"db", x"df", x"de", x"c2", x"a3", x"9b", x"a1", x"ce", x"de", x"dc", x"d8", x"da", 
        x"dc", x"dc", x"dc", x"db", x"dd", x"be", x"cd", x"e0", x"db", x"dc", x"dc", x"db", x"dc", x"d8", x"e1", 
        x"dc", x"b4", x"9b", x"99", x"b5", x"d9", x"e1", x"db", x"df", x"e0", x"dc", x"dc", x"de", x"de", x"db", 
        x"da", x"dd", x"df", x"df", x"dd", x"de", x"de", x"dd", x"dd", x"dd", x"db", x"db", x"d9", x"da", x"db", 
        x"be", x"cb", x"da", x"de", x"cf", x"ac", x"d6", x"dd", x"dc", x"de", x"da", x"dc", x"df", x"d9", x"b4", 
        x"93", x"99", x"ac", x"a4", x"aa", x"d4", x"db", x"db", x"dc", x"db", x"d9", x"e1", x"d0", x"98", x"af", 
        x"d7", x"d9", x"da", x"db", x"dd", x"dd", x"e3", x"b2", x"c9", x"df", x"dd", x"dc", x"dc", x"d9", x"db", 
        x"de", x"cc", x"9b", x"93", x"90", x"b1", x"dc", x"de", x"dd", x"d7", x"db", x"e1", x"e1", x"d1", x"b3", 
        x"da", x"e5", x"db", x"af", x"dc", x"e2", x"e3", x"e6", x"e2", x"dd", x"e2", x"ba", x"95", x"99", x"a3", 
        x"9a", x"b9", x"e0", x"e3", x"e2", x"e2", x"e4", x"e2", x"c2", x"c0", x"e7", x"e2", x"e2", x"e0", x"e1", 
        x"e5", x"db", x"ab", x"95", x"93", x"b7", x"e0", x"e5", x"e1", x"e0", x"e2", x"e7", x"e6", x"e5", x"e6", 
        x"e3", x"e0", x"e1", x"e2", x"e2", x"e2", x"e0", x"e5", x"e3", x"e6", x"cb", x"9c", x"9f", x"9e", x"be", 
        x"e7", x"e4", x"e3", x"e1", x"e0", x"e4", x"bc", x"91", x"9b", x"92", x"b7", x"e3", x"e6", x"e4", x"e3", 
        x"e6", x"b6", x"72", x"9a", x"96", x"a1", x"d2", x"e5", x"e2", x"e3", x"e1", x"e5", x"dd", x"b2", x"9a", 
        x"97", x"99", x"da", x"e6", x"e3", x"dc", x"e4", x"e1", x"a9", x"cc", x"e2", x"e1", x"e1", x"e2", x"e3", 
        x"e4", x"b0", x"c2", x"e2", x"e3", x"e5", x"e5", x"e2", x"b5", x"94", x"95", x"9d", x"d7", x"e7", x"e2", 
        x"e3", x"e6", x"da", x"a7", x"9f", x"96", x"8f", x"d9", x"e2", x"e3", x"e6", x"df", x"b2", x"c5", x"e6", 
        x"e2", x"e1", x"df", x"e6", x"cc", x"9a", x"a2", x"98", x"c5", x"e3", x"e5", x"e3", x"e3", x"e4", x"e3", 
        x"e2", x"e3", x"e6", x"e6", x"e3", x"e3", x"e5", x"e6", x"e2", x"b5", x"a6", x"b0", x"7f", x"be", x"e7", 
        x"e3", x"e5", x"e8", x"c4", x"9f", x"aa", x"9e", x"ce", x"e6", x"e4", x"e3", x"e4", x"e1", x"e2", x"e5", 
        x"e7", x"e6", x"e3", x"e4", x"e5", x"eb", x"b8", x"b8", x"e0", x"e7", x"e5", x"e5", x"e3", x"e5", x"e5", 
        x"e9", x"be", x"a3", x"ac", x"a8", x"d8", x"ea", x"e4", x"e4", x"af", x"c4", x"e6", x"e6", x"e7", x"d1", 
        x"a7", x"b1", x"a6", x"cb", x"e5", x"e1", x"df", x"cd", x"99", x"ab", x"a1", x"d0", x"e5", x"e1", x"e3", 
        x"c2", x"a8", x"e5", x"e0", x"e4", x"d8", x"a5", x"dc", x"e4", x"e0", x"e3", x"c8", x"a6", x"b5", x"9a", 
        x"d6", x"e6", x"e3", x"de", x"b6", x"d5", x"b7", x"c5", x"e4", x"e9", x"da", x"ae", x"e3", x"e6", x"e9", 
        x"ca", x"b0", x"b8", x"91", x"db", x"e7", x"ed", x"d1", x"b0", x"ad", x"a9", x"e0", x"e7", x"e7", x"bb", 
        x"ae", x"bf", x"cc", x"e8", x"e6", x"e6", x"e5", x"e4", x"e6", x"e8", x"e6", x"e4", x"e9", x"cc", x"ab", 
        x"bb", x"bb", x"e4", x"e5", x"e3", x"bb", x"c7", x"eb", x"e4", x"e5", x"e5", x"e6", x"e6", x"e5", x"e5", 
        x"e5", x"e6", x"b6", x"c5", x"c0", x"b4", x"e6", x"ed", x"cc", x"b1", x"ba", x"ca", x"e9", x"e8", x"ea", 
        x"e7", x"e7", x"e5", x"e7", x"e5", x"e7", x"dd", x"b9", x"aa", x"cc", x"e7", x"eb", x"b5", x"b2", x"ae", 
        x"d8", x"e7", x"e9", x"d1", x"b2", x"bc", x"e7", x"ec", x"e9", x"e8", x"e8", x"e8", x"e9", x"eb", x"e1", 
        x"b3", x"ac", x"b4", x"e8", x"ef", x"d2", x"bb", x"bb", x"c3", x"db", x"e1", x"b9", x"bd", x"ba", x"cc", 
        x"e7", x"d2", x"c3", x"de", x"e6", x"b3", x"d2", x"e0", x"c6", x"b9", x"cd", x"da", x"e1", x"d9", x"ab", 
        x"a1", x"c3", x"e5", x"cb", x"c0", x"dd", x"e5", x"c9", x"c3", x"e5", x"c8", x"b7", x"bc", x"c9", x"e2", 
        x"d2", x"bf", x"c2", x"d8", x"ed", x"d6", x"af", x"cf", x"c1", x"3f", x"3d", x"94", x"d0", x"cd", x"d1", 
        x"b2", x"76", x"7a", x"7c", x"6c", x"73", x"67", x"75", x"6b", x"67", x"70", x"6b", x"59", x"66", x"6a", 
        x"60", x"58", x"62", x"67", x"64", x"65", x"56", x"60", x"62", x"51", x"5e", x"57", x"59", x"44", x"20", 
        x"31", x"5a", x"4a", x"45", x"56", x"59", x"3a", x"40", x"50", x"50", x"64", x"7e", x"7e", x"67", x"36", 
        x"26", x"37", x"5c", x"7a", x"75", x"61", x"38", x"34", x"46", x"36", x"2e", x"3e", x"46", x"43", x"41", 
        x"2b", x"21", x"47", x"42", x"30", x"34", x"23", x"22", x"22", x"2e", x"29", x"26", x"60", x"55", x"2d", 
        x"4f", x"5a", x"59", x"62", x"51", x"55", x"6d", x"4a", x"26", x"2a", x"27", x"1c", x"14", x"22", x"49", 
        x"5a", x"9b", x"a8", x"6a", x"1d", x"2b", x"28", x"28", x"3a", x"7a", x"a9", x"ab", x"c1", x"d3", x"aa", 
        x"62", x"6b", x"a8", x"aa", x"70", x"56", x"39", x"24", x"27", x"25", x"1f", x"24", x"23", x"27", x"5b", 
        x"5b", x"55", x"64", x"5a", x"5d", x"6b", x"69", x"6b", x"5e", x"27", x"15", x"28", x"40", x"41", x"1f", 
        x"38", x"47", x"41", x"44", x"a1", x"6f", x"69", x"70", x"53", x"4c", x"46", x"2e", x"3d", x"53", x"3c", 
        x"1e", x"42", x"68", x"72", x"78", x"9f", x"a8", x"a5", x"a4", x"a0", x"af", x"e1", x"e0", x"dc", x"e1", 
        x"df", x"d5", x"d6", x"d6", x"dc", x"e0", x"df", x"e0", x"df", x"da", x"da", x"d9", x"db", x"d8", x"d7", 
        x"d8", x"da", x"db", x"d9", x"da", x"df", x"dd", x"e1", x"dd", x"e4", x"de", x"db", x"db", x"da", x"d7", 
        x"cd", x"db", x"da", x"da", x"d9", x"db", x"e1", x"de", x"dc", x"e0", x"df", x"d9", x"d9", x"d8", x"da", 
        x"db", x"da", x"dc", x"da", x"dd", x"dd", x"dd", x"dc", x"dd", x"da", x"dc", x"db", x"de", x"dc", x"dc", 
        x"e0", x"e2", x"de", x"e1", x"e0", x"e2", x"e0", x"de", x"dd", x"d8", x"db", x"db", x"db", x"dc", x"dc", 
        x"db", x"dd", x"de", x"dc", x"db", x"dd", x"de", x"dc", x"db", x"db", x"db", x"dd", x"da", x"da", x"db", 
        x"de", x"dc", x"d9", x"db", x"dd", x"d8", x"df", x"dc", x"db", x"de", x"db", x"dc", x"dd", x"dd", x"de", 
        x"d1", x"ce", x"db", x"df", x"da", x"d6", x"da", x"db", x"dc", x"dc", x"dc", x"db", x"e4", x"d1", x"d0", 
        x"dd", x"dd", x"dc", x"d8", x"dc", x"dc", x"e0", x"d8", x"da", x"e0", x"dd", x"db", x"da", x"d9", x"d9", 
        x"db", x"df", x"d5", x"cc", x"d0", x"dd", x"dd", x"dd", x"e1", x"d6", x"d7", x"e2", x"e0", x"e2", x"dd", 
        x"e1", x"df", x"e7", x"e0", x"e9", x"e1", x"e1", x"e3", x"e2", x"e2", x"e2", x"e0", x"d2", x"cf", x"de", 
        x"dd", x"d7", x"e4", x"e1", x"de", x"e0", x"e0", x"e4", x"e2", x"e0", x"e3", x"e2", x"e3", x"df", x"e1", 
        x"e4", x"e5", x"e7", x"cf", x"d1", x"e5", x"e5", x"df", x"e3", x"e2", x"e4", x"e6", x"e2", x"e3", x"e5", 
        x"e2", x"e0", x"e1", x"e2", x"e3", x"e4", x"e1", x"e3", x"e4", x"e0", x"e4", x"d9", x"c5", x"d0", x"e1", 
        x"e4", x"e4", x"e1", x"e3", x"e0", x"e6", x"e0", x"c6", x"c7", x"d5", x"e1", x"e7", x"e5", x"e2", x"e5", 
        x"e4", x"be", x"98", x"c3", x"bb", x"d8", x"e8", x"e1", x"e2", x"e6", x"e2", x"de", x"e1", x"e0", x"c3", 
        x"bd", x"db", x"e1", x"e3", x"e2", x"df", x"e4", x"e6", x"d2", x"e1", x"e2", x"e2", x"e5", x"e2", x"e1", 
        x"e5", x"d4", x"d9", x"e2", x"e0", x"e2", x"e2", x"e3", x"db", x"c0", x"b4", x"d2", x"e8", x"e4", x"e1", 
        x"e7", x"e4", x"e8", x"d1", x"b5", x"bf", x"cb", x"e1", x"e4", x"e3", x"e3", x"e3", x"d3", x"da", x"e6", 
        x"e4", x"e1", x"e0", x"e3", x"e5", x"c9", x"a9", x"bd", x"e0", x"e4", x"e2", x"e4", x"e6", x"e5", x"e3", 
        x"e2", x"e2", x"e4", x"e4", x"e3", x"e3", x"e4", x"e3", x"e7", x"df", x"b1", x"aa", x"b6", x"d6", x"e6", 
        x"e3", x"e6", x"e4", x"e1", x"bd", x"a3", x"b7", x"df", x"e2", x"e1", x"e4", x"e5", x"e2", x"e2", x"e3", 
        x"e5", x"e3", x"e2", x"e4", x"e5", x"e8", x"d3", x"d2", x"e4", x"e6", x"e3", x"e5", x"e5", x"e7", x"e3", 
        x"e7", x"de", x"b3", x"9e", x"c7", x"e2", x"e3", x"e4", x"e7", x"cd", x"d5", x"e4", x"e3", x"e5", x"e8", 
        x"c4", x"9d", x"b3", x"d8", x"e2", x"de", x"de", x"dd", x"b7", x"98", x"b2", x"df", x"e4", x"e1", x"e4", 
        x"ce", x"af", x"db", x"e1", x"e2", x"dd", x"c4", x"dd", x"e2", x"e4", x"e2", x"dd", x"ab", x"9a", x"b8", 
        x"e2", x"e0", x"e7", x"dd", x"c9", x"e0", x"ca", x"d1", x"e4", x"e7", x"e1", x"c8", x"e5", x"e5", x"e9", 
        x"df", x"ae", x"a1", x"99", x"d9", x"ef", x"ea", x"e0", x"ae", x"9a", x"bc", x"e3", x"e6", x"e8", x"d8", 
        x"a5", x"9e", x"ce", x"e8", x"e7", x"e7", x"e7", x"e5", x"e6", x"e8", x"e7", x"e4", x"e6", x"dd", x"ac", 
        x"95", x"c0", x"e3", x"e1", x"e3", x"c5", x"c1", x"e2", x"e5", x"e5", x"e6", x"e6", x"e5", x"e5", x"e5", 
        x"e5", x"e9", x"ca", x"9e", x"9e", x"c3", x"e7", x"ea", x"de", x"ad", x"96", x"c4", x"e6", x"e8", x"e6", 
        x"e4", x"e4", x"e4", x"e5", x"e7", x"e6", x"d5", x"a7", x"a1", x"d0", x"e5", x"ea", x"cc", x"a1", x"a0", 
        x"df", x"e7", x"e8", x"c4", x"9e", x"bd", x"e8", x"ec", x"e9", x"e8", x"e8", x"e8", x"e7", x"ea", x"e2", 
        x"b5", x"9a", x"ae", x"e3", x"f1", x"d0", x"97", x"92", x"c9", x"e1", x"e0", x"b5", x"8d", x"9e", x"da", 
        x"e4", x"d0", x"c6", x"de", x"e3", x"b9", x"d0", x"dc", x"d0", x"9c", x"98", x"d0", x"e4", x"db", x"a5", 
        x"94", x"b4", x"e4", x"d3", x"b8", x"d6", x"e2", x"c7", x"c1", x"e4", x"d1", x"a3", x"9c", x"ca", x"e4", 
        x"d3", x"c0", x"c4", x"d7", x"e8", x"d0", x"a5", x"c0", x"c6", x"4a", x"3d", x"8f", x"ce", x"ca", x"cc", 
        x"c4", x"90", x"78", x"7b", x"6b", x"66", x"64", x"72", x"68", x"63", x"6e", x"6c", x"57", x"63", x"66", 
        x"5b", x"50", x"5d", x"69", x"5d", x"4f", x"4e", x"60", x"60", x"51", x"5a", x"58", x"5b", x"46", x"22", 
        x"34", x"5b", x"4e", x"39", x"4d", x"58", x"3f", x"42", x"4d", x"50", x"60", x"6f", x"6f", x"67", x"38", 
        x"26", x"36", x"5c", x"70", x"71", x"66", x"36", x"36", x"47", x"32", x"28", x"39", x"42", x"42", x"41", 
        x"2c", x"24", x"47", x"44", x"2d", x"32", x"23", x"20", x"24", x"2d", x"2d", x"23", x"2f", x"27", x"19", 
        x"32", x"44", x"50", x"67", x"54", x"32", x"30", x"35", x"33", x"2e", x"2c", x"24", x"1e", x"1f", x"60", 
        x"7b", x"9a", x"b1", x"70", x"23", x"27", x"25", x"2a", x"34", x"73", x"a8", x"aa", x"c4", x"d0", x"d8", 
        x"aa", x"51", x"67", x"62", x"49", x"55", x"4f", x"3d", x"2d", x"1d", x"1e", x"29", x"25", x"27", x"59", 
        x"62", x"56", x"64", x"5d", x"5e", x"69", x"68", x"6b", x"61", x"2d", x"19", x"2b", x"42", x"44", x"22", 
        x"3c", x"3d", x"32", x"43", x"7e", x"4c", x"36", x"52", x"56", x"4c", x"35", x"21", x"4d", x"6c", x"33", 
        x"41", x"49", x"30", x"4a", x"56", x"a0", x"aa", x"a6", x"a5", x"a2", x"b2", x"e2", x"e0", x"dd", x"df", 
        x"e0", x"dd", x"d5", x"d6", x"d4", x"d8", x"d7", x"dc", x"de", x"d9", x"da", x"db", x"db", x"dc", x"dd", 
        x"dd", x"dc", x"da", x"dc", x"da", x"dc", x"dd", x"de", x"df", x"de", x"de", x"db", x"db", x"dc", x"da", 
        x"d1", x"dd", x"da", x"d9", x"d6", x"d9", x"dc", x"dd", x"dc", x"dd", x"db", x"dc", x"da", x"d8", x"da", 
        x"d9", x"da", x"dd", x"dc", x"dc", x"df", x"dc", x"db", x"df", x"dc", x"dc", x"db", x"db", x"d9", x"da", 
        x"da", x"dd", x"e1", x"e0", x"de", x"e0", x"da", x"df", x"e0", x"e0", x"dc", x"d9", x"d3", x"d7", x"dc", 
        x"dc", x"da", x"db", x"da", x"da", x"dd", x"de", x"db", x"d9", x"da", x"db", x"dd", x"d8", x"d8", x"d9", 
        x"da", x"db", x"dd", x"da", x"d9", x"de", x"da", x"dd", x"da", x"dc", x"da", x"dc", x"d8", x"d9", x"d8", 
        x"da", x"dc", x"d6", x"da", x"db", x"d5", x"d7", x"d4", x"d6", x"d6", x"db", x"da", x"d7", x"d9", x"db", 
        x"da", x"d7", x"d9", x"d9", x"da", x"da", x"d9", x"da", x"dc", x"db", x"da", x"da", x"d9", x"da", x"da", 
        x"d9", x"d8", x"dc", x"de", x"dc", x"db", x"d7", x"d8", x"d9", x"d4", x"d6", x"e0", x"dd", x"e1", x"e0", 
        x"e1", x"e2", x"df", x"e1", x"e1", x"e2", x"e0", x"e0", x"e2", x"de", x"de", x"e2", x"e2", x"e4", x"e2", 
        x"e3", x"e3", x"e1", x"dd", x"df", x"de", x"e0", x"e1", x"e2", x"e2", x"de", x"df", x"e0", x"e2", x"e2", 
        x"df", x"e1", x"e3", x"e5", x"e3", x"e1", x"e1", x"e0", x"e1", x"e1", x"e2", x"e2", x"e1", x"e2", x"e3", 
        x"e1", x"e0", x"e1", x"e3", x"e3", x"e2", x"e1", x"e2", x"e2", x"e3", x"e1", x"e5", x"e5", x"e6", x"e4", 
        x"e1", x"e4", x"e0", x"e2", x"e3", x"de", x"e5", x"e5", x"e3", x"e7", x"e5", x"e3", x"e3", x"e6", x"e7", 
        x"e3", x"bb", x"a2", x"e2", x"e5", x"e3", x"e3", x"e2", x"e0", x"e0", x"e5", x"e3", x"e1", x"e1", x"e4", 
        x"e5", x"e6", x"e1", x"e1", x"e3", x"de", x"e3", x"e0", x"e0", x"e3", x"e3", x"e3", x"e3", x"e1", x"e2", 
        x"e3", x"e4", x"e3", x"e3", x"e0", x"e2", x"e0", x"e2", x"e4", x"ea", x"e6", x"e5", x"e5", x"e5", x"e0", 
        x"e4", x"e4", x"e4", x"e5", x"df", x"e5", x"e4", x"e5", x"de", x"e1", x"e0", x"e3", x"e4", x"e4", x"e4", 
        x"e2", x"e1", x"de", x"e5", x"e2", x"e2", x"e1", x"e3", x"e2", x"e2", x"e4", x"e3", x"e1", x"e2", x"e2", 
        x"e3", x"e2", x"e2", x"e2", x"e4", x"e5", x"e3", x"e5", x"e8", x"e8", x"e4", x"e0", x"e5", x"e6", x"e7", 
        x"e4", x"e2", x"e4", x"e2", x"e3", x"df", x"e2", x"e5", x"e3", x"e3", x"e2", x"e4", x"e5", x"e3", x"e1", 
        x"e3", x"e1", x"e1", x"e4", x"e4", x"e4", x"e6", x"e3", x"e4", x"e4", x"e4", x"e4", x"e2", x"e6", x"e6", 
        x"e3", x"e1", x"e2", x"dd", x"e6", x"e4", x"e3", x"e3", x"e5", x"e3", x"e2", x"e0", x"e3", x"e2", x"e3", 
        x"e1", x"de", x"e1", x"e2", x"e2", x"e0", x"dd", x"de", x"dd", x"da", x"df", x"e1", x"e0", x"e0", x"e0", 
        x"e1", x"d9", x"dd", x"df", x"df", x"e0", x"dc", x"e0", x"df", x"dd", x"de", x"e5", x"dd", x"d6", x"dd", 
        x"df", x"df", x"e0", x"e0", x"e1", x"e3", x"de", x"df", x"e5", x"e4", x"e7", x"e8", x"e8", x"e6", x"e3", 
        x"e5", x"e3", x"da", x"ab", x"d8", x"ed", x"e7", x"e8", x"e0", x"db", x"e4", x"e6", x"e6", x"e4", x"eb", 
        x"d9", x"da", x"e9", x"e6", x"e5", x"e6", x"e6", x"e4", x"e4", x"e6", x"e5", x"e5", x"e8", x"e8", x"e0", 
        x"d6", x"e4", x"e4", x"e7", x"e6", x"e0", x"dd", x"e4", x"e7", x"e6", x"e5", x"e5", x"e5", x"e5", x"e5", 
        x"e5", x"e5", x"e7", x"d5", x"dc", x"ec", x"ea", x"e5", x"e5", x"d8", x"ce", x"e0", x"e7", x"e6", x"e4", 
        x"e4", x"e4", x"e5", x"e6", x"e6", x"e5", x"e6", x"d6", x"d0", x"e3", x"e5", x"e2", x"e0", x"d3", x"cf", 
        x"e0", x"e3", x"e8", x"e1", x"d4", x"e2", x"ea", x"e9", x"e8", x"e8", x"e9", x"e8", x"e6", x"e8", x"e9", 
        x"da", x"d5", x"da", x"e9", x"ed", x"d3", x"ae", x"cc", x"e4", x"e3", x"e0", x"c0", x"b7", x"d0", x"e1", 
        x"e1", x"e2", x"db", x"e0", x"e2", x"d7", x"dc", x"e0", x"de", x"cb", x"cb", x"de", x"df", x"e1", x"d1", 
        x"c7", x"d3", x"df", x"dd", x"d3", x"d9", x"e2", x"dc", x"d8", x"e0", x"df", x"cb", x"c1", x"de", x"e1", 
        x"d9", x"dc", x"de", x"e2", x"e7", x"dd", x"c4", x"d8", x"d0", x"53", x"42", x"88", x"ce", x"ca", x"cc", 
        x"d1", x"bc", x"86", x"7a", x"75", x"67", x"76", x"76", x"6e", x"6b", x"6f", x"70", x"63", x"6c", x"69", 
        x"69", x"63", x"67", x"6b", x"66", x"57", x"5b", x"64", x"5f", x"5d", x"5d", x"5c", x"60", x"4c", x"26", 
        x"39", x"56", x"57", x"4e", x"51", x"5f", x"53", x"4f", x"4e", x"4f", x"5a", x"70", x"74", x"6f", x"3d", 
        x"28", x"34", x"68", x"6f", x"6e", x"74", x"4d", x"40", x"45", x"3e", x"39", x"41", x"42", x"40", x"3e", 
        x"2a", x"22", x"41", x"47", x"30", x"33", x"22", x"1e", x"26", x"2b", x"2d", x"18", x"17", x"13", x"0c", 
        x"12", x"16", x"20", x"2f", x"24", x"14", x"21", x"32", x"35", x"2c", x"28", x"20", x"1d", x"3c", x"73", 
        x"67", x"81", x"8e", x"3e", x"21", x"28", x"25", x"2d", x"3d", x"74", x"a8", x"a9", x"bf", x"cf", x"d4", 
        x"78", x"22", x"27", x"40", x"3b", x"44", x"58", x"5d", x"4d", x"2e", x"26", x"2e", x"2a", x"2a", x"52", 
        x"64", x"59", x"64", x"5d", x"5b", x"66", x"66", x"69", x"61", x"32", x"1b", x"29", x"40", x"44", x"24", 
        x"2a", x"28", x"28", x"60", x"a6", x"7d", x"5a", x"3c", x"41", x"87", x"65", x"2c", x"47", x"76", x"53", 
        x"6d", x"7c", x"46", x"2c", x"46", x"a1", x"a5", x"a4", x"a5", x"a1", x"b3", x"de", x"df", x"e0", x"e0", 
        x"e5", x"e5", x"dc", x"db", x"de", x"d6", x"e1", x"dc", x"e3", x"e0", x"de", x"e1", x"de", x"df", x"df", 
        x"df", x"dd", x"dd", x"e1", x"de", x"e0", x"e0", x"dc", x"e4", x"e2", x"e3", x"de", x"de", x"e4", x"e1", 
        x"e7", x"e1", x"dd", x"e0", x"d9", x"e4", x"e2", x"e0", x"df", x"df", x"e1", x"e3", x"e1", x"df", x"df", 
        x"df", x"e4", x"e2", x"df", x"e1", x"e3", x"e3", x"e2", x"e3", x"e3", x"e2", x"e0", x"e1", x"e0", x"e1", 
        x"e2", x"e2", x"e3", x"e2", x"e3", x"e2", x"e0", x"e1", x"e2", x"e3", x"e1", x"de", x"d2", x"db", x"e5", 
        x"e6", x"e1", x"e1", x"e3", x"e3", x"e2", x"e3", x"de", x"dd", x"db", x"e2", x"e1", x"e4", x"e3", x"e0", 
        x"d8", x"dd", x"e1", x"e3", x"df", x"e3", x"e3", x"e2", x"e1", x"e2", x"e0", x"e0", x"e0", x"e1", x"e1", 
        x"e1", x"e1", x"e0", x"e1", x"e1", x"e1", x"df", x"de", x"de", x"e0", x"e1", x"e0", x"dd", x"e3", x"e0", 
        x"e0", x"e1", x"e1", x"e1", x"e1", x"e1", x"e1", x"e2", x"e3", x"e2", x"e1", x"e0", x"df", x"e0", x"e2", 
        x"e0", x"e0", x"df", x"df", x"e0", x"e0", x"de", x"dd", x"e0", x"df", x"de", x"e2", x"e1", x"e2", x"e2", 
        x"e3", x"e5", x"e2", x"e1", x"e3", x"e4", x"e3", x"e3", x"e4", x"e3", x"e3", x"e4", x"e2", x"e2", x"e0", 
        x"e1", x"e2", x"e3", x"e2", x"e3", x"e3", x"e4", x"e1", x"e1", x"e2", x"e1", x"e0", x"e2", x"e3", x"e4", 
        x"e1", x"e2", x"e4", x"e3", x"e1", x"e1", x"e0", x"e0", x"e0", x"e0", x"e3", x"e3", x"e2", x"e2", x"e1", 
        x"e2", x"e2", x"e1", x"e1", x"e3", x"e4", x"e7", x"e4", x"e3", x"e3", x"e3", x"e4", x"e5", x"e5", x"e4", 
        x"e5", x"e3", x"e2", x"e5", x"e5", x"e2", x"e4", x"e3", x"e2", x"e4", x"e5", x"e5", x"e6", x"e5", x"e6", 
        x"e6", x"d2", x"cd", x"e2", x"e2", x"e2", x"e3", x"e6", x"e4", x"e3", x"e7", x"e5", x"e5", x"e3", x"e3", 
        x"e5", x"e3", x"e2", x"e3", x"e6", x"e1", x"df", x"e2", x"e7", x"e2", x"e2", x"e3", x"e4", x"e3", x"e2", 
        x"e2", x"e2", x"e2", x"e7", x"e8", x"e6", x"e4", x"e4", x"e3", x"e6", x"e5", x"e4", x"e5", x"e5", x"e5", 
        x"e5", x"e5", x"e2", x"e3", x"e4", x"e7", x"e7", x"e6", x"e5", x"e3", x"e3", x"e5", x"e3", x"e6", x"e6", 
        x"e5", x"e3", x"e4", x"e5", x"e6", x"e4", x"e6", x"e6", x"e3", x"e5", x"e7", x"e4", x"e3", x"e5", x"e5", 
        x"e6", x"e7", x"e5", x"e5", x"e6", x"e7", x"e6", x"e8", x"e7", x"e7", x"e8", x"e7", x"e8", x"e4", x"e6", 
        x"e5", x"e4", x"e4", x"e2", x"e6", x"e7", x"e4", x"e5", x"e5", x"e3", x"e3", x"e7", x"e4", x"e3", x"e5", 
        x"e9", x"e6", x"e4", x"e7", x"e6", x"e4", x"e5", x"e4", x"e1", x"e2", x"e7", x"e6", x"e2", x"e4", x"e5", 
        x"e3", x"e2", x"e7", x"e5", x"e5", x"e6", x"e6", x"e3", x"e6", x"e6", x"e4", x"e5", x"e5", x"e2", x"e2", 
        x"e4", x"e6", x"e6", x"e6", x"e7", x"df", x"dd", x"e2", x"e2", x"e2", x"e2", x"e1", x"df", x"df", x"df", 
        x"e0", x"e0", x"e0", x"df", x"df", x"e1", x"e0", x"df", x"de", x"e0", x"e0", x"e0", x"e1", x"e1", x"e0", 
        x"df", x"e1", x"e0", x"e1", x"e2", x"e0", x"e2", x"e4", x"e5", x"e6", x"e9", x"ea", x"e7", x"e4", x"e2", 
        x"e2", x"e8", x"e5", x"c3", x"d8", x"e6", x"e8", x"e5", x"e7", x"e8", x"e4", x"e3", x"e3", x"e3", x"e5", 
        x"e4", x"e5", x"e4", x"e2", x"e2", x"e5", x"e6", x"e6", x"e4", x"e6", x"e6", x"e2", x"e6", x"e6", x"e5", 
        x"e6", x"e4", x"e3", x"e5", x"e4", x"e3", x"e3", x"e3", x"e5", x"e3", x"e4", x"e5", x"e5", x"e5", x"e4", 
        x"e4", x"e3", x"e7", x"eb", x"f0", x"f1", x"eb", x"e4", x"e7", x"e8", x"e4", x"e5", x"e4", x"e3", x"e2", 
        x"e2", x"e4", x"e4", x"e4", x"e2", x"e2", x"e4", x"e5", x"e4", x"e0", x"e1", x"de", x"e1", x"e4", x"e1", 
        x"e4", x"e4", x"e7", x"e8", x"e9", x"e8", x"e7", x"e8", x"e8", x"e9", x"e7", x"e7", x"e7", x"e9", x"e9", 
        x"e6", x"e8", x"e8", x"ea", x"ec", x"da", x"d0", x"e5", x"e7", x"e3", x"dc", x"cf", x"d4", x"e3", x"de", 
        x"e0", x"e2", x"de", x"dd", x"de", x"dd", x"de", x"de", x"dc", x"e0", x"de", x"df", x"dd", x"dd", x"df", 
        x"e1", x"e1", x"da", x"dd", x"e1", x"dc", x"dc", x"dc", x"dc", x"da", x"de", x"e0", x"dc", x"e1", x"de", 
        x"df", x"e4", x"e3", x"e5", x"e7", x"e5", x"e2", x"eb", x"d2", x"53", x"3d", x"89", x"cc", x"c7", x"cc", 
        x"cd", x"d0", x"a1", x"75", x"75", x"73", x"76", x"73", x"6f", x"6e", x"6d", x"6c", x"6a", x"69", x"67", 
        x"70", x"6e", x"68", x"69", x"6a", x"6b", x"66", x"62", x"5f", x"62", x"5e", x"5c", x"60", x"51", x"2a", 
        x"34", x"56", x"5c", x"58", x"56", x"5e", x"5d", x"54", x"53", x"4f", x"5b", x"75", x"76", x"6f", x"43", 
        x"30", x"3c", x"71", x"8b", x"8d", x"82", x"57", x"3e", x"42", x"42", x"41", x"43", x"3e", x"40", x"3f", 
        x"2e", x"20", x"3d", x"4e", x"2b", x"2b", x"39", x"30", x"2c", x"2b", x"28", x"13", x"0e", x"08", x"07", 
        x"0f", x"1f", x"17", x"15", x"0c", x"0b", x"1c", x"34", x"36", x"2d", x"2a", x"26", x"22", x"5f", x"ad", 
        x"94", x"4c", x"3d", x"23", x"2d", x"2e", x"2d", x"35", x"48", x"71", x"a6", x"ac", x"c0", x"d3", x"d1", 
        x"6d", x"26", x"38", x"38", x"2a", x"48", x"5e", x"60", x"5c", x"37", x"25", x"23", x"23", x"22", x"4f", 
        x"6b", x"63", x"67", x"6b", x"69", x"68", x"68", x"6b", x"64", x"3e", x"23", x"2a", x"44", x"47", x"24", 
        x"2e", x"3b", x"55", x"88", x"b4", x"6d", x"47", x"36", x"5a", x"63", x"31", x"37", x"65", x"5a", x"40", 
        x"4d", x"62", x"51", x"57", x"57", x"97", x"9b", x"90", x"8a", x"8e", x"9c", x"c7", x"d1", x"d2", x"d6", 
        x"d9", x"da", x"da", x"da", x"de", x"d9", x"da", x"d3", x"db", x"d8", x"d3", x"d0", x"ca", x"c7", x"c6", 
        x"c8", x"c8", x"cb", x"d0", x"ca", x"cd", x"d8", x"d4", x"d8", x"da", x"d9", x"d8", x"d6", x"d6", x"d8", 
        x"de", x"d2", x"cc", x"d5", x"d8", x"d6", x"d3", x"d4", x"d3", x"d6", x"d8", x"d3", x"cf", x"d4", x"da", 
        x"d8", x"d3", x"d4", x"da", x"da", x"da", x"db", x"db", x"db", x"da", x"d8", x"d6", x"d9", x"da", x"da", 
        x"dc", x"de", x"df", x"db", x"da", x"dc", x"e1", x"df", x"da", x"da", x"d8", x"d5", x"d5", x"dd", x"dc", 
        x"dc", x"df", x"e1", x"de", x"d9", x"d4", x"d4", x"cf", x"d2", x"d3", x"da", x"dd", x"e0", x"de", x"da", 
        x"d4", x"d8", x"df", x"e0", x"e1", x"e5", x"e3", x"e3", x"e5", x"e1", x"e1", x"e3", x"e1", x"e1", x"e4", 
        x"e3", x"e2", x"e5", x"e4", x"e6", x"e6", x"e5", x"e6", x"e5", x"e5", x"e5", x"e4", x"e4", x"ea", x"e7", 
        x"e8", x"e9", x"e8", x"e8", x"e8", x"e8", x"e8", x"e8", x"e6", x"e6", x"e6", x"e5", x"e3", x"e2", x"e4", 
        x"e6", x"e7", x"e4", x"e5", x"e7", x"e4", x"e5", x"e4", x"e5", x"e6", x"e5", x"e3", x"e4", x"e5", x"e2", 
        x"e4", x"e6", x"e6", x"e3", x"e4", x"e5", x"e6", x"e4", x"e4", x"e5", x"e6", x"e6", x"e6", x"e6", x"e5", 
        x"e6", x"e6", x"e7", x"e4", x"e4", x"e5", x"e7", x"e6", x"e5", x"e4", x"e2", x"e4", x"e6", x"e7", x"e3", 
        x"e5", x"e7", x"e4", x"e6", x"e5", x"e4", x"e6", x"e6", x"e5", x"e3", x"e4", x"e5", x"e2", x"e5", x"e9", 
        x"e9", x"e6", x"e4", x"e3", x"e4", x"e6", x"eb", x"e7", x"e7", x"e6", x"e6", x"e6", x"e8", x"e8", x"e9", 
        x"eb", x"e7", x"e5", x"e7", x"e7", x"e7", x"e7", x"e7", x"e7", x"e7", x"e7", x"e7", x"e8", x"e8", x"e7", 
        x"e8", x"e7", x"e7", x"e9", x"e8", x"e5", x"e4", x"e8", x"e7", x"e6", x"e9", x"e8", x"eb", x"eb", x"ea", 
        x"ea", x"e7", x"e4", x"e7", x"ec", x"e8", x"e5", x"e8", x"ec", x"e8", x"e8", x"e9", x"ea", x"e9", x"e8", 
        x"e8", x"ea", x"e9", x"ea", x"e9", x"e7", x"e6", x"e6", x"ea", x"ec", x"ea", x"e9", x"e8", x"e8", x"e7", 
        x"e7", x"e8", x"e6", x"e7", x"e9", x"ea", x"e9", x"e9", x"ec", x"ea", x"e9", x"e7", x"e3", x"e7", x"e7", 
        x"e7", x"e7", x"e6", x"e4", x"e8", x"e9", x"ea", x"e8", x"e7", x"e9", x"e9", x"e7", x"e7", x"e9", x"e8", 
        x"e7", x"e6", x"e7", x"e8", x"e9", x"e9", x"e8", x"e9", x"e7", x"e7", x"e7", x"e8", x"ed", x"ea", x"ec", 
        x"eb", x"eb", x"e9", x"e6", x"e9", x"e8", x"e7", x"ea", x"e9", x"e7", x"e9", x"ed", x"e8", x"e8", x"eb", 
        x"ee", x"eb", x"e8", x"ea", x"ea", x"e9", x"ea", x"eb", x"e9", x"e8", x"eb", x"ea", x"e9", x"ea", x"ea", 
        x"e7", x"e7", x"ea", x"e6", x"e8", x"ea", x"e9", x"e9", x"ea", x"e8", x"e9", x"ec", x"ea", x"e9", x"ea", 
        x"eb", x"eb", x"eb", x"ed", x"ef", x"ea", x"ea", x"ed", x"ec", x"e9", x"eb", x"ec", x"eb", x"ec", x"eb", 
        x"e9", x"e9", x"ec", x"eb", x"ea", x"ea", x"ea", x"e7", x"e8", x"eb", x"ea", x"e9", x"eb", x"eb", x"e9", 
        x"e9", x"ea", x"eb", x"eb", x"ec", x"ea", x"eb", x"ed", x"ed", x"ef", x"f2", x"f1", x"ef", x"ea", x"e8", 
        x"e7", x"e8", x"e9", x"e5", x"e9", x"e9", x"e9", x"e7", x"e9", x"ea", x"e7", x"e7", x"e8", x"e8", x"e8", 
        x"e7", x"e6", x"e5", x"e5", x"e6", x"e8", x"e9", x"e9", x"e8", x"eb", x"ed", x"e8", x"eb", x"ea", x"e6", 
        x"e5", x"e5", x"e8", x"ea", x"ea", x"e9", x"e9", x"ea", x"ea", x"e7", x"e8", x"e9", x"e9", x"e9", x"e9", 
        x"ea", x"e9", x"ea", x"ed", x"f1", x"f2", x"ef", x"ea", x"ef", x"ee", x"e9", x"e9", x"e7", x"e8", x"ea", 
        x"e9", x"e8", x"e7", x"e7", x"e7", x"e7", x"e7", x"e8", x"e9", x"e8", x"ea", x"e7", x"e8", x"e8", x"e8", 
        x"ec", x"ea", x"eb", x"ed", x"ed", x"eb", x"ec", x"ed", x"ed", x"eb", x"eb", x"eb", x"ec", x"ed", x"ed", 
        x"ec", x"eb", x"ed", x"f1", x"f4", x"ec", x"e7", x"ea", x"ec", x"ea", x"e8", x"e8", x"e7", x"e9", x"e4", 
        x"e7", x"e7", x"e6", x"e7", x"e8", x"e7", x"e5", x"e5", x"e4", x"e9", x"e5", x"e6", x"e6", x"ea", x"e8", 
        x"e8", x"eb", x"ea", x"ec", x"e9", x"e5", x"e5", x"e6", x"e7", x"e5", x"e8", x"e8", x"e6", x"e9", x"e6", 
        x"e8", x"ee", x"ee", x"ed", x"ed", x"eb", x"eb", x"f1", x"d9", x"60", x"3c", x"88", x"d2", x"d0", x"ce", 
        x"cd", x"d3", x"b8", x"7f", x"7e", x"7d", x"7b", x"77", x"77", x"75", x"75", x"77", x"74", x"70", x"6e", 
        x"75", x"77", x"73", x"72", x"70", x"75", x"73", x"6e", x"6b", x"6e", x"6b", x"68", x"6c", x"5a", x"2b", 
        x"2f", x"59", x"69", x"69", x"65", x"69", x"6a", x"63", x"64", x"63", x"6f", x"88", x"8b", x"7c", x"4e", 
        x"30", x"35", x"74", x"89", x"83", x"7b", x"60", x"53", x"57", x"58", x"54", x"54", x"54", x"54", x"50", 
        x"37", x"25", x"3a", x"4c", x"2d", x"2b", x"40", x"38", x"2c", x"2e", x"2b", x"13", x"07", x"04", x"06", 
        x"19", x"4e", x"30", x"1a", x"0a", x"0b", x"1d", x"33", x"35", x"35", x"2b", x"21", x"1a", x"28", x"65", 
        x"82", x"43", x"13", x"11", x"25", x"38", x"3b", x"3c", x"4b", x"74", x"af", x"b3", x"c0", x"d3", x"db", 
        x"73", x"29", x"3f", x"2c", x"2a", x"51", x"60", x"5c", x"58", x"43", x"34", x"34", x"2d", x"29", x"58", 
        x"76", x"73", x"6f", x"71", x"6f", x"6a", x"69", x"6a", x"5e", x"40", x"2a", x"30", x"4b", x"4a", x"27", 
        x"3a", x"67", x"75", x"77", x"a0", x"54", x"29", x"3b", x"67", x"72", x"69", x"69", x"48", x"2d", x"2c", 
        x"36", x"49", x"3c", x"84", x"b5", x"c1", x"c6", x"c5", x"c5", x"c5", x"cb", x"dd", x"d8", x"da", x"db", 
        x"dc", x"dc", x"de", x"dc", x"df", x"e1", x"df", x"da", x"de", x"e0", x"df", x"dd", x"db", x"d6", x"d8", 
        x"df", x"e0", x"e0", x"da", x"cd", x"c9", x"d9", x"dc", x"d5", x"d5", x"d8", x"da", x"da", x"d8", x"df", 
        x"e0", x"da", x"de", x"e4", x"e5", x"df", x"dd", x"e2", x"e2", x"e4", x"e6", x"df", x"e1", x"e4", x"e6", 
        x"e1", x"d4", x"d7", x"e3", x"e4", x"e4", x"e4", x"e3", x"e2", x"e2", x"e3", x"e4", x"e1", x"e2", x"e5", 
        x"e5", x"e5", x"e8", x"e8", x"e4", x"e5", x"e7", x"e4", x"e1", x"e6", x"e3", x"e0", x"e4", x"e5", x"e4", 
        x"e2", x"e4", x"e7", x"e5", x"e1", x"e2", x"e2", x"de", x"df", x"e2", x"e4", x"ea", x"e8", x"e5", x"e3", 
        x"e0", x"e0", x"e7", x"e4", x"e7", x"ea", x"e3", x"e4", x"e6", x"e3", x"e3", x"e6", x"e4", x"e1", x"e4", 
        x"e1", x"e2", x"e6", x"de", x"de", x"e2", x"e5", x"e7", x"e5", x"e6", x"e7", x"e5", x"e7", x"ec", x"e9", 
        x"ec", x"eb", x"eb", x"ec", x"ec", x"ec", x"eb", x"eb", x"e8", x"e7", x"e7", x"e8", x"e6", x"e5", x"e8", 
        x"ec", x"eb", x"e7", x"e8", x"eb", x"e8", x"e9", x"eb", x"e8", x"ec", x"ed", x"e8", x"eb", x"eb", x"e5", 
        x"e5", x"ea", x"ed", x"e8", x"e2", x"e3", x"e9", x"ec", x"eb", x"e9", x"e9", x"e9", x"ea", x"ec", x"ef", 
        x"ec", x"ea", x"ed", x"eb", x"ea", x"e7", x"ec", x"ef", x"eb", x"e5", x"e3", x"e5", x"e8", x"ec", x"e8", 
        x"ea", x"eb", x"e4", x"e5", x"e3", x"e5", x"ea", x"ea", x"ec", x"e8", x"e5", x"e6", x"e6", x"e7", x"e7", 
        x"e8", x"e9", x"ec", x"e9", x"e4", x"ea", x"ef", x"ec", x"ec", x"ec", x"eb", x"ea", x"e7", x"ea", x"ed", 
        x"f1", x"ef", x"ed", x"ee", x"e9", x"eb", x"ed", x"ed", x"ec", x"ec", x"ee", x"ee", x"ec", x"ec", x"ec", 
        x"eb", x"f2", x"f2", x"ee", x"ed", x"eb", x"ec", x"ef", x"ec", x"e9", x"ec", x"ed", x"ef", x"f0", x"ee", 
        x"ee", x"eb", x"e9", x"ea", x"ed", x"ec", x"eb", x"eb", x"ec", x"ea", x"ea", x"ec", x"ef", x"f0", x"f0", 
        x"ee", x"ee", x"f0", x"ee", x"ec", x"ec", x"e8", x"e8", x"ed", x"f0", x"ef", x"ee", x"ed", x"ed", x"ed", 
        x"ed", x"eb", x"e4", x"e7", x"ee", x"ef", x"ee", x"ec", x"ee", x"eb", x"eb", x"ea", x"e8", x"ea", x"eb", 
        x"ea", x"ea", x"e9", x"e9", x"ed", x"ef", x"ef", x"eb", x"e9", x"ec", x"ec", x"e9", x"e8", x"eb", x"eb", 
        x"e7", x"e7", x"e9", x"eb", x"eb", x"ea", x"ea", x"eb", x"ea", x"ea", x"ea", x"eb", x"ef", x"ed", x"f0", 
        x"f2", x"f1", x"ee", x"ec", x"ee", x"eb", x"eb", x"ef", x"ec", x"ec", x"ee", x"f0", x"ec", x"ed", x"ed", 
        x"ee", x"ea", x"e9", x"ed", x"ee", x"ee", x"ed", x"ed", x"ed", x"ec", x"ea", x"e9", x"ea", x"ec", x"ec", 
        x"e8", x"e7", x"ee", x"eb", x"ed", x"ed", x"ed", x"ed", x"ec", x"ea", x"ee", x"f2", x"ef", x"eb", x"ec", 
        x"ec", x"ec", x"ec", x"ed", x"ef", x"ed", x"ec", x"ef", x"ed", x"ea", x"ec", x"ed", x"f0", x"f0", x"ed", 
        x"eb", x"ed", x"ef", x"ee", x"ed", x"ee", x"ed", x"ec", x"ed", x"ee", x"ec", x"eb", x"ef", x"f0", x"ed", 
        x"ec", x"ee", x"ee", x"ee", x"ef", x"ed", x"ed", x"ef", x"ef", x"f1", x"f4", x"f1", x"ee", x"eb", x"e9", 
        x"e9", x"eb", x"ec", x"e4", x"e0", x"e6", x"ea", x"ec", x"ec", x"eb", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ed", x"eb", x"eb", x"ed", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ee", x"ec", x"ed", x"ed", x"ed", 
        x"ed", x"ea", x"eb", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f3", x"f1", x"f0", x"f1", x"f3", x"f4", x"f3", x"f1", x"f2", x"f0", x"ed", x"ed", x"ea", x"eb", x"ee", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"e8", x"eb", x"f0", x"ee", x"ee", x"f0", x"f2", 
        x"f0", x"ed", x"ee", x"f0", x"f1", x"f0", x"f0", x"f1", x"ef", x"ee", x"ef", x"f1", x"f2", x"f0", x"ef", 
        x"ef", x"ee", x"ee", x"f0", x"ef", x"ed", x"ee", x"ee", x"ee", x"f0", x"f3", x"f1", x"ed", x"ec", x"e7", 
        x"ea", x"ec", x"ec", x"ee", x"ee", x"ed", x"ec", x"ea", x"e8", x"ea", x"e8", x"ea", x"ec", x"f2", x"f1", 
        x"ef", x"ef", x"ec", x"ec", x"ed", x"eb", x"eb", x"ef", x"ef", x"ed", x"ef", x"ec", x"eb", x"ed", x"ea", 
        x"eb", x"f3", x"f4", x"f0", x"ef", x"f1", x"f0", x"f3", x"e5", x"78", x"3d", x"84", x"da", x"db", x"d3", 
        x"d4", x"d7", x"d3", x"92", x"80", x"80", x"81", x"7d", x"7f", x"7c", x"7d", x"7f", x"7b", x"79", x"74", 
        x"73", x"76", x"75", x"72", x"6e", x"71", x"73", x"6f", x"6a", x"6a", x"6a", x"6b", x"6d", x"5b", x"2a", 
        x"2a", x"56", x"66", x"5c", x"5a", x"5e", x"60", x"5a", x"5a", x"59", x"55", x"4d", x"4b", x"47", x"3a", 
        x"2a", x"2b", x"3f", x"3d", x"3a", x"4a", x"4d", x"50", x"54", x"4f", x"4b", x"4d", x"49", x"46", x"45", 
        x"33", x"20", x"2f", x"57", x"4c", x"4a", x"58", x"58", x"4a", x"4a", x"41", x"1b", x"03", x"01", x"04", 
        x"0f", x"2f", x"1e", x"1e", x"0e", x"06", x"14", x"2a", x"38", x"2f", x"24", x"26", x"2b", x"25", x"6a", 
        x"95", x"5a", x"0f", x"0b", x"23", x"34", x"3e", x"46", x"4d", x"6e", x"ac", x"b2", x"be", x"d8", x"ca", 
        x"4d", x"1a", x"2f", x"1c", x"29", x"4f", x"5c", x"58", x"56", x"3d", x"30", x"3b", x"36", x"36", x"44", 
        x"4a", x"42", x"40", x"3f", x"3f", x"3e", x"32", x"31", x"30", x"30", x"31", x"33", x"3f", x"42", x"28", 
        x"3e", x"36", x"29", x"66", x"ac", x"58", x"57", x"89", x"76", x"5d", x"62", x"53", x"40", x"39", x"2e", 
        x"2d", x"4a", x"74", x"97", x"d8", x"cf", x"db", x"dc", x"d2", x"cf", x"cb", x"e1", x"e2", x"db", x"dc", 
        x"df", x"e0", x"dc", x"df", x"e6", x"e5", x"e4", x"e1", x"e2", x"e5", x"e5", x"e0", x"de", x"dd", x"dc", 
        x"e2", x"e7", x"e5", x"e1", x"db", x"d5", x"d5", x"de", x"df", x"da", x"da", x"e1", x"e9", x"e1", x"e1", 
        x"e7", x"e0", x"e3", x"e9", x"e5", x"e3", x"e3", x"e6", x"e6", x"e6", x"e7", x"e6", x"e7", x"e6", x"e8", 
        x"eb", x"e2", x"e1", x"e3", x"e6", x"e9", x"e6", x"e1", x"e1", x"e5", x"e6", x"e6", x"e2", x"e0", x"e2", 
        x"e4", x"e5", x"e2", x"e3", x"e0", x"e1", x"e5", x"e3", x"df", x"e2", x"e7", x"e7", x"e6", x"e7", x"e5", 
        x"e3", x"e4", x"e2", x"e3", x"e1", x"e6", x"e7", x"e3", x"df", x"e2", x"e6", x"ea", x"e6", x"e9", x"eb", 
        x"ea", x"e6", x"e7", x"e2", x"e3", x"e8", x"e6", x"e4", x"e6", x"e6", x"e1", x"df", x"de", x"df", x"e5", 
        x"e6", x"e1", x"e1", x"e1", x"e4", x"e5", x"e4", x"e9", x"ea", x"e6", x"e7", x"e5", x"e7", x"e9", x"e8", 
        x"e9", x"e4", x"e5", x"e6", x"e7", x"e8", x"e7", x"e7", x"e9", x"e7", x"e8", x"e8", x"e7", x"e7", x"eb", 
        x"ec", x"e8", x"e6", x"e6", x"e8", x"e5", x"e7", x"e9", x"e7", x"ea", x"ea", x"e9", x"eb", x"e8", x"e5", 
        x"e4", x"e7", x"ea", x"e5", x"df", x"e2", x"eb", x"eb", x"e8", x"e4", x"e3", x"e4", x"e6", x"e8", x"eb", 
        x"e9", x"e8", x"e8", x"e5", x"e8", x"e7", x"e7", x"ea", x"e7", x"e1", x"e1", x"e6", x"e8", x"e9", x"e8", 
        x"e8", x"e8", x"e7", x"e8", x"e7", x"e8", x"e8", x"e8", x"ee", x"eb", x"e7", x"e9", x"ea", x"e7", x"e3", 
        x"e4", x"e7", x"ea", x"e8", x"e4", x"ea", x"ee", x"ea", x"ea", x"ec", x"ea", x"e9", x"e7", x"ea", x"eb", 
        x"ee", x"eb", x"ea", x"ea", x"e5", x"e7", x"eb", x"eb", x"e9", x"e9", x"ed", x"ed", x"ec", x"eb", x"ed", 
        x"eb", x"ea", x"ec", x"ed", x"eb", x"eb", x"ec", x"eb", x"e9", x"e9", x"ed", x"ee", x"ec", x"ea", x"e8", 
        x"eb", x"ea", x"ec", x"ec", x"ef", x"ee", x"ee", x"eb", x"ed", x"ec", x"e9", x"e9", x"eb", x"eb", x"eb", 
        x"ea", x"e9", x"e9", x"e6", x"e9", x"ea", x"e8", x"eb", x"ee", x"ee", x"ee", x"ed", x"ec", x"ec", x"ee", 
        x"ef", x"eb", x"dd", x"e0", x"e8", x"ea", x"ea", x"e7", x"e9", x"ea", x"ea", x"ea", x"e9", x"e7", x"e5", 
        x"e4", x"e8", x"ea", x"e9", x"eb", x"ec", x"ed", x"ed", x"ea", x"ec", x"ed", x"ea", x"e9", x"eb", x"ec", 
        x"e9", x"ea", x"eb", x"ed", x"ec", x"ea", x"eb", x"eb", x"ec", x"ee", x"ee", x"ee", x"ec", x"eb", x"ed", 
        x"ed", x"ed", x"ec", x"ea", x"ea", x"e7", x"e7", x"ed", x"e9", x"ea", x"eb", x"eb", x"e9", x"eb", x"ec", 
        x"ec", x"e9", x"e9", x"ed", x"ec", x"ec", x"ed", x"ec", x"ec", x"ea", x"e9", x"e8", x"e8", x"e8", x"e9", 
        x"e5", x"e2", x"ec", x"ed", x"ef", x"ef", x"ed", x"ee", x"ed", x"ec", x"ee", x"ef", x"f0", x"f0", x"ef", 
        x"ee", x"ed", x"ee", x"ef", x"f0", x"ed", x"ec", x"ef", x"ee", x"ec", x"ee", x"ee", x"ef", x"ef", x"ec", 
        x"ec", x"ef", x"f0", x"ee", x"ed", x"ef", x"ef", x"ee", x"ee", x"f0", x"ed", x"e9", x"eb", x"ef", x"ee", 
        x"ec", x"ef", x"ef", x"ed", x"f0", x"ee", x"ef", x"f1", x"f2", x"f4", x"f7", x"f7", x"f5", x"f1", x"ee", 
        x"ec", x"ed", x"ed", x"e6", x"e5", x"f3", x"f3", x"f3", x"f2", x"ef", x"f1", x"f2", x"f3", x"f3", x"f2", 
        x"f1", x"ef", x"ee", x"ee", x"ef", x"ee", x"ec", x"ec", x"ed", x"ed", x"ec", x"ec", x"ec", x"ed", x"f0", 
        x"f0", x"ee", x"ec", x"ed", x"ef", x"ef", x"f0", x"f0", x"ef", x"ed", x"ef", x"f1", x"f1", x"ef", x"f0", 
        x"f3", x"f2", x"f2", x"f3", x"f3", x"f3", x"f1", x"f0", x"ef", x"ee", x"ef", x"ef", x"ea", x"eb", x"ee", 
        x"ee", x"ef", x"ee", x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ef", x"f0", x"ef", x"f0", x"f0", x"f1", 
        x"f0", x"ed", x"ee", x"f0", x"f2", x"f0", x"f1", x"f0", x"ef", x"f0", x"f0", x"f1", x"f1", x"f0", x"ea", 
        x"eb", x"ed", x"ed", x"f2", x"f2", x"f0", x"f0", x"ed", x"f0", x"f2", x"f0", x"ee", x"eb", x"ea", x"e5", 
        x"e9", x"ec", x"ec", x"ee", x"ee", x"ec", x"eb", x"ec", x"eb", x"ec", x"eb", x"eb", x"eb", x"ed", x"ed", 
        x"ec", x"ec", x"eb", x"ec", x"ed", x"ed", x"ec", x"f1", x"ee", x"ed", x"ef", x"ee", x"eb", x"ec", x"ec", 
        x"ec", x"f2", x"f2", x"ef", x"ef", x"f1", x"f0", x"f2", x"eb", x"8e", x"3c", x"7d", x"d7", x"d8", x"d2", 
        x"d6", x"d4", x"da", x"98", x"82", x"86", x"81", x"80", x"7e", x"7e", x"7c", x"7b", x"77", x"79", x"75", 
        x"71", x"74", x"72", x"6f", x"6c", x"6d", x"6f", x"6b", x"68", x"65", x"64", x"65", x"63", x"58", x"2c", 
        x"28", x"4e", x"60", x"5c", x"59", x"5b", x"5d", x"5a", x"5a", x"59", x"45", x"2c", x"2b", x"2b", x"2e", 
        x"2f", x"3f", x"48", x"3a", x"3b", x"4e", x"53", x"55", x"56", x"50", x"5a", x"5c", x"4b", x"3d", x"39", 
        x"2e", x"23", x"2f", x"53", x"40", x"37", x"3d", x"44", x"3c", x"3b", x"32", x"12", x"01", x"01", x"05", 
        x"10", x"22", x"18", x"23", x"13", x"04", x"0a", x"1d", x"33", x"20", x"1b", x"27", x"2a", x"21", x"57", 
        x"9e", x"72", x"14", x"0d", x"2d", x"3c", x"42", x"50", x"53", x"69", x"a9", x"b2", x"c0", x"d5", x"98", 
        x"1f", x"14", x"20", x"16", x"24", x"4f", x"5c", x"59", x"5b", x"44", x"27", x"32", x"38", x"3a", x"3f", 
        x"3a", x"38", x"3c", x"44", x"45", x"40", x"3b", x"3d", x"3c", x"40", x"40", x"3c", x"3e", x"39", x"25", 
        x"44", x"3c", x"23", x"74", x"c0", x"66", x"78", x"7a", x"34", x"3a", x"55", x"45", x"4b", x"42", x"44", 
        x"45", x"54", x"6d", x"8e", x"da", x"c6", x"cf", x"da", x"ce", x"ce", x"d1", x"e3", x"e5", x"e3", x"df", 
        x"e2", x"e4", x"de", x"e2", x"e4", x"e0", x"e8", x"e5", x"e0", x"e2", x"e2", x"e1", x"e1", x"e5", x"df", 
        x"de", x"de", x"dc", x"de", x"e5", x"e4", x"e4", x"e6", x"df", x"de", x"e4", x"e8", x"ea", x"e4", x"e1", 
        x"e2", x"e2", x"e4", x"e5", x"de", x"e3", x"e5", x"e2", x"e3", x"e3", x"e1", x"e7", x"e7", x"e5", x"e5", 
        x"e8", x"e6", x"e7", x"e7", x"e8", x"e8", x"e2", x"df", x"e4", x"e7", x"e2", x"e7", x"e9", x"e6", x"e0", 
        x"e2", x"e7", x"df", x"e2", x"e5", x"e5", x"e3", x"e4", x"e6", x"e6", x"e8", x"e9", x"e8", x"e6", x"e7", 
        x"e3", x"e2", x"e1", x"e2", x"df", x"e4", x"e6", x"e7", x"e4", x"e8", x"e8", x"e8", x"e3", x"ea", x"ed", 
        x"eb", x"e6", x"e7", x"e5", x"e2", x"e5", x"e8", x"e3", x"e4", x"ed", x"e8", x"e0", x"dd", x"df", x"e4", 
        x"e6", x"e5", x"e5", x"e7", x"e9", x"e6", x"e2", x"eb", x"ee", x"e9", x"e8", x"e7", x"e8", x"e6", x"e7", 
        x"e7", x"e4", x"e5", x"e6", x"e7", x"e8", x"e9", x"e9", x"ea", x"e9", x"ea", x"e9", x"e7", x"e6", x"e8", 
        x"ea", x"e8", x"e8", x"e7", x"e8", x"e4", x"e8", x"eb", x"e9", x"ea", x"e5", x"e9", x"e9", x"e4", x"e6", 
        x"e5", x"e7", x"eb", x"e9", x"e4", x"e8", x"ee", x"e8", x"e8", x"e7", x"e8", x"e9", x"ea", x"eb", x"ea", 
        x"e9", x"e7", x"e3", x"e0", x"e7", x"e7", x"e6", x"eb", x"e9", x"e3", x"e4", x"e8", x"e8", x"e9", x"e7", 
        x"e7", x"e8", x"e5", x"e9", x"ea", x"e9", x"e7", x"e6", x"ec", x"ea", x"e7", x"e9", x"ed", x"eb", x"ea", 
        x"ed", x"ea", x"e8", x"eb", x"ea", x"ec", x"ed", x"e9", x"e8", x"ec", x"ea", x"ea", x"e8", x"eb", x"eb", 
        x"ed", x"eb", x"ec", x"ed", x"ea", x"e9", x"ea", x"eb", x"eb", x"ea", x"e9", x"eb", x"ed", x"ee", x"ef", 
        x"ee", x"e9", x"ec", x"ef", x"ed", x"ec", x"ed", x"ea", x"e9", x"ee", x"f1", x"ee", x"ec", x"eb", x"e9", 
        x"eb", x"ec", x"ef", x"ed", x"ee", x"ec", x"ed", x"ec", x"ed", x"ee", x"ef", x"ed", x"ea", x"e9", x"e9", 
        x"eb", x"ec", x"eb", x"e9", x"ec", x"ec", x"eb", x"ee", x"ef", x"ed", x"ee", x"ed", x"ed", x"ec", x"ed", 
        x"ee", x"ec", x"e1", x"e2", x"ea", x"ea", x"ec", x"ea", x"ea", x"eb", x"ea", x"e9", x"ea", x"e8", x"e8", 
        x"ea", x"ed", x"ec", x"ea", x"eb", x"ee", x"ef", x"ee", x"eb", x"ec", x"ec", x"ea", x"ea", x"ec", x"eb", 
        x"ea", x"ed", x"ec", x"ee", x"ed", x"ea", x"ec", x"ea", x"eb", x"ed", x"ed", x"eb", x"e9", x"ec", x"ee", 
        x"ee", x"ed", x"ef", x"ef", x"ef", x"ea", x"ea", x"ef", x"ec", x"ed", x"ec", x"ed", x"ed", x"ee", x"ee", 
        x"ee", x"ec", x"ec", x"ed", x"ea", x"ea", x"ed", x"ec", x"ea", x"eb", x"ea", x"eb", x"ea", x"e8", x"e9", 
        x"e5", x"df", x"eb", x"ec", x"ef", x"ef", x"ee", x"ef", x"ef", x"f0", x"ed", x"ec", x"f0", x"f0", x"ef", 
        x"ec", x"ec", x"ed", x"ef", x"f0", x"ec", x"eb", x"ef", x"f1", x"ef", x"f1", x"f0", x"ee", x"ed", x"ec", 
        x"ee", x"f0", x"f0", x"ee", x"ed", x"ef", x"ef", x"ee", x"ef", x"f1", x"ee", x"ea", x"ea", x"ef", x"ef", 
        x"ed", x"f1", x"f1", x"ef", x"ef", x"ed", x"ef", x"f2", x"f3", x"f5", x"f8", x"f7", x"f5", x"f1", x"f0", 
        x"ef", x"f0", x"f0", x"e8", x"e5", x"f2", x"ef", x"ed", x"f0", x"ee", x"f0", x"f0", x"f1", x"f2", x"f2", 
        x"f1", x"ef", x"f0", x"f0", x"f1", x"f0", x"ee", x"ed", x"ef", x"ef", x"f0", x"f1", x"ed", x"ee", x"f1", 
        x"f0", x"ee", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"f2", x"ef", x"f2", x"f4", x"f4", x"f1", x"f2", 
        x"f4", x"f2", x"f2", x"f3", x"f4", x"f2", x"f0", x"ee", x"ed", x"ee", x"f0", x"ee", x"e9", x"ea", x"ef", 
        x"f0", x"f2", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", x"ed", x"ee", x"f2", x"f0", x"f0", 
        x"f0", x"ed", x"f0", x"f1", x"f1", x"ef", x"f0", x"f0", x"f0", x"f1", x"f0", x"ef", x"f1", x"f4", x"ef", 
        x"f1", x"f2", x"ef", x"f2", x"f2", x"ef", x"ee", x"ed", x"f0", x"f0", x"ee", x"f0", x"ef", x"eb", x"e4", 
        x"e9", x"eb", x"ed", x"ee", x"ef", x"ef", x"ed", x"ee", x"f0", x"ee", x"ef", x"ec", x"ea", x"e9", x"eb", 
        x"eb", x"ea", x"ee", x"ee", x"eb", x"ed", x"ed", x"ee", x"ea", x"eb", x"ed", x"eb", x"eb", x"ef", x"f0", 
        x"ef", x"f3", x"f2", x"f1", x"f1", x"f0", x"ee", x"f0", x"ec", x"9a", x"39", x"73", x"d6", x"d8", x"d6", 
        x"d9", x"d4", x"da", x"99", x"91", x"97", x"7f", x"80", x"7b", x"7d", x"7d", x"7a", x"79", x"7c", x"79", 
        x"75", x"75", x"70", x"6e", x"6d", x"6d", x"6d", x"6b", x"6d", x"68", x"65", x"65", x"62", x"5c", x"30", 
        x"26", x"49", x"5f", x"5e", x"5b", x"59", x"59", x"5a", x"5a", x"5c", x"4f", x"34", x"34", x"32", x"31", 
        x"2d", x"3f", x"4c", x"38", x"3b", x"4e", x"53", x"53", x"54", x"54", x"60", x"5f", x"51", x"45", x"3b", 
        x"2b", x"22", x"2f", x"4f", x"3d", x"36", x"39", x"3c", x"3a", x"3c", x"2a", x"0c", x"02", x"03", x"09", 
        x"18", x"22", x"18", x"23", x"15", x"07", x"03", x"0e", x"1d", x"26", x"32", x"37", x"30", x"21", x"31", 
        x"89", x"91", x"36", x"0d", x"1b", x"3d", x"44", x"49", x"52", x"65", x"a6", x"af", x"c1", x"cf", x"74", 
        x"12", x"18", x"21", x"18", x"2a", x"56", x"5c", x"59", x"59", x"52", x"31", x"30", x"42", x"41", x"44", 
        x"44", x"42", x"40", x"43", x"40", x"37", x"36", x"3c", x"39", x"3a", x"37", x"37", x"3c", x"36", x"23", 
        x"53", x"45", x"2a", x"7a", x"c4", x"58", x"4b", x"5e", x"61", x"78", x"4e", x"27", x"23", x"51", x"87", 
        x"80", x"53", x"2e", x"80", x"dd", x"c6", x"cb", x"e0", x"ca", x"c7", x"ce", x"e0", x"e3", x"e5", x"e0", 
        x"db", x"db", x"dc", x"dd", x"db", x"e3", x"e4", x"e1", x"de", x"e1", x"e1", x"e2", x"df", x"e0", x"dc", 
        x"e0", x"e3", x"e1", x"e3", x"e6", x"de", x"e3", x"e7", x"e0", x"e4", x"e6", x"e4", x"e8", x"e8", x"e1", 
        x"dc", x"e5", x"e6", x"df", x"dc", x"e3", x"e5", x"df", x"e2", x"e2", x"e0", x"e6", x"e5", x"e7", x"e8", 
        x"e8", x"e7", x"e8", x"e9", x"ea", x"e8", x"e2", x"e2", x"e9", x"e9", x"e1", x"e6", x"e7", x"e6", x"e3", 
        x"e0", x"e7", x"e6", x"e5", x"e8", x"e4", x"cc", x"cd", x"e3", x"e9", x"e8", x"e7", x"e6", x"e6", x"e9", 
        x"e6", x"e3", x"dd", x"e1", x"e1", x"e5", x"e9", x"eb", x"e7", x"e7", x"e8", x"e8", x"e4", x"e8", x"eb", 
        x"e9", x"e7", x"e9", x"e7", x"e5", x"e6", x"e9", x"e5", x"e6", x"ea", x"ea", x"e6", x"e3", x"e5", x"e4", 
        x"e4", x"e4", x"e1", x"df", x"e5", x"eb", x"e9", x"ea", x"eb", x"eb", x"ea", x"ea", x"e9", x"e4", x"e9", 
        x"e7", x"e8", x"e8", x"e8", x"e9", x"ea", x"ea", x"eb", x"ea", x"ec", x"eb", x"e7", x"e6", x"e6", x"e5", 
        x"e5", x"e5", x"e8", x"e5", x"e4", x"e1", x"e5", x"eb", x"ea", x"e9", x"e2", x"e6", x"e8", x"e4", x"e9", 
        x"ea", x"ea", x"ec", x"ec", x"e8", x"e9", x"ec", x"e7", x"e8", x"ea", x"eb", x"eb", x"ea", x"e9", x"e6", 
        x"e2", x"e1", x"e1", x"e2", x"e2", x"d6", x"e1", x"e9", x"e8", x"e6", x"e9", x"ed", x"eb", x"ec", x"e7", 
        x"e7", x"e9", x"e4", x"ea", x"ec", x"ea", x"e8", x"e6", x"eb", x"e9", x"e7", x"ea", x"ec", x"e9", x"e6", 
        x"eb", x"e9", x"e8", x"eb", x"e9", x"ec", x"ed", x"ea", x"e9", x"ed", x"ea", x"ea", x"e8", x"ec", x"eb", 
        x"eb", x"ea", x"eb", x"eb", x"ee", x"ed", x"ea", x"ea", x"ec", x"ea", x"e6", x"e7", x"ea", x"ea", x"ea", 
        x"eb", x"eb", x"ed", x"ee", x"ea", x"ea", x"ee", x"ee", x"ec", x"ec", x"ec", x"ee", x"ec", x"ed", x"ed", 
        x"ed", x"eb", x"ed", x"ea", x"eb", x"ea", x"ec", x"ec", x"ed", x"ed", x"ef", x"ee", x"ec", x"ec", x"ed", 
        x"ed", x"ec", x"eb", x"ec", x"ec", x"ea", x"eb", x"ed", x"ed", x"ed", x"ee", x"ee", x"ed", x"ec", x"eb", 
        x"eb", x"e9", x"de", x"e2", x"ee", x"ec", x"ee", x"ea", x"ec", x"ec", x"eb", x"e9", x"eb", x"ea", x"ed", 
        x"ef", x"ee", x"eb", x"ec", x"ed", x"f1", x"ee", x"ea", x"ea", x"eb", x"eb", x"ea", x"eb", x"ed", x"ea", 
        x"e9", x"ed", x"eb", x"ee", x"ed", x"eb", x"ec", x"e9", x"ea", x"e8", x"e9", x"ea", x"ea", x"f0", x"ef", 
        x"ec", x"ea", x"ec", x"ed", x"ec", x"e9", x"ea", x"ed", x"eb", x"ec", x"e7", x"e9", x"ec", x"eb", x"ec", 
        x"ee", x"ed", x"ef", x"ef", x"ec", x"ee", x"ed", x"e9", x"e9", x"eb", x"ea", x"ec", x"ec", x"ea", x"ec", 
        x"e8", x"e0", x"ec", x"ec", x"ef", x"ef", x"ee", x"f0", x"f0", x"f0", x"ed", x"ec", x"f0", x"ee", x"ec", 
        x"eb", x"ec", x"ed", x"ed", x"ed", x"eb", x"ea", x"ee", x"ef", x"ee", x"ef", x"ed", x"ed", x"ec", x"ec", 
        x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"ed", x"ec", x"ed", x"f0", x"ef", x"eb", x"eb", x"ef", x"ee", 
        x"ed", x"ef", x"f2", x"f1", x"ee", x"ed", x"ef", x"f3", x"f3", x"f3", x"f6", x"f4", x"f2", x"f0", x"ef", 
        x"ee", x"ef", x"ee", x"e8", x"e1", x"ed", x"ed", x"ed", x"f2", x"f2", x"ef", x"ef", x"f0", x"f1", x"f1", 
        x"f0", x"ef", x"ef", x"f1", x"f1", x"f1", x"f0", x"f0", x"ef", x"ef", x"f1", x"f2", x"ee", x"ef", x"f2", 
        x"f0", x"ef", x"f1", x"ef", x"ee", x"ef", x"f0", x"f1", x"f1", x"ef", x"f2", x"f5", x"f4", x"f1", x"f0", 
        x"f1", x"f0", x"f1", x"f3", x"f3", x"f1", x"f0", x"ef", x"ee", x"ee", x"ef", x"ec", x"e6", x"ea", x"f0", 
        x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"ee", x"ec", x"ee", x"f1", x"ee", x"ef", 
        x"ef", x"ee", x"f1", x"f0", x"ef", x"ec", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"f1", x"f6", x"f2", 
        x"f1", x"f1", x"f0", x"f0", x"f2", x"f1", x"f2", x"ee", x"eb", x"ef", x"f0", x"f0", x"ef", x"ed", x"e6", 
        x"ec", x"ee", x"ed", x"ed", x"f0", x"f1", x"ef", x"ee", x"ed", x"e8", x"eb", x"eb", x"ec", x"eb", x"e8", 
        x"eb", x"ef", x"f1", x"ea", x"eb", x"ef", x"f1", x"ee", x"ec", x"ef", x"ee", x"ec", x"ed", x"f1", x"ef", 
        x"ef", x"f2", x"f1", x"f2", x"f3", x"f0", x"ef", x"f0", x"ed", x"a4", x"3a", x"6b", x"cf", x"d6", x"d7", 
        x"d9", x"d6", x"d9", x"98", x"97", x"b3", x"82", x"7a", x"7c", x"7e", x"7f", x"7a", x"79", x"7a", x"78", 
        x"78", x"76", x"70", x"70", x"6e", x"6b", x"6b", x"68", x"6c", x"68", x"65", x"66", x"62", x"5e", x"31", 
        x"22", x"47", x"62", x"5e", x"5e", x"5b", x"5b", x"5c", x"58", x"5b", x"57", x"3d", x"39", x"38", x"35", 
        x"2e", x"3b", x"4e", x"34", x"3b", x"4f", x"54", x"52", x"4f", x"4d", x"49", x"3f", x"40", x"40", x"3d", 
        x"2c", x"21", x"2d", x"4c", x"3f", x"36", x"36", x"3b", x"40", x"3e", x"21", x"05", x"04", x"04", x"08", 
        x"1d", x"30", x"1e", x"1e", x"19", x"12", x"05", x"09", x"1a", x"23", x"2d", x"3c", x"2b", x"18", x"21", 
        x"73", x"a4", x"6d", x"18", x"0b", x"39", x"4f", x"4e", x"5d", x"6a", x"a6", x"ac", x"c4", x"ca", x"5e", 
        x"0e", x"17", x"25", x"1a", x"33", x"57", x"55", x"58", x"58", x"5a", x"46", x"32", x"3a", x"3e", x"40", 
        x"3a", x"39", x"3a", x"3b", x"36", x"37", x"39", x"39", x"35", x"36", x"39", x"37", x"31", x"2b", x"1c", 
        x"4b", x"32", x"25", x"6f", x"c9", x"68", x"49", x"52", x"59", x"7b", x"50", x"3e", x"4b", x"6e", x"78", 
        x"6c", x"43", x"25", x"7d", x"dd", x"c3", x"cc", x"e0", x"ca", x"c5", x"cf", x"e4", x"e2", x"df", x"e0", 
        x"db", x"e0", x"e5", x"d3", x"c4", x"e0", x"e1", x"e2", x"e4", x"e9", x"e9", x"ea", x"e3", x"e1", x"e1", 
        x"e5", x"e5", x"e4", x"e2", x"df", x"de", x"e0", x"e7", x"e7", x"e2", x"e4", x"e5", x"e6", x"e5", x"e6", 
        x"e3", x"e4", x"e8", x"e6", x"e8", x"e6", x"e3", x"e2", x"e6", x"e8", x"e6", x"e5", x"e7", x"e4", x"e6", 
        x"e8", x"ea", x"e5", x"e4", x"e9", x"e7", x"e5", x"e5", x"e5", x"e4", x"e5", x"e7", x"e7", x"ea", x"e3", 
        x"db", x"e5", x"ec", x"e6", x"e5", x"e7", x"d4", x"d2", x"e2", x"e5", x"e5", x"e7", x"e7", x"e4", x"e9", 
        x"e8", x"df", x"d8", x"e3", x"e2", x"e4", x"e8", x"ea", x"e7", x"e5", x"e7", x"ec", x"e9", x"e7", x"e8", 
        x"e7", x"e8", x"e9", x"e7", x"ea", x"e7", x"e6", x"e7", x"e8", x"e3", x"e8", x"ea", x"e5", x"e7", x"e6", 
        x"e8", x"ed", x"ec", x"e6", x"e9", x"ea", x"e5", x"e7", x"ea", x"e9", x"e8", x"ea", x"e8", x"e2", x"e9", 
        x"e6", x"e9", x"e8", x"e8", x"e7", x"e7", x"e7", x"e8", x"e9", x"ec", x"e8", x"e2", x"e4", x"ea", x"eb", 
        x"e8", x"ea", x"ef", x"e9", x"e8", x"e6", x"e9", x"ee", x"e6", x"e6", x"e3", x"e3", x"eb", x"eb", x"ec", 
        x"e9", x"e8", x"ea", x"eb", x"e8", x"e7", x"e8", x"ea", x"ea", x"e9", x"e9", x"e9", x"e9", x"e8", x"e8", 
        x"eb", x"eb", x"e6", x"e5", x"e7", x"da", x"e4", x"ea", x"e7", x"e6", x"e9", x"ec", x"ea", x"eb", x"ec", 
        x"ea", x"e9", x"ea", x"e9", x"e8", x"ec", x"ea", x"e6", x"e9", x"e9", x"ea", x"ed", x"ed", x"ea", x"ea", 
        x"eb", x"e4", x"e4", x"ed", x"ec", x"ea", x"ea", x"e9", x"e7", x"ec", x"e8", x"e7", x"e6", x"ea", x"ea", 
        x"e9", x"e8", x"e9", x"e6", x"e9", x"ec", x"ed", x"eb", x"e8", x"e8", x"ea", x"ed", x"e6", x"e3", x"e9", 
        x"ea", x"ed", x"ef", x"ef", x"ec", x"e8", x"ed", x"f0", x"ef", x"ea", x"e7", x"f0", x"ed", x"ee", x"ed", 
        x"ec", x"e9", x"ea", x"ea", x"ed", x"ec", x"ef", x"f0", x"f1", x"ee", x"ec", x"ea", x"e9", x"ea", x"eb", 
        x"ec", x"eb", x"ec", x"ed", x"ec", x"ec", x"ed", x"ea", x"e9", x"ec", x"ee", x"ed", x"ec", x"ed", x"ed", 
        x"ec", x"ea", x"dd", x"e3", x"ef", x"e8", x"e8", x"e8", x"ec", x"eb", x"ea", x"ea", x"ed", x"ec", x"ee", 
        x"f0", x"ec", x"ea", x"eb", x"e8", x"e9", x"e9", x"ea", x"eb", x"ec", x"eb", x"ec", x"ee", x"ee", x"eb", 
        x"e7", x"ea", x"e9", x"ed", x"ee", x"ec", x"ec", x"e9", x"ea", x"e4", x"e7", x"ee", x"f0", x"f1", x"ed", 
        x"ef", x"eb", x"eb", x"eb", x"ec", x"ea", x"ec", x"ee", x"ed", x"ee", x"e8", x"ea", x"ef", x"ec", x"ea", 
        x"ec", x"ec", x"ec", x"ec", x"eb", x"f0", x"ec", x"e7", x"eb", x"ed", x"e9", x"eb", x"ef", x"ec", x"ec", 
        x"e9", x"e0", x"ed", x"ed", x"f1", x"ef", x"ec", x"ef", x"ec", x"ec", x"ec", x"ed", x"f0", x"ec", x"ed", 
        x"ee", x"ef", x"f0", x"ef", x"ed", x"f0", x"ef", x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"ee", x"ec", 
        x"ed", x"ed", x"ec", x"ee", x"ef", x"ee", x"ee", x"ec", x"ee", x"f1", x"f2", x"ee", x"eb", x"ef", x"f1", 
        x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f3", x"f6", x"f5", x"f4", x"f5", x"f4", x"f2", x"f1", x"ef", 
        x"ef", x"f0", x"f0", x"e9", x"e1", x"ed", x"f1", x"ef", x"f0", x"f2", x"f0", x"f1", x"f2", x"f2", x"f1", 
        x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f1", x"f1", x"ee", x"ed", x"ef", x"f0", x"ec", x"ef", x"f1", 
        x"ee", x"f0", x"f2", x"f0", x"ee", x"ee", x"ef", x"f1", x"f1", x"ef", x"f3", x"f7", x"f6", x"f1", x"ef", 
        x"f0", x"ee", x"ee", x"f0", x"f1", x"ef", x"ef", x"f1", x"ee", x"ed", x"ef", x"ed", x"e7", x"ea", x"ef", 
        x"ed", x"ed", x"ed", x"ee", x"ef", x"f0", x"f1", x"f1", x"ee", x"f1", x"f0", x"f0", x"f1", x"ed", x"f0", 
        x"f0", x"f0", x"f3", x"f1", x"ee", x"ec", x"ee", x"ee", x"ed", x"ee", x"ef", x"f1", x"f2", x"f1", x"f0", 
        x"ed", x"f1", x"f3", x"ee", x"ed", x"f0", x"f2", x"ee", x"ec", x"f0", x"f0", x"ef", x"f0", x"f0", x"ec", 
        x"ef", x"f2", x"ef", x"ed", x"ee", x"f0", x"ed", x"ed", x"ee", x"e9", x"ed", x"ea", x"ea", x"eb", x"e9", 
        x"f0", x"d9", x"a0", x"6c", x"82", x"c2", x"eb", x"f0", x"f0", x"ef", x"eb", x"ee", x"f1", x"f1", x"eb", 
        x"eb", x"f1", x"f1", x"f1", x"f1", x"ef", x"ef", x"f2", x"ef", x"ad", x"40", x"6b", x"cf", x"db", x"d8", 
        x"d7", x"d8", x"dc", x"95", x"8a", x"d6", x"98", x"7a", x"81", x"7d", x"79", x"79", x"79", x"77", x"74", 
        x"78", x"77", x"73", x"75", x"72", x"6c", x"6c", x"68", x"69", x"67", x"65", x"64", x"60", x"5e", x"31", 
        x"20", x"45", x"60", x"5b", x"5d", x"5a", x"58", x"5a", x"55", x"58", x"56", x"45", x"3b", x"38", x"33", 
        x"2e", x"39", x"52", x"35", x"39", x"4b", x"4f", x"4b", x"49", x"4e", x"48", x"3d", x"3f", x"3d", x"44", 
        x"36", x"26", x"2a", x"45", x"46", x"42", x"44", x"44", x"49", x"49", x"27", x"0b", x"0b", x"08", x"04", 
        x"14", x"20", x"16", x"17", x"18", x"17", x"07", x"0e", x"1b", x"28", x"33", x"3b", x"2a", x"23", x"1c", 
        x"60", x"96", x"90", x"38", x"06", x"22", x"4c", x"4f", x"5a", x"66", x"a4", x"ab", x"c5", x"ba", x"40", 
        x"0f", x"19", x"25", x"1a", x"39", x"56", x"53", x"5a", x"59", x"5a", x"51", x"31", x"3c", x"43", x"2d", 
        x"18", x"16", x"26", x"3b", x"3c", x"3d", x"38", x"39", x"3b", x"3d", x"3f", x"2d", x"14", x"0c", x"0f", 
        x"38", x"3d", x"35", x"69", x"cd", x"80", x"3f", x"31", x"42", x"6e", x"56", x"3a", x"41", x"5c", x"66", 
        x"72", x"4b", x"2d", x"7a", x"e2", x"c9", x"cf", x"e0", x"cd", x"ca", x"d5", x"e6", x"e0", x"e3", x"e6", 
        x"e0", x"e2", x"e5", x"db", x"ce", x"e1", x"de", x"dd", x"e8", x"e8", x"e7", x"e6", x"e1", x"e4", x"de", 
        x"df", x"e2", x"e5", x"e4", x"e4", x"e1", x"df", x"e3", x"e4", x"e2", x"e3", x"e5", x"e5", x"e2", x"e7", 
        x"e8", x"e6", x"e4", x"e5", x"e7", x"e6", x"e4", x"e5", x"e7", x"ea", x"e7", x"e5", x"e6", x"e6", x"e7", 
        x"e7", x"e6", x"e5", x"e6", x"e9", x"e9", x"e6", x"e3", x"e5", x"e4", x"e6", x"e7", x"e5", x"ea", x"e1", 
        x"e2", x"eb", x"ec", x"e2", x"e1", x"e6", x"e4", x"e3", x"e3", x"e4", x"e7", x"e5", x"e4", x"e3", x"e2", 
        x"e3", x"de", x"da", x"e8", x"de", x"e3", x"eb", x"ea", x"eb", x"ec", x"ea", x"ea", x"e8", x"e7", x"e6", 
        x"e5", x"e7", x"e6", x"e9", x"ea", x"e8", x"e5", x"e5", x"e9", x"e9", x"e5", x"e6", x"ea", x"ea", x"e8", 
        x"e6", x"e6", x"e8", x"e8", x"eb", x"eb", x"e4", x"e4", x"e7", x"eb", x"ea", x"ea", x"e9", x"e4", x"e8", 
        x"e5", x"e3", x"e8", x"e8", x"e4", x"e8", x"e5", x"e8", x"e9", x"e9", x"e7", x"e4", x"e4", x"e6", x"e6", 
        x"e5", x"e8", x"ed", x"e8", x"ea", x"ec", x"ea", x"e8", x"e3", x"e7", x"e8", x"e8", x"eb", x"ec", x"ec", 
        x"eb", x"e9", x"e8", x"e6", x"e4", x"e4", x"e8", x"ed", x"eb", x"e6", x"e6", x"e8", x"e9", x"e8", x"e6", 
        x"ec", x"e9", x"e7", x"e4", x"e9", x"e5", x"e5", x"e9", x"e7", x"eb", x"ec", x"e9", x"e8", x"ec", x"e9", 
        x"e7", x"e9", x"ea", x"ea", x"eb", x"ee", x"eb", x"e8", x"e9", x"eb", x"eb", x"ea", x"ec", x"ec", x"ed", 
        x"ec", x"e5", x"e6", x"ef", x"ee", x"ea", x"ed", x"ed", x"e9", x"ea", x"ec", x"ec", x"e9", x"ea", x"ea", 
        x"ea", x"ed", x"ec", x"eb", x"ed", x"eb", x"ee", x"ea", x"e6", x"e9", x"ed", x"ef", x"e5", x"e7", x"ed", 
        x"ec", x"e8", x"e9", x"ea", x"eb", x"ea", x"ec", x"ec", x"ec", x"ec", x"ed", x"f0", x"ed", x"eb", x"ec", 
        x"ee", x"eb", x"ed", x"ed", x"ed", x"ef", x"ef", x"ee", x"f0", x"ee", x"ed", x"eb", x"ea", x"e8", x"ea", 
        x"eb", x"ef", x"ed", x"ea", x"eb", x"ed", x"ed", x"ec", x"ea", x"ea", x"eb", x"ec", x"ee", x"ee", x"ec", 
        x"ec", x"ec", x"e1", x"e5", x"ed", x"e7", x"e6", x"e7", x"ef", x"ed", x"ea", x"eb", x"ed", x"ed", x"f0", 
        x"ef", x"e9", x"e7", x"eb", x"ea", x"e8", x"e9", x"ec", x"ed", x"ed", x"ec", x"ee", x"eb", x"eb", x"ec", 
        x"ed", x"eb", x"eb", x"ea", x"eb", x"ec", x"ee", x"ea", x"ea", x"e8", x"ea", x"ee", x"ef", x"ee", x"ec", 
        x"ed", x"ec", x"ec", x"ec", x"ed", x"ed", x"ed", x"eb", x"ee", x"ed", x"e9", x"e8", x"ec", x"ed", x"eb", 
        x"eb", x"ec", x"eb", x"ea", x"ef", x"f1", x"ec", x"e9", x"ea", x"eb", x"e9", x"e8", x"ec", x"ec", x"eb", 
        x"e7", x"df", x"eb", x"ee", x"ef", x"ef", x"ed", x"ec", x"ea", x"ec", x"f0", x"ec", x"e1", x"ea", x"ec", 
        x"ec", x"ef", x"ee", x"ee", x"ee", x"f0", x"ef", x"ef", x"ee", x"ef", x"f0", x"f0", x"ee", x"ef", x"ec", 
        x"ee", x"ef", x"ee", x"ef", x"f0", x"f1", x"f0", x"ec", x"ed", x"ee", x"ef", x"f0", x"ed", x"ee", x"f0", 
        x"ef", x"ef", x"ee", x"ed", x"f0", x"f0", x"f2", x"f4", x"f5", x"f5", x"f5", x"f5", x"f3", x"f1", x"f1", 
        x"f0", x"ef", x"f0", x"e9", x"e2", x"ef", x"ed", x"ee", x"ef", x"f1", x"f2", x"f2", x"f0", x"f1", x"f1", 
        x"ef", x"ee", x"ee", x"f0", x"ef", x"f0", x"f1", x"ef", x"ec", x"ec", x"ee", x"f0", x"ef", x"ef", x"f0", 
        x"f1", x"f3", x"f1", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f0", x"f5", x"f7", x"f5", x"f2", x"f0", 
        x"f0", x"ee", x"f0", x"f0", x"ef", x"eb", x"ea", x"ee", x"ec", x"ed", x"ee", x"ed", x"e9", x"e9", x"ee", 
        x"f0", x"f0", x"ef", x"ed", x"ed", x"ee", x"f0", x"f0", x"ed", x"ee", x"f0", x"f1", x"f1", x"f0", x"f2", 
        x"ef", x"ef", x"f1", x"f1", x"f0", x"ef", x"f0", x"ef", x"ee", x"ef", x"f0", x"f1", x"f3", x"f4", x"f1", 
        x"ed", x"ee", x"f0", x"ee", x"ec", x"ef", x"ef", x"ee", x"f0", x"f0", x"f2", x"ef", x"f1", x"e8", x"b5", 
        x"9f", x"be", x"ea", x"ed", x"ee", x"ef", x"f0", x"ed", x"ec", x"ec", x"f0", x"ee", x"eb", x"ee", x"ed", 
        x"e6", x"89", x"2c", x"12", x"21", x"58", x"ce", x"ef", x"ea", x"eb", x"e9", x"ee", x"f4", x"f3", x"ee", 
        x"ec", x"f1", x"f2", x"f1", x"f1", x"ee", x"ef", x"f2", x"f1", x"b3", x"40", x"67", x"cd", x"de", x"d9", 
        x"d7", x"d6", x"db", x"9c", x"87", x"e5", x"bf", x"87", x"7e", x"7e", x"79", x"7a", x"7b", x"76", x"72", 
        x"75", x"79", x"75", x"74", x"72", x"6e", x"6a", x"66", x"69", x"67", x"66", x"61", x"62", x"5e", x"33", 
        x"27", x"39", x"3b", x"34", x"4a", x"59", x"52", x"5a", x"58", x"55", x"58", x"4b", x"42", x"3f", x"3c", 
        x"32", x"36", x"55", x"47", x"43", x"4f", x"4e", x"4c", x"4b", x"4f", x"4c", x"42", x"41", x"46", x"4f", 
        x"41", x"26", x"26", x"48", x"4e", x"45", x"47", x"45", x"48", x"4b", x"38", x"1a", x"0d", x"07", x"05", 
        x"18", x"19", x"17", x"1d", x"18", x"13", x"09", x"17", x"20", x"34", x"46", x"35", x"21", x"2d", x"25", 
        x"63", x"90", x"9e", x"58", x"09", x"0d", x"33", x"48", x"54", x"62", x"a3", x"ac", x"c6", x"a5", x"26", 
        x"0e", x"1d", x"23", x"1e", x"3b", x"55", x"51", x"59", x"5a", x"57", x"4c", x"28", x"3d", x"33", x"12", 
        x"05", x"06", x"12", x"33", x"39", x"36", x"2e", x"38", x"3b", x"31", x"32", x"1c", x"04", x"02", x"0b", 
        x"38", x"3e", x"3e", x"66", x"be", x"68", x"21", x"3a", x"75", x"69", x"42", x"25", x"34", x"4f", x"5f", 
        x"44", x"1f", x"20", x"65", x"dc", x"cd", x"cb", x"dc", x"cc", x"c9", x"cf", x"e3", x"e0", x"de", x"df", 
        x"e0", x"de", x"e2", x"e5", x"db", x"df", x"df", x"de", x"e8", x"e5", x"e3", x"e0", x"dd", x"ec", x"e1", 
        x"de", x"e2", x"e4", x"e1", x"e6", x"ea", x"e6", x"e0", x"df", x"e3", x"e3", x"e5", x"e5", x"df", x"e3", 
        x"e8", x"ea", x"e6", x"e7", x"e7", x"e5", x"e8", x"e8", x"e5", x"e6", x"e6", x"e9", x"e8", x"e7", x"e6", 
        x"e5", x"e5", x"e4", x"e4", x"e6", x"e8", x"e5", x"e2", x"e8", x"e6", x"e6", x"e8", x"e4", x"ea", x"df", 
        x"e1", x"e7", x"e9", x"e5", x"e3", x"e4", x"e6", x"e7", x"e3", x"e3", x"e7", x"e4", x"e4", x"e9", x"e8", 
        x"e2", x"da", x"db", x"e7", x"dd", x"e6", x"ef", x"e8", x"e8", x"e7", x"e7", x"e5", x"e9", x"ea", x"e7", 
        x"e6", x"e5", x"e7", x"e8", x"e4", x"ea", x"ea", x"e4", x"e1", x"e8", x"e3", x"e5", x"ef", x"eb", x"e8", 
        x"e9", x"e6", x"e4", x"e4", x"e9", x"ec", x"e9", x"eb", x"e9", x"e3", x"e6", x"e8", x"e9", x"e6", x"e6", 
        x"e3", x"e3", x"e8", x"ea", x"e8", x"eb", x"e7", x"eb", x"e7", x"e1", x"e2", x"e7", x"e8", x"e6", x"e5", 
        x"df", x"e2", x"ea", x"e6", x"e9", x"ed", x"eb", x"e7", x"e5", x"e8", x"e9", x"e9", x"e9", x"ea", x"e9", 
        x"ea", x"ea", x"e8", x"e6", x"e6", x"e8", x"ea", x"ea", x"ea", x"e4", x"e5", x"e7", x"e8", x"eb", x"ea", 
        x"e8", x"e0", x"e2", x"e6", x"ea", x"dd", x"df", x"e6", x"e4", x"ea", x"e8", x"e1", x"df", x"ec", x"eb", 
        x"e8", x"eb", x"ea", x"eb", x"e9", x"e9", x"e9", x"eb", x"ed", x"ed", x"ed", x"eb", x"ec", x"eb", x"ef", 
        x"ef", x"ea", x"e9", x"ec", x"ed", x"ed", x"f1", x"ef", x"e8", x"e6", x"ea", x"e8", x"ed", x"ec", x"e9", 
        x"e7", x"ec", x"ea", x"eb", x"ee", x"eb", x"ed", x"ea", x"e9", x"ec", x"ee", x"ee", x"e6", x"ea", x"ea", 
        x"ec", x"ec", x"ec", x"eb", x"ea", x"eb", x"e9", x"e8", x"eb", x"eb", x"eb", x"ee", x"eb", x"e7", x"eb", 
        x"ee", x"ed", x"ef", x"ed", x"eb", x"ec", x"eb", x"e9", x"ec", x"ec", x"eb", x"e9", x"eb", x"ea", x"eb", 
        x"eb", x"ef", x"ec", x"e9", x"eb", x"ee", x"ee", x"ee", x"ed", x"ec", x"eb", x"eb", x"ec", x"ec", x"ea", 
        x"ed", x"ed", x"de", x"e1", x"ea", x"ea", x"ea", x"e6", x"eb", x"ec", x"ec", x"ed", x"e9", x"e6", x"eb", 
        x"ed", x"e9", x"e6", x"ec", x"ec", x"ea", x"e9", x"e9", x"e8", x"e9", x"e9", x"eb", x"e7", x"e9", x"eb", 
        x"ed", x"eb", x"ee", x"eb", x"ec", x"ed", x"ee", x"e9", x"ea", x"e9", x"ea", x"eb", x"ec", x"eb", x"eb", 
        x"ec", x"eb", x"eb", x"eb", x"eb", x"eb", x"ea", x"ea", x"ef", x"ee", x"ed", x"eb", x"ed", x"ee", x"ee", 
        x"ec", x"ee", x"ec", x"e9", x"f0", x"ee", x"ec", x"ed", x"ed", x"ee", x"ee", x"ed", x"ed", x"ed", x"ea", 
        x"e6", x"de", x"ea", x"ee", x"ee", x"f2", x"f2", x"ef", x"ed", x"ef", x"f4", x"f3", x"e6", x"ef", x"ee", 
        x"ec", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ee", x"f0", x"f0", x"ee", x"f1", x"ed", 
        x"ee", x"ef", x"ec", x"ed", x"ed", x"f2", x"f1", x"ee", x"ee", x"ed", x"ef", x"f1", x"ee", x"ed", x"ef", 
        x"ef", x"f0", x"f1", x"ee", x"ee", x"ef", x"f2", x"f4", x"f5", x"f5", x"f4", x"f6", x"f3", x"f2", x"f2", 
        x"f0", x"ee", x"ef", x"e9", x"e2", x"ef", x"eb", x"ee", x"ee", x"f0", x"f0", x"ee", x"ed", x"f0", x"f0", 
        x"ef", x"ef", x"ee", x"f0", x"ef", x"f0", x"f1", x"ef", x"ed", x"ed", x"ed", x"ee", x"ee", x"ec", x"eb", 
        x"ed", x"f0", x"f2", x"f0", x"f1", x"f1", x"f0", x"f0", x"f2", x"f0", x"f5", x"f7", x"f4", x"f1", x"f0", 
        x"ee", x"ec", x"ef", x"f0", x"ef", x"eb", x"ea", x"ee", x"ed", x"ed", x"ee", x"ed", x"ea", x"e9", x"ee", 
        x"ef", x"f0", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", x"f1", x"f2", x"f0", x"ef", x"f0", 
        x"ee", x"ef", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f0", x"f2", x"f5", x"f3", 
        x"ef", x"ed", x"ef", x"ef", x"ee", x"f0", x"ef", x"ec", x"f0", x"ee", x"ed", x"f0", x"ec", x"aa", x"3a", 
        x"29", x"40", x"b3", x"ed", x"eb", x"ef", x"ef", x"ed", x"ec", x"ed", x"f0", x"ef", x"ed", x"ed", x"ee", 
        x"c9", x"53", x"14", x"09", x"0c", x"14", x"a4", x"ed", x"ed", x"ee", x"ee", x"f1", x"f5", x"f4", x"f0", 
        x"ee", x"f2", x"f3", x"f1", x"f0", x"ed", x"ed", x"ef", x"ef", x"b5", x"3c", x"60", x"c6", x"db", x"d7", 
        x"d6", x"d6", x"dc", x"a6", x"85", x"e6", x"d8", x"9c", x"78", x"81", x"7e", x"7a", x"7f", x"7c", x"77", 
        x"74", x"79", x"76", x"72", x"70", x"71", x"6c", x"66", x"64", x"59", x"59", x"54", x"51", x"4e", x"33", 
        x"21", x"2d", x"4c", x"46", x"2d", x"42", x"52", x"4b", x"48", x"4e", x"5e", x"61", x"59", x"4f", x"49", 
        x"33", x"39", x"5f", x"54", x"4a", x"49", x"4d", x"4e", x"51", x"4b", x"4a", x"47", x"43", x"43", x"45", 
        x"3b", x"24", x"27", x"49", x"4e", x"42", x"45", x"43", x"46", x"4a", x"45", x"2b", x"0d", x"03", x"05", 
        x"19", x"18", x"15", x"15", x"16", x"17", x"11", x"1e", x"13", x"25", x"30", x"19", x"0d", x"25", x"30", 
        x"74", x"94", x"a2", x"62", x"09", x"04", x"1b", x"40", x"57", x"61", x"9c", x"aa", x"c5", x"90", x"16", 
        x"0e", x"20", x"23", x"1f", x"3a", x"54", x"50", x"5a", x"5c", x"57", x"4e", x"2a", x"3a", x"24", x"08", 
        x"06", x"07", x"11", x"30", x"34", x"30", x"31", x"32", x"23", x"0e", x"0d", x"07", x"02", x"04", x"0b", 
        x"3e", x"31", x"2c", x"56", x"b7", x"89", x"75", x"8a", x"7b", x"71", x"4b", x"1e", x"37", x"44", x"2b", 
        x"29", x"3d", x"1f", x"65", x"d1", x"cc", x"cc", x"dd", x"ce", x"c8", x"ca", x"dc", x"dc", x"dc", x"df", 
        x"e7", x"e1", x"e0", x"e5", x"df", x"e1", x"e3", x"e7", x"eb", x"e3", x"dc", x"e2", x"e5", x"e9", x"e3", 
        x"e4", x"eb", x"ec", x"e5", x"e2", x"e4", x"e8", x"e7", x"e4", x"e5", x"e5", x"e7", x"e6", x"df", x"e7", 
        x"eb", x"e6", x"e5", x"e8", x"e7", x"e2", x"e5", x"e5", x"e4", x"e7", x"e7", x"e8", x"e6", x"e6", x"e5", 
        x"e4", x"e3", x"e6", x"e8", x"e5", x"e6", x"e8", x"e9", x"ea", x"e4", x"e0", x"eb", x"e8", x"ea", x"e4", 
        x"e7", x"e7", x"e5", x"e5", x"e5", x"e4", x"e5", x"ea", x"e7", x"e3", x"e4", x"e3", x"e4", x"ea", x"eb", 
        x"e6", x"e0", x"e0", x"e3", x"de", x"e4", x"eb", x"e9", x"e9", x"e5", x"e5", x"e3", x"eb", x"ed", x"e8", 
        x"e9", x"e6", x"e5", x"e6", x"e5", x"ee", x"ed", x"e7", x"e6", x"e5", x"df", x"df", x"e4", x"e0", x"e2", 
        x"e6", x"e8", x"ea", x"e9", x"e9", x"e8", x"e9", x"ea", x"e7", x"e4", x"e8", x"eb", x"ec", x"e8", x"e7", 
        x"e6", x"e8", x"e6", x"e4", x"e7", x"ea", x"e9", x"eb", x"ec", x"e9", x"e8", x"e6", x"e5", x"e5", x"e8", 
        x"e4", x"e5", x"e9", x"e5", x"e6", x"ea", x"ea", x"e8", x"e8", x"e9", x"ea", x"ea", x"eb", x"ec", x"eb", 
        x"e9", x"e9", x"e7", x"e6", x"e8", x"eb", x"ea", x"e8", x"e7", x"e5", x"e7", x"e8", x"e8", x"ed", x"ed", 
        x"e4", x"e2", x"e4", x"e3", x"e7", x"df", x"e3", x"e8", x"e3", x"e7", x"e7", x"e7", x"e9", x"ed", x"ea", 
        x"e9", x"ec", x"ed", x"ee", x"e9", x"e2", x"e2", x"ea", x"ec", x"ea", x"eb", x"ec", x"ee", x"ec", x"ec", 
        x"ec", x"ec", x"ea", x"e9", x"e9", x"e9", x"ef", x"ec", x"e5", x"e6", x"ec", x"ea", x"e6", x"e7", x"e7", 
        x"e8", x"ed", x"eb", x"eb", x"ea", x"e9", x"eb", x"ea", x"eb", x"ea", x"eb", x"ef", x"eb", x"eb", x"e8", 
        x"ea", x"ed", x"ec", x"e9", x"ea", x"eb", x"e9", x"e9", x"ee", x"ec", x"e9", x"f1", x"ed", x"e8", x"e9", 
        x"ea", x"e9", x"ec", x"ee", x"eb", x"eb", x"ea", x"eb", x"ee", x"ed", x"eb", x"e9", x"ec", x"eb", x"eb", 
        x"ea", x"ec", x"eb", x"ec", x"ed", x"ed", x"ee", x"ec", x"eb", x"ec", x"ed", x"ee", x"ef", x"ee", x"eb", 
        x"ea", x"ea", x"dc", x"df", x"eb", x"ee", x"f1", x"ed", x"ed", x"eb", x"ea", x"ed", x"e9", x"e4", x"e8", 
        x"ed", x"e8", x"e3", x"e8", x"e7", x"e6", x"e7", x"e8", x"e6", x"e9", x"ea", x"ec", x"e8", x"ea", x"eb", 
        x"ec", x"ec", x"ee", x"ec", x"ed", x"eb", x"ea", x"eb", x"ed", x"eb", x"ec", x"ed", x"ee", x"ee", x"ec", 
        x"eb", x"ec", x"ed", x"ed", x"ec", x"eb", x"ea", x"eb", x"ec", x"ec", x"ee", x"ee", x"ee", x"e9", x"eb", 
        x"ea", x"ed", x"ec", x"eb", x"ef", x"ee", x"ed", x"ef", x"ef", x"ed", x"ed", x"ed", x"ec", x"eb", x"eb", 
        x"e8", x"e0", x"ea", x"ef", x"ef", x"f1", x"ee", x"ed", x"eb", x"ea", x"ed", x"f2", x"ef", x"f1", x"ef", 
        x"ec", x"ed", x"ee", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ee", x"ed", x"f0", x"ee", 
        x"ef", x"f1", x"ee", x"ef", x"ee", x"f0", x"f0", x"ee", x"ef", x"ef", x"ef", x"f1", x"ec", x"ec", x"ee", 
        x"ee", x"ef", x"f1", x"ee", x"ed", x"f0", x"f2", x"f5", x"f5", x"f5", x"f5", x"f4", x"f3", x"f2", x"f0", 
        x"ee", x"ed", x"f0", x"ea", x"e2", x"ef", x"ee", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", 
        x"ed", x"eb", x"eb", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", x"ee", x"f0", x"ef", x"ef", x"ee", x"ee", 
        x"ee", x"f0", x"f2", x"f1", x"f1", x"f2", x"f1", x"f0", x"f2", x"f3", x"f7", x"f7", x"f3", x"f1", x"f1", 
        x"f1", x"ee", x"f0", x"f1", x"f1", x"ef", x"ee", x"ef", x"ef", x"f0", x"ee", x"ee", x"ec", x"eb", x"f0", 
        x"ee", x"ee", x"f0", x"f1", x"f2", x"f1", x"ef", x"ee", x"ed", x"ee", x"f0", x"f2", x"f3", x"f2", x"f2", 
        x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"ed", x"ed", x"ef", x"ef", x"f0", x"f0", x"f2", x"f4", x"f2", 
        x"f0", x"ee", x"f0", x"f0", x"ef", x"f1", x"f1", x"f0", x"f2", x"f0", x"e8", x"f2", x"de", x"71", x"28", 
        x"60", x"6f", x"a2", x"e2", x"f0", x"ef", x"ea", x"ed", x"ef", x"ee", x"ee", x"ed", x"ee", x"f2", x"ef", 
        x"e1", x"93", x"41", x"2d", x"2b", x"11", x"8f", x"e8", x"ee", x"ea", x"ef", x"f1", x"f2", x"f3", x"f0", 
        x"ee", x"f2", x"f2", x"ef", x"f1", x"f2", x"f1", x"f0", x"f1", x"bf", x"41", x"5d", x"c1", x"dd", x"d6", 
        x"d5", x"d5", x"dc", x"aa", x"7f", x"e4", x"dc", x"aa", x"7c", x"81", x"7c", x"78", x"7e", x"7c", x"79", 
        x"75", x"77", x"73", x"72", x"71", x"6f", x"6c", x"68", x"5b", x"3f", x"3a", x"3c", x"40", x"3b", x"2c", 
        x"2e", x"53", x"9d", x"ac", x"5f", x"3c", x"41", x"43", x"45", x"50", x"4c", x"31", x"36", x"4d", x"38", 
        x"1a", x"14", x"31", x"45", x"46", x"49", x"46", x"43", x"45", x"41", x"43", x"46", x"43", x"40", x"45", 
        x"3d", x"24", x"23", x"41", x"4b", x"44", x"46", x"45", x"47", x"49", x"4c", x"3d", x"10", x"02", x"06", 
        x"13", x"16", x"11", x"11", x"1a", x"23", x"20", x"13", x"08", x"23", x"4f", x"3c", x"22", x"23", x"2d", 
        x"6b", x"93", x"a8", x"65", x"0b", x"05", x"08", x"24", x"51", x"65", x"9d", x"ae", x"aa", x"6a", x"10", 
        x"0e", x"1f", x"1e", x"15", x"33", x"4f", x"45", x"56", x"56", x"54", x"52", x"35", x"3a", x"20", x"05", 
        x"03", x"04", x"12", x"31", x"37", x"2f", x"36", x"31", x"16", x"03", x"01", x"0b", x"0b", x"04", x"0d", 
        x"44", x"2a", x"25", x"58", x"bc", x"8c", x"6b", x"8b", x"94", x"69", x"22", x"40", x"7f", x"54", x"34", 
        x"47", x"58", x"26", x"89", x"d4", x"d0", x"d5", x"dd", x"cf", x"ca", x"ce", x"e2", x"e5", x"e2", x"dd", 
        x"e6", x"e3", x"e0", x"e1", x"e2", x"e8", x"e3", x"e2", x"e5", x"e4", x"e1", x"e5", x"e3", x"e3", x"e0", 
        x"e1", x"e6", x"e8", x"e3", x"dc", x"dd", x"e7", x"ea", x"e8", x"e7", x"e5", x"e5", x"e8", x"e7", x"ea", 
        x"ec", x"e5", x"e4", x"e5", x"e3", x"e3", x"e5", x"e3", x"e1", x"e4", x"e3", x"e4", x"e4", x"e2", x"e1", 
        x"e3", x"e6", x"e7", x"e6", x"e7", x"e5", x"e4", x"e3", x"e3", x"e1", x"e0", x"e5", x"e2", x"e5", x"e4", 
        x"e5", x"e2", x"e4", x"e9", x"ea", x"e6", x"e3", x"e6", x"e4", x"e2", x"e4", x"e5", x"e7", x"e6", x"e5", 
        x"e5", x"e4", x"e4", x"e6", x"df", x"dd", x"e0", x"e4", x"e7", x"e6", x"e6", x"e4", x"e7", x"e6", x"e2", 
        x"e4", x"e5", x"e8", x"e7", x"e3", x"e9", x"eb", x"e8", x"e6", x"e9", x"e4", x"e2", x"e5", x"e8", x"eb", 
        x"e9", x"e9", x"e7", x"e6", x"e8", x"e6", x"e6", x"e8", x"e9", x"e8", x"e9", x"e8", x"e5", x"e3", x"e5", 
        x"e7", x"e7", x"e4", x"e1", x"e8", x"ea", x"ea", x"e6", x"ea", x"e9", x"e3", x"de", x"e4", x"eb", x"e9", 
        x"ea", x"e9", x"ea", x"e8", x"e8", x"ea", x"e6", x"e5", x"e8", x"ea", x"ec", x"ee", x"ef", x"ef", x"ee", 
        x"ed", x"ea", x"e6", x"e4", x"e4", x"e6", x"e8", x"eb", x"e9", x"e8", x"ec", x"eb", x"e9", x"ec", x"eb", 
        x"e6", x"e8", x"e9", x"e4", x"e8", x"e9", x"e5", x"e7", x"e5", x"eb", x"ea", x"eb", x"eb", x"ea", x"eb", 
        x"ec", x"ec", x"ec", x"ec", x"e8", x"e3", x"e4", x"eb", x"ed", x"eb", x"ed", x"ef", x"f0", x"f0", x"ea", 
        x"e7", x"eb", x"eb", x"e9", x"eb", x"ea", x"ee", x"ee", x"e7", x"e7", x"eb", x"eb", x"e9", x"ea", x"e9", 
        x"e9", x"ea", x"e8", x"e8", x"e9", x"eb", x"ea", x"e8", x"ea", x"e8", x"e8", x"ec", x"e9", x"ec", x"ec", 
        x"ed", x"ea", x"ea", x"e7", x"ea", x"eb", x"e8", x"e7", x"eb", x"ea", x"e9", x"ef", x"eb", x"ea", x"ec", 
        x"ec", x"ec", x"ed", x"eb", x"e9", x"e8", x"e8", x"e9", x"ea", x"eb", x"ee", x"ee", x"ed", x"ed", x"eb", 
        x"ea", x"ec", x"eb", x"ed", x"ed", x"ec", x"ee", x"eb", x"eb", x"ec", x"ec", x"ed", x"ef", x"ee", x"ec", 
        x"ea", x"e8", x"d8", x"d9", x"e5", x"e8", x"eb", x"eb", x"ec", x"ef", x"e8", x"ea", x"ec", x"eb", x"ed", 
        x"ee", x"ea", x"e5", x"e8", x"e8", x"e7", x"ea", x"eb", x"eb", x"eb", x"ea", x"ed", x"e9", x"eb", x"eb", 
        x"ec", x"ee", x"ed", x"e9", x"eb", x"eb", x"ea", x"eb", x"e9", x"e9", x"e9", x"e9", x"e9", x"eb", x"eb", 
        x"eb", x"ed", x"ee", x"ee", x"ed", x"ec", x"eb", x"eb", x"ec", x"eb", x"ee", x"ed", x"ec", x"e9", x"ee", 
        x"ec", x"ec", x"eb", x"e9", x"ec", x"ec", x"ec", x"ef", x"ee", x"e8", x"e8", x"eb", x"ea", x"ea", x"ed", 
        x"ec", x"e2", x"ea", x"ed", x"ed", x"f0", x"ed", x"ef", x"ef", x"ed", x"ed", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ed", x"ef", x"ee", x"ef", x"f0", x"f0", x"ef", x"f0", x"ee", x"ee", x"ed", x"ef", x"ee", 
        x"ee", x"ef", x"ed", x"ed", x"ee", x"f1", x"ef", x"ed", x"ee", x"ef", x"f0", x"f2", x"ee", x"ee", x"f0", 
        x"ee", x"ef", x"f1", x"ef", x"ee", x"f0", x"f2", x"f4", x"f5", x"f6", x"f5", x"f2", x"f3", x"f3", x"f0", 
        x"ed", x"ed", x"ef", x"eb", x"e1", x"ef", x"f0", x"f2", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f1", 
        x"f0", x"ee", x"ec", x"ee", x"ef", x"ed", x"ee", x"f0", x"f0", x"ef", x"f2", x"f1", x"f1", x"f1", x"f2", 
        x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f2", x"ef", x"f0", x"f5", x"f8", x"f6", x"f1", x"f0", x"f2", 
        x"f2", x"f1", x"f1", x"f0", x"f1", x"f0", x"ef", x"ee", x"ef", x"f0", x"ee", x"ed", x"ec", x"ec", x"f0", 
        x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ed", x"ed", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"ef", x"ed", x"ed", x"ed", x"ec", x"ec", x"ee", x"f0", x"f2", x"f4", x"f6", x"f2", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"f0", x"ed", x"ef", x"f2", x"ee", x"f5", x"e0", x"74", x"31", 
        x"76", x"85", x"a8", x"e5", x"ef", x"ef", x"ea", x"ec", x"ee", x"ee", x"ef", x"ee", x"ec", x"e9", x"f1", 
        x"e2", x"99", x"77", x"8d", x"72", x"24", x"98", x"e9", x"ec", x"ea", x"f1", x"f3", x"f1", x"f2", x"f1", 
        x"ef", x"f1", x"f1", x"ee", x"f0", x"f1", x"f1", x"ee", x"f1", x"c7", x"45", x"55", x"bb", x"e1", x"d9", 
        x"d9", x"d8", x"de", x"af", x"78", x"e1", x"d8", x"ae", x"8f", x"83", x"78", x"7b", x"7e", x"7a", x"79", 
        x"77", x"78", x"72", x"6f", x"6d", x"6d", x"70", x"70", x"60", x"3e", x"39", x"3b", x"38", x"35", x"2d", 
        x"30", x"4e", x"89", x"98", x"7e", x"47", x"3f", x"43", x"4b", x"50", x"26", x"1d", x"2b", x"2c", x"24", 
        x"22", x"35", x"32", x"45", x"40", x"42", x"46", x"42", x"41", x"46", x"48", x"48", x"45", x"43", x"48", 
        x"42", x"27", x"23", x"40", x"4c", x"46", x"43", x"44", x"44", x"44", x"4c", x"4b", x"19", x"04", x"09", 
        x"10", x"16", x"12", x"15", x"2d", x"44", x"56", x"1f", x"0b", x"20", x"49", x"3f", x"2d", x"2d", x"35", 
        x"5d", x"78", x"8f", x"5b", x"09", x"03", x"03", x"0a", x"3e", x"61", x"98", x"ae", x"99", x"4a", x"09", 
        x"0e", x"20", x"19", x"11", x"31", x"4c", x"3b", x"4f", x"4f", x"50", x"56", x"3f", x"3e", x"20", x"08", 
        x"04", x"0c", x"16", x"2d", x"3f", x"3c", x"39", x"3c", x"21", x"07", x"04", x"14", x"16", x"08", x"12", 
        x"4f", x"3c", x"30", x"5f", x"b8", x"77", x"82", x"89", x"45", x"22", x"16", x"48", x"8d", x"6f", x"48", 
        x"4b", x"34", x"31", x"90", x"d1", x"c8", x"d1", x"d8", x"ce", x"c6", x"ce", x"e5", x"e1", x"db", x"df", 
        x"e1", x"e5", x"e5", x"de", x"df", x"e5", x"e4", x"dd", x"df", x"e3", x"e5", x"dc", x"d3", x"e3", x"e3", 
        x"e1", x"e6", x"e4", x"dd", x"d8", x"de", x"e4", x"e2", x"e2", x"e6", x"e7", x"e6", x"e8", x"e7", x"e3", 
        x"e5", x"e5", x"e5", x"e5", x"df", x"e1", x"e7", x"e7", x"e2", x"e3", x"e4", x"e8", x"e3", x"e1", x"e2", 
        x"e5", x"e7", x"e7", x"e6", x"e8", x"e5", x"e4", x"e4", x"e4", x"e6", x"e6", x"e7", x"e4", x"e3", x"e4", 
        x"e8", x"e6", x"e9", x"e9", x"e9", x"e6", x"e1", x"e2", x"e2", x"e3", x"e5", x"e6", x"e9", x"e9", x"e9", 
        x"e9", x"e7", x"e7", x"e6", x"e0", x"dc", x"df", x"e4", x"e6", x"e9", x"eb", x"eb", x"e7", x"e6", x"e4", 
        x"e2", x"e8", x"e8", x"ec", x"e8", x"e6", x"e7", x"e7", x"e7", x"e9", x"e6", x"e3", x"e6", x"eb", x"ec", 
        x"e5", x"e7", x"ea", x"e9", x"e4", x"df", x"e7", x"e8", x"e7", x"e9", x"ea", x"e9", x"e6", x"e6", x"e8", 
        x"e9", x"e5", x"e8", x"e6", x"e8", x"e8", x"eb", x"e6", x"e9", x"e9", x"e6", x"e2", x"e7", x"ec", x"ec", 
        x"e9", x"e8", x"eb", x"ec", x"e9", x"ea", x"e7", x"e5", x"e7", x"e8", x"e9", x"eb", x"ec", x"ec", x"ea", 
        x"e5", x"e3", x"e7", x"ea", x"e8", x"eb", x"ef", x"ed", x"ed", x"eb", x"ec", x"e9", x"e7", x"ea", x"eb", 
        x"e9", x"e8", x"e9", x"eb", x"eb", x"eb", x"e6", x"e7", x"e6", x"ea", x"e7", x"e9", x"e8", x"e6", x"eb", 
        x"ed", x"ec", x"eb", x"ea", x"e9", x"e8", x"e5", x"e7", x"e8", x"e6", x"ea", x"ea", x"e9", x"ed", x"eb", 
        x"e8", x"ea", x"e9", x"e9", x"ec", x"e8", x"ea", x"ed", x"ea", x"e6", x"e8", x"e9", x"ec", x"ec", x"e7", 
        x"e6", x"e8", x"e9", x"ec", x"ec", x"ed", x"e9", x"e8", x"eb", x"ea", x"eb", x"ea", x"e8", x"ee", x"ed", 
        x"eb", x"e8", x"e9", x"ea", x"ef", x"ec", x"e9", x"e9", x"ea", x"e9", x"ea", x"ec", x"e9", x"ec", x"ef", 
        x"ed", x"ec", x"ed", x"ed", x"ee", x"ed", x"ee", x"ee", x"ed", x"ee", x"ec", x"eb", x"eb", x"ec", x"ea", 
        x"e9", x"eb", x"ea", x"ec", x"ec", x"ec", x"ee", x"ec", x"ec", x"ed", x"ea", x"ea", x"ea", x"ea", x"ec", 
        x"ed", x"eb", x"db", x"dd", x"ea", x"e9", x"ec", x"ed", x"ef", x"f1", x"e8", x"e9", x"ed", x"ee", x"ee", 
        x"ee", x"ed", x"e9", x"eb", x"e9", x"e8", x"eb", x"eb", x"ed", x"eb", x"e6", x"ea", x"e9", x"e9", x"e9", 
        x"ed", x"ee", x"eb", x"e9", x"eb", x"eb", x"ea", x"ec", x"eb", x"ec", x"ec", x"ea", x"ea", x"ec", x"ed", 
        x"ea", x"ec", x"ed", x"ec", x"e9", x"e7", x"e8", x"ed", x"ef", x"ef", x"f0", x"ec", x"ec", x"ed", x"f0", 
        x"ee", x"ec", x"e9", x"e8", x"eb", x"ec", x"ec", x"ee", x"ed", x"e9", x"ea", x"ee", x"ed", x"ec", x"ee", 
        x"ed", x"e2", x"ea", x"ee", x"ed", x"ef", x"ed", x"ed", x"ee", x"f0", x"ef", x"ed", x"ec", x"ec", x"ef", 
        x"f1", x"ed", x"e7", x"eb", x"ed", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"eb", x"eb", x"eb", 
        x"eb", x"ee", x"ec", x"ec", x"ef", x"f2", x"f0", x"ed", x"ef", x"ee", x"ee", x"f1", x"f2", x"f2", x"f3", 
        x"f0", x"f0", x"f1", x"ee", x"ef", x"f0", x"f1", x"f3", x"f4", x"f5", x"f4", x"ef", x"f2", x"f3", x"f1", 
        x"ee", x"ee", x"ee", x"eb", x"e1", x"ed", x"f0", x"f0", x"ed", x"ee", x"f0", x"f1", x"f1", x"f0", x"f1", 
        x"ef", x"ed", x"ec", x"ef", x"f0", x"ef", x"ed", x"ee", x"ef", x"ee", x"f0", x"ee", x"ef", x"f0", x"f1", 
        x"ef", x"ee", x"f0", x"ef", x"f1", x"f3", x"f1", x"f0", x"f0", x"f3", x"f6", x"f5", x"f1", x"ef", x"ef", 
        x"ee", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ed", x"ec", x"eb", x"eb", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"ee", x"ed", x"ed", x"ed", x"ed", x"ef", x"ef", x"ef", x"f0", x"f0", x"ee", 
        x"f0", x"f2", x"f3", x"f3", x"f1", x"f1", x"f1", x"ee", x"ed", x"ef", x"f1", x"f4", x"f6", x"f6", x"f1", 
        x"ef", x"ef", x"ef", x"ef", x"f0", x"ef", x"f1", x"f0", x"ef", x"f1", x"f1", x"ee", x"e7", x"9d", x"46", 
        x"62", x"4f", x"76", x"d8", x"ec", x"ed", x"ec", x"eb", x"eb", x"ed", x"f0", x"ef", x"ed", x"ef", x"eb", 
        x"e0", x"92", x"7a", x"af", x"9c", x"5c", x"b1", x"ea", x"eb", x"ee", x"f2", x"f1", x"f0", x"f2", x"f1", 
        x"ef", x"f1", x"f0", x"ef", x"f0", x"ef", x"ee", x"ed", x"f0", x"cd", x"48", x"4b", x"b2", x"e2", x"d9", 
        x"da", x"d9", x"de", x"b6", x"7a", x"de", x"d8", x"ad", x"a7", x"94", x"77", x"7d", x"80", x"7c", x"7b", 
        x"78", x"78", x"75", x"72", x"70", x"70", x"6b", x"64", x"58", x"3f", x"3e", x"3f", x"39", x"3e", x"33", 
        x"28", x"55", x"9d", x"a8", x"a3", x"4c", x"3d", x"47", x"4a", x"3a", x"15", x"42", x"5b", x"33", x"40", 
        x"73", x"a2", x"94", x"8c", x"50", x"49", x"4f", x"49", x"46", x"4b", x"4b", x"47", x"46", x"41", x"3e", 
        x"3f", x"28", x"22", x"40", x"4d", x"43", x"3d", x"40", x"40", x"40", x"43", x"49", x"2a", x"0a", x"06", 
        x"0b", x"0e", x"0b", x"23", x"86", x"be", x"c5", x"3a", x"05", x"0b", x"26", x"41", x"51", x"43", x"4f", 
        x"82", x"82", x"85", x"65", x"14", x"05", x"05", x"03", x"31", x"63", x"93", x"b1", x"aa", x"46", x"06", 
        x"10", x"20", x"18", x"18", x"3b", x"51", x"3e", x"4e", x"4d", x"4f", x"59", x"44", x"3b", x"1c", x"08", 
        x"05", x"13", x"18", x"12", x"2b", x"36", x"38", x"3e", x"27", x"09", x"03", x"0a", x"0b", x"04", x"0e", 
        x"49", x"39", x"30", x"4f", x"9c", x"6a", x"55", x"3b", x"2a", x"21", x"1d", x"1c", x"4b", x"6b", x"56", 
        x"77", x"7e", x"62", x"7f", x"d5", x"d0", x"dc", x"dc", x"cd", x"c6", x"cf", x"e2", x"e0", x"dd", x"e4", 
        x"df", x"e2", x"e7", x"e2", x"e5", x"e5", x"df", x"e0", x"e5", x"e2", x"db", x"d8", x"de", x"e8", x"e2", 
        x"df", x"e7", x"e6", x"e1", x"e3", x"e4", x"e5", x"e4", x"e2", x"e4", x"e4", x"e4", x"e3", x"e3", x"e3", 
        x"e6", x"e5", x"e6", x"e6", x"e9", x"e3", x"e4", x"e6", x"e7", x"e8", x"e8", x"eb", x"e7", x"e8", x"ea", 
        x"ea", x"e9", x"e8", x"e7", x"e8", x"e8", x"e9", x"ea", x"e9", x"ea", x"e6", x"e2", x"e2", x"df", x"e3", 
        x"e8", x"e3", x"e3", x"e1", x"e4", x"e5", x"e2", x"e3", x"e4", x"e5", x"e6", x"e5", x"e5", x"e7", x"ea", 
        x"e6", x"e5", x"e9", x"e4", x"df", x"e2", x"e7", x"e6", x"e2", x"e7", x"eb", x"ed", x"e9", x"ec", x"ec", 
        x"e7", x"ec", x"e6", x"ee", x"ed", x"e8", x"e6", x"e7", x"e9", x"e8", x"e8", x"e9", x"eb", x"eb", x"e8", 
        x"e4", x"e8", x"e6", x"e9", x"ea", x"e6", x"ea", x"ea", x"e7", x"e2", x"e5", x"e7", x"e5", x"e4", x"e1", 
        x"e1", x"e1", x"e9", x"eb", x"e5", x"e1", x"e8", x"e8", x"ee", x"ee", x"ef", x"ed", x"ea", x"e9", x"ed", 
        x"ea", x"e9", x"ec", x"ea", x"e1", x"e6", x"eb", x"eb", x"e9", x"e6", x"e5", x"e5", x"e7", x"e8", x"ea", 
        x"e9", x"e9", x"ef", x"ee", x"e7", x"e4", x"e9", x"eb", x"ef", x"ec", x"e9", x"e6", x"e6", x"ec", x"ea", 
        x"e7", x"e9", x"ea", x"eb", x"e6", x"e8", x"e6", x"e6", x"e6", x"e9", x"e7", x"ec", x"eb", x"e5", x"e9", 
        x"eb", x"eb", x"eb", x"ea", x"eb", x"f0", x"eb", x"e9", x"eb", x"e9", x"ec", x"eb", x"e9", x"eb", x"ea", 
        x"eb", x"ec", x"eb", x"e7", x"e4", x"e1", x"e4", x"ea", x"ea", x"e5", x"e7", x"e8", x"eb", x"ee", x"ea", 
        x"e9", x"e8", x"e7", x"ea", x"e8", x"e8", x"e4", x"e6", x"e8", x"ea", x"ed", x"e9", x"ea", x"ef", x"e9", 
        x"e6", x"e8", x"ed", x"ec", x"f0", x"ea", x"e9", x"ec", x"ee", x"ec", x"ea", x"ea", x"e8", x"ed", x"ef", 
        x"eb", x"ea", x"eb", x"eb", x"ee", x"ed", x"ec", x"eb", x"e9", x"eb", x"ea", x"ea", x"ec", x"ef", x"ed", 
        x"ec", x"ed", x"ec", x"eb", x"eb", x"ec", x"ec", x"ed", x"ed", x"ed", x"ec", x"eb", x"e9", x"ea", x"eb", 
        x"ea", x"e7", x"d8", x"db", x"eb", x"e9", x"eb", x"ea", x"e9", x"ed", x"e9", x"eb", x"eb", x"ea", x"eb", 
        x"ea", x"ec", x"e9", x"eb", x"e8", x"ea", x"ed", x"eb", x"eb", x"ea", x"e5", x"ea", x"ea", x"ed", x"ec", 
        x"ed", x"eb", x"e8", x"eb", x"ec", x"ed", x"eb", x"e9", x"e8", x"ea", x"ea", x"e9", x"e8", x"e9", x"eb", 
        x"e9", x"eb", x"ed", x"ec", x"ea", x"ea", x"eb", x"ec", x"ee", x"ee", x"ee", x"e8", x"e9", x"ed", x"ee", 
        x"ee", x"eb", x"e8", x"ea", x"ed", x"ee", x"ec", x"ed", x"ed", x"ed", x"ed", x"ed", x"ec", x"eb", x"ec", 
        x"ec", x"e1", x"ea", x"f0", x"ef", x"f0", x"f0", x"f0", x"ef", x"f1", x"f3", x"ef", x"f0", x"ee", x"ee", 
        x"f0", x"ea", x"e4", x"ea", x"ec", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ec", x"ed", x"ee", 
        x"ee", x"f2", x"f1", x"f0", x"f1", x"f1", x"f0", x"ef", x"f2", x"ef", x"ec", x"ef", x"f3", x"f2", x"f4", 
        x"f2", x"f1", x"f1", x"ed", x"ef", x"ef", x"f0", x"f3", x"f5", x"f3", x"f1", x"ef", x"f1", x"f1", x"ef", 
        x"ef", x"ef", x"ee", x"ec", x"e1", x"ed", x"f0", x"ec", x"ec", x"ef", x"ec", x"e9", x"ec", x"ee", x"f1", 
        x"f2", x"f1", x"f0", x"ee", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ef", x"f2", x"f3", 
        x"f2", x"f1", x"f1", x"ef", x"f0", x"f1", x"f0", x"f1", x"f3", x"f5", x"f7", x"f7", x"f5", x"f3", x"f1", 
        x"ed", x"f1", x"f0", x"f1", x"ee", x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"ec", x"eb", x"e9", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"f0", x"f3", x"f4", x"f2", x"ef", x"ee", x"eb", x"e8", 
        x"ea", x"ed", x"ef", x"f0", x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", x"f2", x"f3", x"f4", x"f3", x"f1", 
        x"f0", x"f1", x"f0", x"f1", x"f2", x"f0", x"ef", x"ed", x"ec", x"ec", x"ee", x"ec", x"ec", x"bb", x"79", 
        x"7e", x"62", x"77", x"d5", x"f2", x"f0", x"ef", x"eb", x"ea", x"ec", x"f0", x"f0", x"ec", x"ec", x"ee", 
        x"f2", x"c8", x"73", x"79", x"a4", x"cf", x"e2", x"e9", x"eb", x"ea", x"f4", x"f3", x"f1", x"f1", x"f0", 
        x"ee", x"f0", x"f1", x"f0", x"f2", x"ef", x"ef", x"f1", x"f2", x"d9", x"51", x"45", x"aa", x"e4", x"d7", 
        x"d9", x"d7", x"dc", x"ba", x"7d", x"d5", x"d8", x"ad", x"b9", x"b4", x"79", x"76", x"7c", x"7a", x"79", 
        x"74", x"75", x"77", x"74", x"70", x"6e", x"59", x"43", x"42", x"43", x"45", x"41", x"42", x"4d", x"3d", 
        x"24", x"30", x"78", x"ba", x"9b", x"45", x"3b", x"4f", x"4b", x"36", x"12", x"3a", x"47", x"30", x"41", 
        x"59", x"7d", x"a1", x"a6", x"4d", x"3f", x"40", x"3a", x"45", x"4c", x"4a", x"44", x"45", x"45", x"3f", 
        x"3f", x"29", x"21", x"42", x"4f", x"45", x"40", x"44", x"43", x"40", x"3e", x"49", x"50", x"28", x"07", 
        x"05", x"05", x"20", x"71", x"a5", x"be", x"e4", x"57", x"09", x"06", x"08", x"32", x"53", x"47", x"45", 
        x"64", x"73", x"6e", x"65", x"28", x"06", x"03", x"02", x"1f", x"5e", x"90", x"ab", x"9a", x"2a", x"03", 
        x"0d", x"19", x"16", x"29", x"48", x"57", x"48", x"52", x"51", x"54", x"5a", x"46", x"2c", x"0e", x"03", 
        x"02", x"10", x"22", x"15", x"24", x"34", x"3e", x"2f", x"18", x"06", x"04", x"03", x"02", x"02", x"06", 
        x"4f", x"37", x"2a", x"51", x"c3", x"9d", x"3c", x"2a", x"2a", x"24", x"21", x"24", x"35", x"32", x"36", 
        x"51", x"60", x"3c", x"79", x"cf", x"c0", x"d0", x"db", x"ca", x"c1", x"cb", x"df", x"e4", x"e0", x"da", 
        x"de", x"de", x"e1", x"e1", x"e6", x"e3", x"df", x"e0", x"e3", x"e5", x"dc", x"db", x"e4", x"e7", x"e5", 
        x"e0", x"e3", x"e3", x"e6", x"e8", x"e4", x"e2", x"e2", x"e4", x"e9", x"e7", x"e7", x"e7", x"e2", x"e4", 
        x"e6", x"e9", x"e5", x"d4", x"e3", x"e7", x"e3", x"e6", x"e6", x"e4", x"e1", x"e7", x"ea", x"e9", x"e9", 
        x"e9", x"e8", x"e5", x"e2", x"e2", x"e4", x"e4", x"e4", x"e4", x"e8", x"e2", x"de", x"e6", x"e6", x"e7", 
        x"e6", x"e1", x"e6", x"e3", x"e4", x"e5", x"e2", x"e4", x"e6", x"e7", x"e6", x"e6", x"e5", x"e3", x"e6", 
        x"e4", x"e0", x"e6", x"e7", x"df", x"e1", x"e6", x"e1", x"db", x"e5", x"e9", x"e9", x"e9", x"ec", x"ea", 
        x"e5", x"e5", x"e5", x"e9", x"e7", x"e7", x"e9", x"e9", x"ea", x"e9", x"e9", x"e9", x"ea", x"e9", x"e6", 
        x"e6", x"eb", x"ea", x"ef", x"ec", x"e5", x"eb", x"e8", x"e5", x"e7", x"e9", x"ea", x"e8", x"e7", x"e2", 
        x"e2", x"e4", x"e8", x"ea", x"e6", x"e3", x"e8", x"e9", x"eb", x"ea", x"ea", x"e8", x"e8", x"e8", x"eb", 
        x"ec", x"ec", x"ee", x"ed", x"e3", x"e6", x"eb", x"eb", x"ea", x"e7", x"e7", x"e9", x"eb", x"eb", x"e9", 
        x"e4", x"e8", x"ee", x"ee", x"e8", x"e7", x"eb", x"ec", x"ec", x"e9", x"eb", x"ee", x"ee", x"ee", x"ea", 
        x"e5", x"ec", x"eb", x"ea", x"e8", x"e8", x"e5", x"e7", x"e7", x"ea", x"e7", x"ed", x"ea", x"e9", x"eb", 
        x"e9", x"ea", x"ed", x"e7", x"e4", x"eb", x"e8", x"e9", x"ee", x"eb", x"ec", x"eb", x"ea", x"ec", x"ed", 
        x"ee", x"ec", x"e9", x"e6", x"e2", x"e7", x"e9", x"e9", x"e5", x"e3", x"e8", x"ea", x"e5", x"ea", x"e8", 
        x"ea", x"ea", x"ea", x"ec", x"ea", x"e8", x"e5", x"e7", x"e7", x"ea", x"ec", x"e9", x"ea", x"eb", x"eb", 
        x"ea", x"e9", x"ee", x"ea", x"ec", x"ec", x"e9", x"e9", x"ed", x"ec", x"ea", x"ec", x"e9", x"ef", x"f0", 
        x"eb", x"ec", x"ed", x"ed", x"f1", x"ef", x"ec", x"ea", x"e8", x"ed", x"ef", x"ef", x"ee", x"f0", x"ed", 
        x"ec", x"ed", x"ef", x"eb", x"ec", x"ec", x"eb", x"ed", x"ec", x"eb", x"eb", x"ea", x"e8", x"ea", x"ed", 
        x"ee", x"eb", x"dd", x"da", x"e8", x"e9", x"ed", x"ec", x"e9", x"eb", x"ea", x"ec", x"eb", x"ea", x"eb", 
        x"eb", x"ea", x"e9", x"ea", x"e8", x"ea", x"ec", x"e9", x"e7", x"ea", x"e7", x"e7", x"e8", x"ed", x"e9", 
        x"ea", x"e9", x"e5", x"eb", x"ec", x"ee", x"ec", x"eb", x"ec", x"eb", x"ec", x"ed", x"ee", x"ed", x"eb", 
        x"e9", x"eb", x"ec", x"eb", x"ea", x"eb", x"ed", x"ed", x"ec", x"ec", x"ee", x"e9", x"e8", x"ea", x"ec", 
        x"f0", x"ef", x"ea", x"ec", x"ee", x"ec", x"ec", x"ec", x"eb", x"ed", x"ee", x"ed", x"ee", x"ed", x"ed", 
        x"ec", x"e0", x"ea", x"f1", x"ed", x"ed", x"ed", x"ee", x"ec", x"ec", x"ef", x"ea", x"ed", x"ee", x"ec", 
        x"ef", x"ee", x"ec", x"f3", x"f0", x"ef", x"ef", x"ee", x"ed", x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", 
        x"ed", x"ef", x"ee", x"ec", x"ef", x"f0", x"ee", x"ee", x"f1", x"f0", x"ee", x"f0", x"f0", x"f0", x"f3", 
        x"f3", x"f2", x"f1", x"ec", x"ee", x"ef", x"f1", x"f5", x"f6", x"f2", x"ed", x"ef", x"f1", x"ef", x"ec", 
        x"ee", x"f0", x"ef", x"ee", x"e3", x"ee", x"f0", x"eb", x"ec", x"f1", x"f1", x"ee", x"f1", x"f0", x"f2", 
        x"f2", x"ee", x"ee", x"ed", x"ee", x"f1", x"f1", x"ef", x"f0", x"f1", x"f0", x"f0", x"f2", x"f3", x"f3", 
        x"f3", x"f2", x"ef", x"ed", x"f0", x"f2", x"f2", x"f2", x"f4", x"f7", x"f8", x"f6", x"f2", x"f2", x"f1", 
        x"ef", x"ef", x"ef", x"f2", x"f0", x"f0", x"f0", x"ef", x"ef", x"ee", x"ee", x"ed", x"eb", x"e9", x"ee", 
        x"ef", x"f0", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"f0", x"f2", x"f2", x"ef", x"f1", x"f0", x"ed", 
        x"ef", x"f0", x"f0", x"ed", x"ec", x"ee", x"f2", x"ef", x"ee", x"ef", x"f1", x"f3", x"f4", x"f2", x"ef", 
        x"ee", x"f0", x"ee", x"ef", x"f1", x"ef", x"ed", x"ee", x"ef", x"ef", x"ee", x"f0", x"d9", x"83", x"5e", 
        x"5a", x"50", x"61", x"b1", x"eb", x"f0", x"ef", x"ee", x"ed", x"ee", x"ef", x"ef", x"ed", x"ed", x"e9", 
        x"ef", x"e5", x"bb", x"89", x"96", x"c6", x"d6", x"d6", x"e1", x"ec", x"f4", x"f1", x"f0", x"f1", x"f0", 
        x"ee", x"f0", x"f1", x"f2", x"f4", x"ef", x"f0", x"f4", x"f1", x"dd", x"57", x"43", x"a7", x"e6", x"d6", 
        x"d8", x"d7", x"df", x"c1", x"79", x"d4", x"d6", x"a8", x"b7", x"d7", x"9b", x"83", x"82", x"7d", x"7d", 
        x"77", x"75", x"74", x"74", x"71", x"71", x"54", x"34", x"34", x"36", x"3c", x"3d", x"3e", x"45", x"38", 
        x"1f", x"24", x"7f", x"c7", x"b1", x"55", x"17", x"2b", x"45", x"45", x"14", x"16", x"2c", x"4a", x"56", 
        x"3d", x"53", x"9f", x"b1", x"4a", x"15", x"16", x"16", x"21", x"2f", x"42", x"43", x"39", x"3c", x"44", 
        x"46", x"2c", x"23", x"42", x"4f", x"46", x"41", x"44", x"42", x"46", x"45", x"45", x"67", x"51", x"15", 
        x"05", x"04", x"30", x"96", x"bd", x"ac", x"d1", x"53", x"0a", x"07", x"04", x"0d", x"21", x"2f", x"31", 
        x"59", x"68", x"2f", x"28", x"19", x"07", x"03", x"03", x"10", x"4b", x"92", x"b1", x"98", x"29", x"04", 
        x"0b", x"12", x"13", x"35", x"4c", x"53", x"4d", x"50", x"52", x"59", x"5a", x"48", x"21", x"08", x"06", 
        x"08", x"09", x"1b", x"21", x"15", x"1d", x"31", x"16", x"07", x"03", x"04", x"04", x"05", x"03", x"04", 
        x"33", x"33", x"2a", x"4f", x"ba", x"89", x"40", x"2e", x"21", x"24", x"1f", x"25", x"28", x"2f", x"3a", 
        x"50", x"2f", x"25", x"74", x"d1", x"c6", x"cd", x"dd", x"cc", x"c3", x"cc", x"e2", x"e4", x"e2", x"e2", 
        x"e5", x"e3", x"e4", x"e2", x"e2", x"e1", x"e3", x"e2", x"e1", x"e6", x"dc", x"db", x"e1", x"e7", x"ea", 
        x"e5", x"e3", x"e6", x"e8", x"e4", x"e6", x"e1", x"e0", x"e9", x"eb", x"e8", x"e8", x"e5", x"df", x"e3", 
        x"e4", x"e7", x"e5", x"d5", x"dc", x"e9", x"e5", x"e8", x"e7", x"e1", x"e2", x"e6", x"e4", x"e7", x"e8", 
        x"e4", x"e2", x"e6", x"e6", x"e0", x"df", x"e5", x"e5", x"e2", x"e4", x"e0", x"e2", x"e9", x"e7", x"e6", 
        x"e5", x"e0", x"e3", x"e3", x"e5", x"e5", x"e2", x"e7", x"e6", x"e8", x"e7", x"e5", x"e7", x"e2", x"e7", 
        x"e3", x"dc", x"e8", x"e8", x"dd", x"e1", x"e7", x"e5", x"e2", x"e4", x"e7", x"e8", x"e9", x"eb", x"e8", 
        x"e4", x"e5", x"e4", x"e8", x"e8", x"e9", x"eb", x"ea", x"ef", x"ec", x"ea", x"e9", x"eb", x"ea", x"e6", 
        x"e9", x"ec", x"e9", x"ea", x"ea", x"e8", x"e6", x"e8", x"e8", x"e4", x"e6", x"ea", x"e9", x"e9", x"e3", 
        x"e5", x"ec", x"e9", x"ea", x"ea", x"ea", x"e9", x"e9", x"e7", x"ea", x"eb", x"e6", x"e5", x"e6", x"e9", 
        x"eb", x"ea", x"e6", x"ea", x"e5", x"e8", x"ec", x"eb", x"ea", x"e9", x"ea", x"e9", x"eb", x"ed", x"e9", 
        x"e4", x"e8", x"eb", x"eb", x"ea", x"ec", x"ed", x"ed", x"ec", x"ea", x"ec", x"ee", x"e9", x"eb", x"eb", 
        x"e7", x"eb", x"e9", x"ec", x"eb", x"e6", x"ea", x"ee", x"ec", x"ec", x"e8", x"ec", x"ea", x"eb", x"e8", 
        x"ea", x"ea", x"ea", x"eb", x"e7", x"e9", x"e9", x"e8", x"ef", x"ed", x"ed", x"ee", x"ea", x"e9", x"ed", 
        x"eb", x"e9", x"e9", x"e9", x"e7", x"ec", x"ea", x"ea", x"e8", x"e7", x"ec", x"e8", x"e5", x"ec", x"e9", 
        x"e9", x"e8", x"e9", x"eb", x"ed", x"ed", x"ea", x"ea", x"ea", x"ec", x"ed", x"ee", x"ed", x"ea", x"ec", 
        x"ed", x"e9", x"e9", x"e7", x"eb", x"ec", x"eb", x"e8", x"eb", x"e9", x"eb", x"f0", x"ea", x"ee", x"f0", 
        x"ed", x"eb", x"ed", x"ea", x"ed", x"e9", x"eb", x"ea", x"e8", x"ec", x"ec", x"ec", x"eb", x"ec", x"eb", 
        x"eb", x"ec", x"ee", x"eb", x"ec", x"ed", x"eb", x"eb", x"eb", x"ec", x"eb", x"ea", x"ea", x"ea", x"ed", 
        x"ee", x"ee", x"df", x"d9", x"e6", x"e9", x"ed", x"ee", x"ea", x"ea", x"ec", x"ea", x"e9", x"ec", x"ee", 
        x"ed", x"eb", x"e9", x"ea", x"e9", x"e8", x"ea", x"e8", x"e9", x"ec", x"ea", x"e8", x"e7", x"eb", x"e6", 
        x"e9", x"eb", x"ea", x"ec", x"eb", x"eb", x"e9", x"ec", x"ec", x"ea", x"ee", x"ef", x"ec", x"ea", x"ea", 
        x"eb", x"ec", x"ec", x"ea", x"e9", x"eb", x"ee", x"ee", x"ec", x"eb", x"ec", x"eb", x"ea", x"eb", x"eb", 
        x"ef", x"ef", x"eb", x"e9", x"ea", x"ea", x"ec", x"ec", x"eb", x"ed", x"ed", x"ed", x"f0", x"ed", x"eb", 
        x"ed", x"dd", x"e8", x"ef", x"ee", x"ee", x"ef", x"f1", x"ef", x"ee", x"ef", x"ec", x"ed", x"ee", x"eb", 
        x"ed", x"f0", x"f0", x"f1", x"ef", x"ee", x"ee", x"ed", x"ee", x"f0", x"f1", x"ef", x"ee", x"ee", x"ee", 
        x"ed", x"f0", x"ef", x"ee", x"ef", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"f2", 
        x"f1", x"f0", x"ee", x"ec", x"ed", x"ef", x"f3", x"f5", x"f6", x"f3", x"ed", x"f0", x"f2", x"ef", x"ed", 
        x"ef", x"f1", x"f0", x"ed", x"e4", x"ee", x"f1", x"ec", x"ed", x"f1", x"f0", x"ef", x"f3", x"f4", x"f3", 
        x"f1", x"ef", x"ee", x"ee", x"f0", x"f1", x"f0", x"f0", x"ef", x"f1", x"f0", x"f0", x"f2", x"f3", x"f3", 
        x"f1", x"ef", x"ee", x"ee", x"f1", x"f2", x"f0", x"ef", x"f2", x"f7", x"f7", x"f3", x"ef", x"f0", x"f1", 
        x"ef", x"ed", x"ec", x"ef", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"f1", x"ee", x"ec", x"e9", x"ed", 
        x"ee", x"ef", x"ef", x"ed", x"ed", x"ee", x"ed", x"ee", x"f0", x"f0", x"ef", x"ef", x"f1", x"f1", x"ef", 
        x"ef", x"ee", x"ed", x"ec", x"eb", x"ee", x"f1", x"ee", x"ec", x"ed", x"f1", x"f3", x"f3", x"f1", x"ef", 
        x"ef", x"f0", x"ef", x"ef", x"f0", x"ee", x"eb", x"ef", x"f0", x"f1", x"f1", x"e8", x"a7", x"65", x"49", 
        x"46", x"70", x"64", x"85", x"d0", x"ec", x"ef", x"ef", x"ec", x"eb", x"ed", x"ee", x"eb", x"f1", x"ef", 
        x"ed", x"ee", x"f3", x"cb", x"9d", x"b7", x"dc", x"d9", x"d7", x"ea", x"f2", x"ee", x"ef", x"f0", x"ef", 
        x"ee", x"f0", x"f2", x"f3", x"f4", x"f2", x"f2", x"f2", x"f1", x"e2", x"5d", x"3e", x"a4", x"e8", x"d5", 
        x"d8", x"d7", x"de", x"ca", x"79", x"d7", x"d7", x"aa", x"b1", x"d3", x"9f", x"76", x"75", x"85", x"84", 
        x"78", x"77", x"74", x"6e", x"67", x"6c", x"54", x"35", x"34", x"37", x"3a", x"39", x"3c", x"46", x"37", 
        x"15", x"23", x"90", x"cb", x"c8", x"77", x"15", x"0f", x"24", x"38", x"37", x"23", x"32", x"56", x"52", 
        x"30", x"1d", x"74", x"8e", x"2c", x"07", x"09", x"0a", x"06", x"0b", x"21", x"46", x"52", x"4f", x"46", 
        x"43", x"2e", x"23", x"41", x"52", x"44", x"40", x"41", x"42", x"47", x"42", x"3b", x"63", x"6a", x"46", 
        x"2b", x"0f", x"23", x"59", x"b4", x"ce", x"df", x"65", x"15", x"1d", x"22", x"18", x"09", x"12", x"24", 
        x"6c", x"97", x"61", x"2e", x"10", x"09", x"0a", x"07", x"05", x"2d", x"8a", x"b2", x"a3", x"3f", x"06", 
        x"14", x"14", x"15", x"36", x"47", x"50", x"4b", x"49", x"4f", x"5d", x"5c", x"4c", x"20", x"08", x"07", 
        x"09", x"08", x"10", x"1d", x"0c", x"0f", x"1a", x"0a", x"07", x"08", x"0d", x"0c", x"0b", x"07", x"0a", 
        x"1e", x"2e", x"30", x"51", x"b2", x"7d", x"48", x"2f", x"20", x"18", x"13", x"28", x"2b", x"2c", x"37", 
        x"5b", x"42", x"43", x"7c", x"cd", x"c3", x"cd", x"db", x"c4", x"c3", x"ce", x"e0", x"df", x"e3", x"e5", 
        x"e3", x"dd", x"df", x"e3", x"e3", x"e4", x"e1", x"e1", x"e3", x"e7", x"de", x"e0", x"e9", x"e7", x"e8", 
        x"e1", x"dd", x"e4", x"e2", x"db", x"e1", x"e3", x"e5", x"ed", x"eb", x"e9", x"e9", x"e1", x"df", x"dd", 
        x"d0", x"d5", x"df", x"ea", x"e9", x"ea", x"e5", x"e6", x"e8", x"e3", x"e5", x"e6", x"e6", x"e9", x"e7", 
        x"e2", x"e2", x"e9", x"e9", x"db", x"d9", x"e1", x"df", x"de", x"e5", x"e5", x"de", x"de", x"e2", x"e3", 
        x"e5", x"e6", x"e5", x"e5", x"e6", x"e5", x"e2", x"e6", x"e1", x"e3", x"e4", x"e1", x"e5", x"e2", x"e2", 
        x"e1", x"dd", x"e8", x"e6", x"de", x"e6", x"e9", x"e7", x"e8", x"e0", x"e6", x"e9", x"ea", x"e9", x"e6", 
        x"e5", x"e7", x"e9", x"e9", x"e6", x"e5", x"eb", x"ea", x"ee", x"e5", x"e3", x"e4", x"e9", x"e7", x"e5", 
        x"e9", x"ec", x"ec", x"e8", x"e7", x"e9", x"e2", x"eb", x"ee", x"e7", x"e6", x"e8", x"ec", x"eb", x"e3", 
        x"e5", x"e7", x"e7", x"e9", x"ed", x"ee", x"e6", x"e6", x"e5", x"eb", x"ec", x"e7", x"ea", x"e9", x"e8", 
        x"e4", x"e6", x"e1", x"e9", x"e5", x"e6", x"ed", x"ed", x"e7", x"e5", x"e6", x"e4", x"e6", x"ea", x"ed", 
        x"ed", x"ee", x"ea", x"ed", x"ec", x"ea", x"e8", x"ea", x"ea", x"ec", x"ed", x"e8", x"e3", x"ea", x"ef", 
        x"ec", x"e9", x"ea", x"eb", x"ea", x"e8", x"e6", x"ec", x"eb", x"ea", x"e6", x"ea", x"eb", x"ea", x"e4", 
        x"eb", x"ec", x"e7", x"e8", x"e5", x"e6", x"e9", x"e6", x"ea", x"eb", x"ed", x"ed", x"eb", x"eb", x"ed", 
        x"e7", x"e9", x"e7", x"e8", x"e9", x"ef", x"e7", x"eb", x"ee", x"e8", x"ea", x"e5", x"e3", x"ea", x"e6", 
        x"e8", x"ea", x"ec", x"ec", x"e9", x"ed", x"ef", x"e3", x"e5", x"e9", x"e8", x"eb", x"eb", x"e9", x"e7", 
        x"e3", x"e3", x"e7", x"e9", x"e9", x"e8", x"ea", x"ea", x"ed", x"e9", x"eb", x"ed", x"ea", x"ea", x"eb", 
        x"ed", x"ee", x"ef", x"ea", x"ec", x"e7", x"ed", x"eb", x"ea", x"ea", x"ea", x"ea", x"eb", x"ec", x"ec", 
        x"ee", x"ef", x"ed", x"ea", x"ea", x"ec", x"ed", x"ed", x"ed", x"ee", x"ec", x"eb", x"ed", x"ec", x"ea", 
        x"eb", x"ed", x"e1", x"dc", x"e9", x"eb", x"ec", x"ec", x"e8", x"e9", x"ec", x"e6", x"e4", x"e9", x"e9", 
        x"e8", x"ec", x"ed", x"eb", x"ec", x"eb", x"ec", x"ec", x"ec", x"ee", x"ef", x"ed", x"eb", x"ec", x"eb", 
        x"ea", x"eb", x"ed", x"ea", x"eb", x"eb", x"e8", x"ed", x"ec", x"ea", x"eb", x"e9", x"eb", x"ed", x"ec", 
        x"ef", x"ed", x"ec", x"ec", x"ed", x"ed", x"ed", x"ee", x"e9", x"e7", x"e4", x"e9", x"ec", x"ef", x"ed", 
        x"ee", x"ef", x"ec", x"e9", x"e9", x"ec", x"eb", x"eb", x"ee", x"f0", x"ed", x"ec", x"eb", x"e8", x"e9", 
        x"ef", x"de", x"e9", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", x"ec", 
        x"eb", x"ed", x"ec", x"e9", x"ec", x"ee", x"ef", x"ee", x"ed", x"ef", x"f1", x"ef", x"f0", x"f1", x"ef", 
        x"f0", x"f1", x"f1", x"f3", x"ef", x"f2", x"f2", x"f4", x"f3", x"ef", x"f1", x"f1", x"f2", x"f2", x"f3", 
        x"f1", x"ed", x"ec", x"ee", x"ee", x"f0", x"f4", x"f4", x"f4", x"f4", x"ef", x"ee", x"f1", x"ef", x"ed", 
        x"ef", x"ef", x"ee", x"eb", x"e4", x"ed", x"f2", x"ee", x"ee", x"ef", x"ee", x"ed", x"f0", x"f3", x"f0", 
        x"ed", x"ee", x"ef", x"f0", x"f1", x"ef", x"ee", x"f0", x"ef", x"ee", x"ee", x"ef", x"f1", x"f3", x"f4", 
        x"f1", x"ef", x"f0", x"ef", x"f0", x"ef", x"ec", x"ed", x"f3", x"f8", x"f7", x"f3", x"f0", x"f2", x"f2", 
        x"ef", x"ef", x"ed", x"ee", x"f2", x"f2", x"ef", x"ee", x"ef", x"f0", x"f2", x"f0", x"ed", x"e7", x"ea", 
        x"eb", x"ef", x"ee", x"ed", x"f0", x"f0", x"ee", x"f1", x"f2", x"ef", x"ed", x"ed", x"ee", x"ee", x"ee", 
        x"f0", x"ef", x"f0", x"f2", x"f1", x"f3", x"f1", x"f0", x"ed", x"ec", x"f1", x"f3", x"f1", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"ee", x"ef", x"f1", x"f2", x"e7", x"ab", x"76", x"7f", x"66", 
        x"61", x"8d", x"5e", x"6f", x"b8", x"d8", x"e6", x"f2", x"ed", x"ea", x"ec", x"ed", x"e8", x"ec", x"ed", 
        x"ef", x"f0", x"f3", x"af", x"91", x"cb", x"e3", x"d7", x"c4", x"d7", x"f2", x"f0", x"ee", x"f2", x"f1", 
        x"ef", x"ef", x"f1", x"ef", x"f0", x"f5", x"f3", x"ed", x"f0", x"e4", x"60", x"3c", x"9b", x"e7", x"d6", 
        x"db", x"d9", x"db", x"cf", x"7f", x"ce", x"df", x"ba", x"95", x"69", x"33", x"29", x"32", x"67", x"80", 
        x"73", x"76", x"7a", x"64", x"4f", x"54", x"4d", x"41", x"41", x"44", x"43", x"3f", x"46", x"38", x"1a", 
        x"0d", x"12", x"4a", x"7d", x"a3", x"7b", x"1f", x"0e", x"07", x"10", x"38", x"6f", x"81", x"7a", x"6b", 
        x"43", x"12", x"21", x"26", x"08", x"09", x"07", x"0a", x"0a", x"06", x"0a", x"67", x"ba", x"b4", x"72", 
        x"39", x"2e", x"28", x"42", x"54", x"46", x"3f", x"40", x"47", x"46", x"42", x"3d", x"57", x"70", x"5e", 
        x"42", x"18", x"23", x"3d", x"75", x"c3", x"ea", x"6e", x"19", x"2e", x"48", x"45", x"2f", x"24", x"4e", 
        x"88", x"ae", x"9f", x"48", x"27", x"38", x"3c", x"2a", x"0b", x"16", x"7c", x"aa", x"a7", x"5c", x"2f", 
        x"57", x"2a", x"10", x"28", x"35", x"49", x"44", x"44", x"50", x"5d", x"5a", x"4b", x"2b", x"12", x"0e", 
        x"12", x"19", x"15", x"13", x"13", x"14", x"13", x"17", x"1c", x"1b", x"23", x"27", x"2e", x"36", x"3a", 
        x"31", x"39", x"32", x"50", x"be", x"90", x"38", x"30", x"26", x"16", x"28", x"43", x"32", x"27", x"31", 
        x"49", x"45", x"43", x"86", x"d0", x"b9", x"c3", x"d9", x"c2", x"c3", x"ce", x"dc", x"da", x"dd", x"e2", 
        x"e2", x"de", x"e1", x"e4", x"e3", x"e3", x"e4", x"e0", x"e1", x"e4", x"e1", x"e0", x"e7", x"e9", x"e3", 
        x"df", x"d7", x"da", x"e7", x"e0", x"e0", x"ea", x"e5", x"e3", x"e5", x"e4", x"e6", x"e1", x"e6", x"e5", 
        x"d8", x"e1", x"e7", x"e8", x"e6", x"e9", x"e8", x"e7", x"e8", x"e6", x"e5", x"e3", x"e7", x"eb", x"e8", 
        x"e6", x"e9", x"e4", x"e4", x"e1", x"e3", x"e4", x"df", x"e1", x"e8", x"e9", x"e2", x"dc", x"e2", x"e2", 
        x"e2", x"e6", x"e4", x"e8", x"e8", x"e6", x"e5", x"e6", x"e2", x"e1", x"e1", x"e1", x"e6", x"e2", x"dc", 
        x"e3", x"e1", x"e2", x"e7", x"e0", x"e5", x"e6", x"e4", x"e9", x"e5", x"e8", x"e8", x"ea", x"e9", x"e9", 
        x"ec", x"e7", x"e6", x"e4", x"e4", x"e8", x"ee", x"eb", x"eb", x"e9", x"e8", x"e5", x"e8", x"ea", x"e8", 
        x"e3", x"e8", x"ed", x"ea", x"ea", x"e9", x"e2", x"e9", x"eb", x"e8", x"e2", x"de", x"e8", x"ea", x"e5", 
        x"e9", x"ea", x"e8", x"e6", x"e7", x"e7", x"e2", x"e5", x"e5", x"ea", x"ea", x"e4", x"e7", x"e8", x"e9", 
        x"e9", x"ea", x"eb", x"f1", x"eb", x"e7", x"e6", x"eb", x"e8", x"e5", x"e6", x"e5", x"e7", x"e9", x"e8", 
        x"e8", x"ed", x"e9", x"ee", x"ed", x"e8", x"e9", x"eb", x"eb", x"eb", x"ee", x"e9", x"e8", x"eb", x"ec", 
        x"e9", x"e9", x"eb", x"eb", x"eb", x"e9", x"e7", x"eb", x"ec", x"e9", x"e5", x"ec", x"ec", x"ec", x"eb", 
        x"ee", x"ef", x"ec", x"e9", x"e6", x"e9", x"eb", x"ea", x"eb", x"ea", x"ed", x"eb", x"eb", x"ed", x"ec", 
        x"e8", x"ea", x"e5", x"ea", x"ee", x"ee", x"e8", x"e9", x"e9", x"e5", x"eb", x"ec", x"ed", x"ed", x"e7", 
        x"ea", x"ea", x"e9", x"ed", x"ea", x"ea", x"eb", x"d8", x"de", x"e8", x"e8", x"ea", x"ea", x"ec", x"e9", 
        x"e5", x"e4", x"e7", x"ea", x"ea", x"ea", x"eb", x"ea", x"ee", x"ea", x"ea", x"ea", x"eb", x"eb", x"ea", 
        x"eb", x"eb", x"eb", x"ec", x"f0", x"eb", x"ec", x"ea", x"eb", x"e9", x"ea", x"eb", x"eb", x"eb", x"eb", 
        x"ed", x"f0", x"ef", x"ec", x"ea", x"eb", x"ee", x"f0", x"ed", x"eb", x"ed", x"ec", x"eb", x"ef", x"ec", 
        x"eb", x"ef", x"df", x"db", x"e8", x"eb", x"ed", x"ed", x"ea", x"e9", x"ed", x"ea", x"e8", x"eb", x"ea", 
        x"e8", x"ea", x"ee", x"ed", x"eb", x"e9", x"eb", x"ea", x"e8", x"ec", x"ef", x"ed", x"ec", x"ed", x"ef", 
        x"ed", x"ec", x"eb", x"e7", x"ea", x"ea", x"e7", x"eb", x"ea", x"e8", x"e3", x"e0", x"e7", x"ec", x"e9", 
        x"ee", x"eb", x"eb", x"ec", x"ed", x"eb", x"e8", x"ea", x"e8", x"e9", x"e9", x"eb", x"eb", x"ea", x"ee", 
        x"ee", x"ed", x"ec", x"ed", x"ed", x"ec", x"ea", x"ea", x"ee", x"ef", x"ec", x"ea", x"e8", x"e8", x"ea", 
        x"ef", x"df", x"e8", x"ef", x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ec", x"ec", 
        x"ee", x"ed", x"ea", x"eb", x"ee", x"ed", x"ef", x"f0", x"ee", x"ed", x"ef", x"f0", x"f0", x"ef", x"ec", 
        x"ee", x"ef", x"ef", x"f0", x"ee", x"ef", x"ef", x"f1", x"f0", x"ee", x"f0", x"f1", x"f2", x"f2", x"f3", 
        x"f1", x"ee", x"ed", x"f0", x"f0", x"f2", x"f3", x"f1", x"f1", x"f1", x"ee", x"ee", x"ef", x"ec", x"eb", 
        x"ec", x"ee", x"ee", x"ed", x"e6", x"ed", x"f2", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"ef", x"ee", 
        x"ed", x"ee", x"ef", x"ef", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"ef", x"f1", x"f3", x"f4", x"f4", 
        x"f2", x"f0", x"f1", x"ef", x"ee", x"ee", x"ed", x"f0", x"f5", x"f8", x"f6", x"f2", x"f0", x"f2", x"f2", 
        x"ef", x"ee", x"ed", x"ee", x"f1", x"f2", x"f0", x"ee", x"ee", x"ef", x"f1", x"ef", x"ee", x"e7", x"ec", 
        x"ec", x"ef", x"ef", x"ed", x"ef", x"f0", x"ee", x"ef", x"ef", x"ed", x"ec", x"ed", x"ef", x"f0", x"f1", 
        x"f2", x"f1", x"f1", x"f2", x"f0", x"f2", x"f1", x"f1", x"ee", x"ed", x"f1", x"f3", x"f1", x"ed", x"ef", 
        x"f0", x"f0", x"f0", x"f1", x"f2", x"f0", x"f0", x"ed", x"ee", x"ee", x"b6", x"71", x"61", x"69", x"6a", 
        x"6f", x"75", x"74", x"91", x"c5", x"ce", x"d0", x"ea", x"ef", x"ed", x"ed", x"ee", x"f0", x"ee", x"ec", 
        x"eb", x"ef", x"e6", x"a8", x"b0", x"d4", x"dd", x"d9", x"c0", x"ca", x"ed", x"f4", x"f0", x"f3", x"f2", 
        x"ef", x"ef", x"f1", x"ef", x"ef", x"f2", x"f2", x"ef", x"f1", x"e6", x"61", x"40", x"96", x"e2", x"d8", 
        x"db", x"d8", x"dd", x"d0", x"7d", x"c1", x"e1", x"c3", x"74", x"2c", x"0e", x"11", x"19", x"3b", x"68", 
        x"78", x"72", x"75", x"64", x"44", x"3c", x"40", x"44", x"40", x"3b", x"3b", x"3e", x"43", x"21", x"07", 
        x"09", x"04", x"21", x"6d", x"bd", x"a1", x"2f", x"12", x"0b", x"06", x"18", x"4f", x"6b", x"8b", x"b2", 
        x"92", x"33", x"0a", x"07", x"07", x"07", x"04", x"04", x"07", x"06", x"07", x"33", x"80", x"a1", x"97", 
        x"54", x"2e", x"26", x"3d", x"50", x"46", x"40", x"44", x"46", x"46", x"49", x"47", x"5c", x"6b", x"4e", 
        x"32", x"1e", x"24", x"41", x"4a", x"95", x"dd", x"5b", x"0d", x"19", x"3c", x"53", x"4f", x"5a", x"98", 
        x"a9", x"b5", x"a2", x"47", x"2b", x"39", x"39", x"31", x"1b", x"19", x"56", x"6c", x"6b", x"4c", x"3d", 
        x"53", x"21", x"1a", x"32", x"3e", x"3c", x"45", x"45", x"4d", x"5b", x"59", x"56", x"57", x"55", x"52", 
        x"51", x"55", x"56", x"56", x"5d", x"59", x"55", x"5e", x"61", x"5c", x"5a", x"5c", x"60", x"66", x"64", 
        x"3e", x"39", x"2d", x"42", x"ba", x"a4", x"34", x"31", x"2f", x"24", x"34", x"39", x"25", x"31", x"2c", 
        x"37", x"32", x"2a", x"83", x"cf", x"c2", x"c6", x"d8", x"c5", x"c6", x"d1", x"e4", x"e2", x"e1", x"e6", 
        x"e0", x"dd", x"e2", x"e4", x"e3", x"e3", x"e1", x"e0", x"e2", x"e0", x"dc", x"da", x"e1", x"e8", x"e0", 
        x"e7", x"e0", x"db", x"e8", x"db", x"d7", x"e3", x"e3", x"e4", x"e7", x"e2", x"e5", x"e5", x"e7", x"e7", 
        x"de", x"e1", x"e8", x"eb", x"e7", x"ea", x"ed", x"e9", x"e7", x"e8", x"e6", x"df", x"e1", x"e6", x"e3", 
        x"e1", x"e2", x"ca", x"ca", x"e6", x"e6", x"e3", x"e4", x"e5", x"e5", x"e7", x"e6", x"df", x"e5", x"e6", 
        x"e5", x"e8", x"e7", x"eb", x"ea", x"e7", x"e5", x"e6", x"e5", x"e5", x"e6", x"e9", x"ed", x"e6", x"e3", 
        x"e7", x"e3", x"e6", x"e8", x"df", x"e1", x"e4", x"e6", x"ec", x"e9", x"e8", x"e8", x"ea", x"ea", x"ea", 
        x"ec", x"e8", x"e6", x"e6", x"e8", x"ec", x"ec", x"e9", x"eb", x"eb", x"ea", x"e4", x"e8", x"f0", x"f2", 
        x"e9", x"e2", x"e1", x"e5", x"ec", x"eb", x"e8", x"eb", x"eb", x"ee", x"e6", x"de", x"e5", x"e4", x"e1", 
        x"e4", x"e9", x"e8", x"e8", x"e9", x"e9", x"e5", x"e9", x"e3", x"e7", x"e7", x"e2", x"e5", x"e6", x"e9", 
        x"ec", x"eb", x"ea", x"eb", x"e9", x"e9", x"e6", x"eb", x"e9", x"e8", x"ea", x"e8", x"e8", x"e9", x"e7", 
        x"e6", x"ee", x"e9", x"ee", x"ed", x"e5", x"ea", x"ea", x"ea", x"e8", x"ec", x"eb", x"eb", x"ed", x"e9", 
        x"e8", x"ea", x"ec", x"eb", x"eb", x"ea", x"eb", x"ec", x"ee", x"ec", x"ea", x"ee", x"e6", x"e4", x"ea", 
        x"e9", x"e6", x"e8", x"e9", x"e8", x"ea", x"eb", x"eb", x"ed", x"eb", x"ec", x"e9", x"e9", x"eb", x"e9", 
        x"ea", x"ee", x"e9", x"ed", x"ef", x"ef", x"ec", x"e9", x"e4", x"e4", x"e8", x"e6", x"ea", x"e7", x"e3", 
        x"e6", x"e8", x"e7", x"eb", x"e8", x"e8", x"ed", x"e3", x"e5", x"e9", x"ec", x"ea", x"e7", x"e7", x"e8", 
        x"eb", x"eb", x"eb", x"ed", x"ed", x"ed", x"ec", x"eb", x"ed", x"ea", x"e9", x"ea", x"e7", x"eb", x"f1", 
        x"ef", x"eb", x"ea", x"e9", x"ee", x"ec", x"ec", x"eb", x"ec", x"eb", x"e6", x"e8", x"eb", x"eb", x"ea", 
        x"eb", x"ed", x"ef", x"ef", x"ec", x"eb", x"ee", x"f0", x"ed", x"eb", x"ee", x"ed", x"eb", x"ed", x"eb", 
        x"ea", x"ee", x"e0", x"dc", x"e8", x"ea", x"ec", x"ee", x"e9", x"e8", x"ed", x"ed", x"eb", x"ec", x"ec", 
        x"eb", x"ea", x"ed", x"ee", x"eb", x"ea", x"ea", x"ea", x"e9", x"ec", x"ee", x"eb", x"e9", x"eb", x"ec", 
        x"ea", x"eb", x"ec", x"e9", x"e9", x"e6", x"e4", x"eb", x"ee", x"ee", x"ed", x"e8", x"e8", x"ee", x"ee", 
        x"ed", x"ec", x"ec", x"eb", x"eb", x"ea", x"ea", x"ec", x"ea", x"eb", x"eb", x"eb", x"e9", x"e7", x"ed", 
        x"ec", x"ea", x"ec", x"ee", x"ed", x"ed", x"ed", x"ed", x"f0", x"f0", x"ec", x"ec", x"ee", x"eb", x"e9", 
        x"eb", x"dd", x"e5", x"ee", x"f0", x"f2", x"f2", x"f2", x"f0", x"f0", x"f1", x"f1", x"f2", x"ef", x"ee", 
        x"f2", x"f1", x"ee", x"f0", x"f2", x"ec", x"ee", x"f2", x"f0", x"ee", x"ee", x"ee", x"ef", x"f0", x"ed", 
        x"ef", x"f0", x"f1", x"f1", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"f0", x"f1", x"f2", x"f3", x"f3", 
        x"f2", x"ef", x"ef", x"f0", x"f1", x"f3", x"f3", x"f0", x"f0", x"ef", x"ed", x"f0", x"ef", x"ee", x"ed", 
        x"ed", x"ef", x"ef", x"ef", x"e6", x"ec", x"f2", x"f1", x"f1", x"ef", x"ef", x"f0", x"ef", x"f1", x"f2", 
        x"ef", x"ee", x"ef", x"ee", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f0", x"f1", x"f4", x"f4", x"f4", 
        x"f2", x"f1", x"f2", x"ef", x"ee", x"f0", x"f0", x"f2", x"f6", x"f7", x"f4", x"f1", x"f0", x"f2", x"f1", 
        x"ef", x"ee", x"ed", x"ed", x"ef", x"f0", x"ee", x"ed", x"ed", x"ed", x"ef", x"ee", x"ee", x"e8", x"ed", 
        x"ee", x"ef", x"ed", x"ed", x"ee", x"ee", x"ec", x"ed", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"f0", 
        x"f2", x"f1", x"f0", x"f1", x"ef", x"f1", x"ef", x"ef", x"ef", x"ef", x"f2", x"f3", x"f1", x"ed", x"f0", 
        x"f1", x"ef", x"f0", x"f0", x"f1", x"ee", x"ef", x"ef", x"f1", x"da", x"81", x"6a", x"5c", x"4c", x"51", 
        x"6c", x"56", x"94", x"bb", x"ce", x"cb", x"c1", x"d8", x"ee", x"eb", x"ed", x"ea", x"f1", x"f0", x"ec", 
        x"ec", x"ef", x"ce", x"8b", x"b7", x"ce", x"d6", x"e0", x"cb", x"ce", x"e9", x"f3", x"f2", x"f3", x"f1", 
        x"ef", x"ef", x"f2", x"f1", x"f0", x"f0", x"f2", x"f0", x"f3", x"e9", x"64", x"44", x"90", x"de", x"d4", 
        x"d5", x"d3", x"da", x"d0", x"7f", x"c1", x"e2", x"c4", x"56", x"1e", x"14", x"15", x"1c", x"1d", x"50", 
        x"79", x"71", x"73", x"6a", x"4a", x"37", x"3a", x"3f", x"3d", x"3b", x"3d", x"42", x"3e", x"18", x"03", 
        x"08", x"07", x"15", x"62", x"d8", x"c5", x"43", x"12", x"0b", x"08", x"0d", x"15", x"17", x"28", x"62", 
        x"a3", x"97", x"36", x"0a", x"07", x"06", x"05", x"07", x"08", x"09", x"0a", x"1b", x"3f", x"53", x"67", 
        x"53", x"3a", x"27", x"3e", x"54", x"4a", x"48", x"4d", x"4a", x"4c", x"4b", x"3c", x"4e", x"6e", x"52", 
        x"30", x"1c", x"1a", x"2f", x"37", x"74", x"d3", x"5c", x"10", x"17", x"23", x"3c", x"48", x"73", x"af", 
        x"b7", x"b9", x"7f", x"35", x"3d", x"5a", x"5d", x"64", x"6a", x"68", x"77", x"76", x"75", x"7a", x"77", 
        x"58", x"23", x"2f", x"3c", x"4d", x"34", x"35", x"39", x"43", x"56", x"59", x"63", x"68", x"67", x"64", 
        x"57", x"4c", x"4e", x"4d", x"4b", x"42", x"39", x"3b", x"35", x"2f", x"2e", x"2f", x"24", x"23", x"21", 
        x"26", x"35", x"31", x"44", x"a3", x"83", x"3d", x"23", x"1f", x"20", x"20", x"1c", x"16", x"31", x"30", 
        x"2f", x"31", x"4b", x"ab", x"d1", x"c9", x"d2", x"dc", x"ca", x"c7", x"ce", x"e1", x"dd", x"dc", x"e4", 
        x"e3", x"df", x"dc", x"e2", x"e6", x"e0", x"dd", x"e1", x"e7", x"e5", x"e1", x"dd", x"e0", x"e6", x"e6", 
        x"ea", x"e8", x"e6", x"e6", x"de", x"de", x"e4", x"e6", x"e8", x"e5", x"e3", x"e7", x"e5", x"e6", x"e8", 
        x"e8", x"e4", x"e4", x"e9", x"e7", x"e6", x"ea", x"e6", x"e3", x"e7", x"e6", x"e1", x"e3", x"e8", x"e6", 
        x"e6", x"e9", x"ce", x"cc", x"e4", x"e2", x"e1", x"e5", x"e2", x"de", x"e1", x"e6", x"e6", x"e7", x"e6", 
        x"e7", x"e5", x"e6", x"e7", x"ea", x"e8", x"e3", x"e5", x"e2", x"e0", x"e4", x"e5", x"e6", x"e3", x"e3", 
        x"df", x"dd", x"e8", x"e5", x"df", x"e1", x"e7", x"e8", x"eb", x"ea", x"e9", x"ec", x"eb", x"ea", x"e7", 
        x"e4", x"e8", x"e9", x"e9", x"eb", x"eb", x"e8", x"e7", x"e9", x"eb", x"ee", x"eb", x"e9", x"e9", x"ea", 
        x"e8", x"e7", x"e6", x"e8", x"ec", x"e9", x"ea", x"eb", x"eb", x"eb", x"e9", x"e7", x"e8", x"e8", x"ea", 
        x"e9", x"ec", x"ea", x"e8", x"e8", x"e7", x"e2", x"e6", x"e4", x"e9", x"eb", x"e8", x"e9", x"e6", x"e7", 
        x"ea", x"ed", x"ef", x"ea", x"e4", x"e7", x"e5", x"e8", x"e5", x"e9", x"ed", x"e8", x"e7", x"ea", x"ea", 
        x"e8", x"ea", x"e3", x"ea", x"ec", x"e5", x"eb", x"e9", x"e9", x"e6", x"e7", x"eb", x"ea", x"ed", x"ed", 
        x"eb", x"e9", x"e9", x"e9", x"ec", x"ef", x"ea", x"e9", x"eb", x"eb", x"ec", x"ec", x"e4", x"e5", x"ee", 
        x"eb", x"e9", x"ec", x"ec", x"ea", x"ea", x"e9", x"e9", x"ef", x"ed", x"eb", x"e8", x"eb", x"ec", x"ea", 
        x"eb", x"ef", x"ec", x"eb", x"e7", x"e7", x"e4", x"e8", x"ea", x"eb", x"eb", x"ea", x"ee", x"ee", x"ea", 
        x"eb", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"eb", x"e6", x"e9", x"f2", x"ed", x"eb", x"ea", x"e8", 
        x"e9", x"e8", x"e9", x"ee", x"ed", x"ef", x"ed", x"eb", x"ee", x"eb", x"eb", x"ee", x"e8", x"e9", x"ee", 
        x"ec", x"eb", x"ec", x"e8", x"e9", x"eb", x"ed", x"eb", x"eb", x"ec", x"e9", x"ea", x"ec", x"eb", x"e9", 
        x"e9", x"ea", x"eb", x"ee", x"ed", x"eb", x"ec", x"ef", x"ef", x"ed", x"ea", x"ec", x"ed", x"e9", x"ea", 
        x"eb", x"eb", x"e0", x"dc", x"e9", x"ea", x"eb", x"ec", x"ea", x"eb", x"ed", x"ed", x"eb", x"eb", x"ec", 
        x"eb", x"ec", x"ec", x"ed", x"ed", x"eb", x"ea", x"eb", x"ed", x"ed", x"ea", x"e8", x"e9", x"eb", x"e9", 
        x"e9", x"ec", x"eb", x"ea", x"eb", x"eb", x"ec", x"ec", x"e7", x"e8", x"ed", x"ea", x"e6", x"ea", x"ec", 
        x"ed", x"ec", x"eb", x"ea", x"ea", x"ec", x"ed", x"ed", x"eb", x"ed", x"ed", x"ee", x"eb", x"e9", x"ee", 
        x"ed", x"ec", x"ee", x"ee", x"ed", x"ee", x"ef", x"ef", x"f0", x"ef", x"ec", x"ed", x"ee", x"ec", x"e9", 
        x"ec", x"e1", x"e7", x"ee", x"ec", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"f1", x"f0", x"ec", 
        x"ee", x"f1", x"f0", x"f0", x"f0", x"ed", x"ee", x"f1", x"f1", x"f1", x"ee", x"ed", x"ef", x"f0", x"ef", 
        x"f1", x"f1", x"f2", x"f1", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"f1", x"f2", x"f2", x"f3", x"f3", 
        x"f1", x"f0", x"f0", x"ef", x"ef", x"f2", x"f2", x"f1", x"f1", x"ee", x"ed", x"f1", x"f0", x"f1", x"f0", 
        x"ee", x"ee", x"ee", x"ef", x"e6", x"ea", x"f0", x"f0", x"f0", x"ee", x"ef", x"f0", x"ef", x"f0", x"f3", 
        x"ef", x"ef", x"f1", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f3", x"f4", x"f4", x"f3", 
        x"f2", x"f1", x"f1", x"ee", x"ef", x"f1", x"f2", x"f3", x"f7", x"f6", x"f3", x"f0", x"f0", x"f1", x"f1", 
        x"ef", x"f1", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"f0", x"ef", x"ee", x"e6", x"ec", 
        x"ef", x"f1", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", x"f1", x"f0", x"ef", x"ee", x"ed", x"ed", x"ee", 
        x"f2", x"f1", x"f0", x"f1", x"ef", x"f1", x"ef", x"ed", x"ef", x"f1", x"f2", x"f0", x"f0", x"ef", x"f0", 
        x"ee", x"ef", x"ef", x"f0", x"f2", x"f0", x"ef", x"ef", x"eb", x"a4", x"67", x"7c", x"6e", x"5f", x"5b", 
        x"77", x"63", x"8c", x"c1", x"c7", x"cb", x"b9", x"c1", x"eb", x"ee", x"ee", x"ea", x"ed", x"ed", x"ec", 
        x"ed", x"f4", x"d1", x"83", x"b1", x"ce", x"d3", x"d6", x"c2", x"ce", x"e6", x"f3", x"f2", x"f3", x"f1", 
        x"ee", x"ee", x"f0", x"ef", x"f0", x"f2", x"f4", x"ef", x"f1", x"e9", x"69", x"43", x"90", x"e4", x"d6", 
        x"d8", x"d7", x"d7", x"d0", x"82", x"bf", x"e1", x"c2", x"53", x"20", x"22", x"2e", x"46", x"47", x"60", 
        x"75", x"68", x"5c", x"5a", x"4a", x"44", x"49", x"45", x"46", x"4b", x"47", x"48", x"4d", x"35", x"0f", 
        x"04", x"0a", x"0c", x"46", x"cc", x"cc", x"57", x"14", x"17", x"36", x"1a", x"05", x"07", x"0b", x"12", 
        x"66", x"bf", x"86", x"1f", x"07", x"03", x"0b", x"0c", x"07", x"06", x"06", x"31", x"4f", x"40", x"3c", 
        x"3c", x"34", x"25", x"35", x"41", x"3d", x"41", x"46", x"49", x"48", x"47", x"46", x"5b", x"75", x"5a", 
        x"36", x"27", x"56", x"66", x"4d", x"59", x"bb", x"92", x"46", x"36", x"2f", x"22", x"2c", x"85", x"af", 
        x"b7", x"a4", x"3d", x"28", x"52", x"70", x"6b", x"66", x"69", x"69", x"5c", x"50", x"48", x"46", x"3c", 
        x"2c", x"1d", x"20", x"4a", x"6c", x"3e", x"62", x"7e", x"97", x"74", x"2d", x"1c", x"1b", x"1a", x"1b", 
        x"21", x"12", x"0f", x"0e", x"0e", x"10", x"11", x"12", x"0a", x"0b", x"18", x"21", x"12", x"0c", x"09", 
        x"21", x"2c", x"26", x"4f", x"b8", x"91", x"46", x"30", x"23", x"28", x"29", x"27", x"16", x"1c", x"29", 
        x"2d", x"2e", x"3e", x"99", x"d4", x"c8", x"d0", x"db", x"cb", x"c7", x"cf", x"e0", x"e0", x"e1", x"e0", 
        x"e7", x"e8", x"e3", x"e3", x"e6", x"e3", x"e3", x"e4", x"e5", x"e5", x"e2", x"e1", x"df", x"df", x"de", 
        x"e5", x"e5", x"e2", x"e4", x"e1", x"db", x"db", x"e1", x"e7", x"e8", x"e8", x"e6", x"e2", x"e9", x"ea", 
        x"ea", x"e7", x"e2", x"e3", x"e8", x"e8", x"e9", x"e7", x"e5", x"e6", x"e6", x"e5", x"e4", x"e5", x"e3", 
        x"e5", x"eb", x"e1", x"df", x"e5", x"e8", x"e8", x"e5", x"dd", x"de", x"e0", x"e4", x"e8", x"e4", x"e3", 
        x"e9", x"e9", x"e9", x"e5", x"eb", x"ea", x"e6", x"e8", x"e4", x"df", x"e5", x"e4", x"e5", x"e8", x"e3", 
        x"dc", x"e1", x"e9", x"e8", x"e3", x"e1", x"e3", x"e3", x"e8", x"ea", x"e7", x"ea", x"ea", x"e9", x"e7", 
        x"e4", x"eb", x"ea", x"ea", x"ea", x"ea", x"e7", x"e7", x"e5", x"e9", x"ed", x"ea", x"e9", x"ea", x"ec", 
        x"ec", x"ea", x"e8", x"e8", x"ea", x"e8", x"ec", x"ec", x"eb", x"e8", x"ea", x"ea", x"e9", x"e9", x"eb", 
        x"e9", x"ea", x"e7", x"e4", x"e6", x"e8", x"e6", x"ec", x"e8", x"ea", x"eb", x"e9", x"e9", x"e4", x"e3", 
        x"e7", x"ea", x"ed", x"ee", x"ec", x"ec", x"e7", x"e8", x"e8", x"ed", x"ef", x"e8", x"e5", x"e7", x"e6", 
        x"e4", x"e9", x"e5", x"ea", x"ea", x"e6", x"e9", x"ea", x"ed", x"e8", x"e6", x"ea", x"e7", x"ea", x"ed", 
        x"ed", x"ed", x"eb", x"e9", x"ec", x"ef", x"ec", x"ec", x"ee", x"ec", x"ec", x"ea", x"e9", x"ec", x"ee", 
        x"e6", x"e9", x"e9", x"e8", x"e6", x"e9", x"e8", x"e8", x"ee", x"ed", x"ea", x"e9", x"ea", x"eb", x"ed", 
        x"e9", x"e6", x"e3", x"eb", x"e9", x"e3", x"e3", x"e6", x"e7", x"ed", x"eb", x"e7", x"e3", x"e5", x"e5", 
        x"e6", x"ed", x"ef", x"ef", x"ee", x"ee", x"eb", x"eb", x"e8", x"e9", x"ec", x"eb", x"f0", x"ef", x"e9", 
        x"e7", x"e5", x"e8", x"ec", x"ea", x"ee", x"eb", x"eb", x"ef", x"ee", x"e9", x"e6", x"e8", x"e9", x"ea", 
        x"ea", x"eb", x"eb", x"eb", x"e9", x"ec", x"ed", x"ea", x"ea", x"eb", x"ec", x"ed", x"ed", x"eb", x"ea", 
        x"eb", x"ed", x"ed", x"ed", x"ed", x"eb", x"eb", x"ec", x"ef", x"ec", x"e6", x"ea", x"ec", x"e7", x"ea", 
        x"ee", x"ec", x"de", x"da", x"ea", x"ec", x"ea", x"ed", x"ec", x"eb", x"eb", x"ec", x"eb", x"ea", x"ed", 
        x"ec", x"ee", x"eb", x"ec", x"ed", x"ec", x"ea", x"eb", x"ef", x"ed", x"e9", x"e7", x"ea", x"ec", x"ea", 
        x"ec", x"ee", x"e6", x"e4", x"e9", x"ea", x"ec", x"ed", x"eb", x"ea", x"ed", x"ec", x"ed", x"ec", x"ea", 
        x"ee", x"ec", x"ea", x"eb", x"ec", x"ee", x"ed", x"eb", x"eb", x"ef", x"f0", x"f1", x"ec", x"e9", x"ee", 
        x"ec", x"ec", x"ed", x"ea", x"e8", x"ea", x"ee", x"ed", x"ee", x"ee", x"eb", x"ea", x"e8", x"ea", x"ec", 
        x"ed", x"e4", x"e8", x"f0", x"f0", x"f1", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f1", x"f0", x"ec", 
        x"ec", x"ef", x"f0", x"ef", x"ee", x"f1", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ef", x"ef", 
        x"f0", x"f0", x"ef", x"f0", x"ee", x"ed", x"ef", x"ee", x"ee", x"f0", x"f1", x"f3", x"f3", x"f4", x"f3", 
        x"f1", x"f0", x"ef", x"ee", x"ed", x"f1", x"f1", x"f2", x"f2", x"ef", x"ef", x"f1", x"ed", x"f0", x"f0", 
        x"ec", x"ed", x"ec", x"ef", x"e7", x"eb", x"f0", x"ef", x"f0", x"ee", x"ee", x"f0", x"ee", x"ec", x"f0", 
        x"ec", x"ee", x"f3", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"f0", x"f1", x"f3", x"f4", x"f3", x"f2", 
        x"f1", x"f1", x"f0", x"ef", x"f0", x"f2", x"f2", x"f3", x"f6", x"f6", x"f2", x"f0", x"f1", x"f1", x"f0", 
        x"ef", x"f0", x"f0", x"ef", x"ed", x"ee", x"ef", x"ed", x"ee", x"ef", x"ef", x"ef", x"ee", x"e6", x"eb", 
        x"ef", x"ef", x"ed", x"ef", x"ee", x"ef", x"ef", x"ed", x"ef", x"f0", x"ef", x"ef", x"ed", x"ed", x"ef", 
        x"f2", x"f1", x"f1", x"f2", x"f0", x"f2", x"f0", x"ed", x"ef", x"f3", x"f2", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"e5", x"88", x"68", x"82", x"7a", x"75", x"7a", 
        x"72", x"7f", x"6f", x"b0", x"bf", x"cb", x"b6", x"af", x"e3", x"ef", x"ed", x"f1", x"f2", x"ed", x"ec", 
        x"ec", x"ef", x"c9", x"85", x"b1", x"c8", x"d2", x"d5", x"c1", x"cf", x"e2", x"f2", x"f3", x"f4", x"f2", 
        x"ef", x"ef", x"f2", x"f2", x"f0", x"f1", x"f3", x"f0", x"f1", x"e9", x"6e", x"3a", x"86", x"db", x"ca", 
        x"ca", x"cd", x"ce", x"ca", x"7e", x"b5", x"e3", x"cc", x"93", x"5b", x"60", x"79", x"a5", x"ae", x"90", 
        x"6b", x"52", x"42", x"4d", x"4e", x"4f", x"4d", x"46", x"48", x"4f", x"47", x"45", x"49", x"47", x"24", 
        x"07", x"0b", x"0c", x"30", x"b7", x"d3", x"5f", x"0d", x"18", x"35", x"10", x"03", x"02", x"05", x"04", 
        x"1a", x"5f", x"97", x"3e", x"0b", x"0b", x"15", x"15", x"03", x"05", x"0a", x"1d", x"44", x"57", x"5b", 
        x"5e", x"60", x"67", x"78", x"7e", x"84", x"85", x"88", x"8a", x"89", x"81", x"7d", x"7f", x"80", x"61", 
        x"3b", x"2e", x"61", x"6b", x"4d", x"42", x"86", x"b8", x"6a", x"4c", x"3b", x"25", x"41", x"95", x"b5", 
        x"c5", x"97", x"24", x"23", x"22", x"1b", x"14", x"10", x"1d", x"28", x"16", x"0e", x"0b", x"12", x"18", 
        x"17", x"2b", x"2c", x"33", x"3f", x"40", x"b1", x"c5", x"c6", x"76", x"1d", x"18", x"1b", x"20", x"1f", 
        x"2c", x"15", x"0d", x"13", x"16", x"15", x"10", x"13", x"15", x"17", x"1e", x"27", x"1d", x"1c", x"1b", 
        x"16", x"1e", x"17", x"42", x"be", x"a5", x"3d", x"39", x"1b", x"1f", x"1e", x"1b", x"14", x"23", x"34", 
        x"45", x"32", x"26", x"83", x"d8", x"c1", x"c9", x"de", x"d0", x"c4", x"c8", x"d9", x"da", x"de", x"db", 
        x"df", x"e4", x"e2", x"e4", x"e7", x"e3", x"e4", x"e6", x"e3", x"e4", x"e2", x"e1", x"d9", x"cc", x"cd", 
        x"e3", x"e6", x"e3", x"e9", x"e4", x"e3", x"dc", x"d7", x"de", x"e5", x"e5", x"e0", x"e2", x"e8", x"e7", 
        x"ea", x"e4", x"e7", x"e9", x"e8", x"e9", x"e8", x"ea", x"e8", x"e6", x"e4", x"ea", x"eb", x"e9", x"e5", 
        x"e4", x"e6", x"e5", x"e1", x"e0", x"e5", x"e6", x"e0", x"d9", x"e3", x"e7", x"e9", x"e1", x"d8", x"e3", 
        x"e9", x"e6", x"e6", x"e3", x"e8", x"e8", x"e7", x"e8", x"e9", x"e5", x"e4", x"e2", x"e5", x"e7", x"e2", 
        x"e0", x"e3", x"e3", x"e7", x"e2", x"df", x"e3", x"e4", x"e7", x"ea", x"eb", x"eb", x"ea", x"e8", x"e7", 
        x"e7", x"e8", x"e5", x"e9", x"eb", x"e8", x"e4", x"ea", x"ea", x"ec", x"ea", x"e5", x"e9", x"ed", x"ed", 
        x"ea", x"e9", x"ea", x"ea", x"e9", x"e7", x"e8", x"e3", x"e7", x"ea", x"eb", x"e8", x"e8", x"eb", x"e7", 
        x"e8", x"ea", x"e9", x"e8", x"eb", x"ec", x"e7", x"e9", x"e9", x"e8", x"e8", x"e7", x"e9", x"e5", x"e5", 
        x"ec", x"e9", x"e5", x"eb", x"ea", x"e5", x"e1", x"e4", x"e5", x"e9", x"ec", x"e8", x"e8", x"ea", x"eb", 
        x"eb", x"ef", x"eb", x"eb", x"e9", x"e9", x"e7", x"e7", x"ee", x"eb", x"ea", x"eb", x"ea", x"e9", x"eb", 
        x"ee", x"f0", x"ee", x"ea", x"ea", x"eb", x"eb", x"ed", x"ed", x"eb", x"ed", x"e5", x"e4", x"ed", x"ee", 
        x"e5", x"ea", x"e8", x"e9", x"e7", x"e8", x"ea", x"ea", x"eb", x"e9", x"e9", x"eb", x"e8", x"e3", x"e9", 
        x"eb", x"e7", x"e2", x"ea", x"e7", x"df", x"e4", x"e5", x"e3", x"eb", x"eb", x"e9", x"e9", x"ea", x"ea", 
        x"e8", x"ec", x"eb", x"ec", x"eb", x"ea", x"eb", x"e7", x"e4", x"e9", x"ee", x"eb", x"ec", x"e9", x"e5", 
        x"ea", x"e9", x"ea", x"ed", x"ea", x"ee", x"eb", x"ec", x"f0", x"ef", x"e9", x"e5", x"e8", x"eb", x"ef", 
        x"ee", x"ee", x"ed", x"ef", x"eb", x"ec", x"ea", x"ea", x"ed", x"ec", x"ed", x"ed", x"ed", x"ec", x"eb", 
        x"ec", x"ed", x"ef", x"ed", x"ea", x"ea", x"eb", x"ec", x"ed", x"ea", x"e9", x"ec", x"eb", x"e9", x"eb", 
        x"ed", x"ef", x"e1", x"db", x"ec", x"ec", x"e8", x"e9", x"eb", x"e9", x"e7", x"ea", x"ea", x"e9", x"eb", 
        x"ea", x"ec", x"ea", x"ea", x"ea", x"ec", x"ec", x"ea", x"ed", x"ee", x"ed", x"eb", x"ec", x"ec", x"e9", 
        x"e9", x"ea", x"e4", x"e3", x"e7", x"e6", x"e7", x"ea", x"ed", x"ec", x"ec", x"eb", x"ed", x"eb", x"e8", 
        x"ec", x"ed", x"ec", x"eb", x"ea", x"eb", x"ec", x"ec", x"ea", x"ec", x"ec", x"ee", x"ee", x"ee", x"ed", 
        x"e8", x"e8", x"ec", x"eb", x"ea", x"ec", x"f0", x"ee", x"ed", x"ed", x"ec", x"ec", x"e9", x"ec", x"ed", 
        x"ec", x"e3", x"e7", x"f0", x"f2", x"f2", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ef", 
        x"ef", x"f1", x"ef", x"ed", x"f0", x"f1", x"f1", x"f2", x"f2", x"ee", x"ed", x"f1", x"ee", x"ef", x"f0", 
        x"f1", x"ef", x"ee", x"f0", x"ee", x"eb", x"ee", x"ee", x"ee", x"f1", x"f0", x"f3", x"f4", x"f5", x"f3", 
        x"f0", x"f0", x"ef", x"ed", x"ee", x"f1", x"f0", x"f1", x"f2", x"f0", x"f1", x"f0", x"ea", x"ee", x"ee", 
        x"eb", x"ee", x"ee", x"f1", x"e8", x"ec", x"f1", x"f0", x"f0", x"ef", x"ee", x"f1", x"ef", x"ee", x"f0", 
        x"ec", x"ed", x"f3", x"f0", x"ef", x"f1", x"f1", x"ef", x"ef", x"f0", x"f1", x"f2", x"f3", x"f1", x"f0", 
        x"f0", x"f0", x"f1", x"f0", x"f1", x"f1", x"ef", x"f2", x"f7", x"f6", x"f1", x"ef", x"f0", x"f0", x"ef", 
        x"ef", x"ed", x"ee", x"ee", x"ed", x"ee", x"ee", x"ea", x"ed", x"ef", x"ee", x"ef", x"ee", x"e5", x"eb", 
        x"ee", x"ec", x"ec", x"ee", x"ed", x"ee", x"ef", x"ed", x"f0", x"f1", x"f1", x"ef", x"ec", x"ec", x"ed", 
        x"f1", x"f0", x"f1", x"f2", x"f0", x"f3", x"f1", x"ef", x"f1", x"f2", x"f1", x"f1", x"f1", x"ed", x"ed", 
        x"ef", x"f1", x"f0", x"ee", x"ed", x"ef", x"ef", x"f0", x"e6", x"91", x"76", x"8a", x"8f", x"84", x"99", 
        x"7f", x"87", x"69", x"9b", x"bd", x"be", x"ae", x"a7", x"e2", x"ef", x"eb", x"ed", x"f0", x"f0", x"ec", 
        x"ef", x"ee", x"b8", x"7a", x"b1", x"c7", x"cd", x"d8", x"cd", x"d3", x"df", x"f1", x"f1", x"f1", x"ef", 
        x"eb", x"eb", x"ee", x"ee", x"ec", x"ee", x"ef", x"ec", x"ee", x"eb", x"79", x"3a", x"83", x"d4", x"c6", 
        x"c2", x"c5", x"c8", x"c4", x"86", x"aa", x"c2", x"a6", x"98", x"77", x"7d", x"af", x"b7", x"8e", x"6e", 
        x"5e", x"54", x"48", x"46", x"48", x"47", x"41", x"43", x"42", x"42", x"41", x"43", x"40", x"49", x"28", 
        x"07", x"07", x"0c", x"28", x"a9", x"d1", x"60", x"0d", x"10", x"15", x"05", x"02", x"01", x"04", x"07", 
        x"0a", x"46", x"af", x"65", x"10", x"0c", x"10", x"15", x"1a", x"35", x"35", x"2f", x"52", x"64", x"68", 
        x"64", x"62", x"5d", x"5a", x"51", x"48", x"40", x"49", x"41", x"3c", x"36", x"2d", x"36", x"6f", x"64", 
        x"40", x"1f", x"1c", x"1f", x"3e", x"52", x"51", x"75", x"37", x"16", x"13", x"1e", x"5b", x"9e", x"b7", 
        x"cf", x"87", x"21", x"32", x"25", x"0e", x"10", x"0c", x"1a", x"2c", x"1e", x"1d", x"23", x"22", x"1e", 
        x"1d", x"45", x"82", x"74", x"36", x"4e", x"ad", x"b1", x"bf", x"83", x"38", x"30", x"31", x"3e", x"3a", 
        x"43", x"38", x"3b", x"4a", x"4e", x"4a", x"41", x"42", x"4b", x"4f", x"4e", x"51", x"4f", x"53", x"4d", 
        x"1d", x"19", x"12", x"3d", x"ae", x"9b", x"38", x"43", x"24", x"19", x"1a", x"1f", x"28", x"30", x"3b", 
        x"46", x"2b", x"24", x"76", x"d2", x"c0", x"cc", x"e4", x"d7", x"c6", x"ca", x"dd", x"de", x"dd", x"da", 
        x"e1", x"e4", x"e1", x"e6", x"e5", x"d8", x"e1", x"e5", x"e4", x"e7", x"e3", x"e0", x"db", x"df", x"df", 
        x"e5", x"e4", x"e1", x"e5", x"e5", x"e9", x"e4", x"db", x"e3", x"eb", x"e3", x"e1", x"e6", x"e4", x"e2", 
        x"e7", x"e0", x"e4", x"e3", x"df", x"e5", x"e6", x"e9", x"e7", x"e6", x"e7", x"ea", x"e5", x"e4", x"e7", 
        x"e7", x"e3", x"e6", x"e4", x"e5", x"e2", x"e4", x"e2", x"de", x"e5", x"e7", x"ea", x"dd", x"d5", x"e5", 
        x"e8", x"e5", x"e8", x"e7", x"e9", x"e6", x"e4", x"e5", x"e7", x"e3", x"e2", x"e4", x"ea", x"e7", x"e7", 
        x"ea", x"eb", x"e7", x"e3", x"df", x"e1", x"e9", x"ea", x"e9", x"e7", x"eb", x"ea", x"e8", x"e6", x"e8", 
        x"e8", x"e7", x"e3", x"e7", x"ed", x"ee", x"e8", x"eb", x"ea", x"ea", x"e8", x"e4", x"e8", x"eb", x"e8", 
        x"e5", x"e9", x"ed", x"eb", x"ea", x"e9", x"ed", x"e9", x"ea", x"eb", x"ed", x"e8", x"e9", x"ea", x"e5", 
        x"e8", x"e7", x"e5", x"e4", x"e5", x"ea", x"e9", x"e9", x"ea", x"e9", x"e6", x"ea", x"ec", x"eb", x"ee", 
        x"ee", x"e9", x"e4", x"e8", x"e6", x"e2", x"e5", x"ea", x"e7", x"e7", x"e8", x"e5", x"e5", x"e6", x"e6", 
        x"e8", x"e7", x"e6", x"e9", x"eb", x"ec", x"ed", x"e9", x"ed", x"ed", x"ee", x"ea", x"e9", x"e8", x"eb", 
        x"ed", x"eb", x"e9", x"e7", x"e5", x"e5", x"e9", x"ea", x"eb", x"ec", x"ed", x"e4", x"e2", x"e8", x"eb", 
        x"e7", x"ec", x"ea", x"ec", x"e6", x"e7", x"ec", x"e8", x"e8", x"ea", x"e9", x"e9", x"e8", x"df", x"e3", 
        x"ec", x"ee", x"eb", x"eb", x"e7", x"e9", x"e9", x"ec", x"eb", x"ea", x"ea", x"ec", x"eb", x"ea", x"ea", 
        x"e9", x"ea", x"e9", x"ec", x"ea", x"e6", x"eb", x"ec", x"ec", x"ed", x"eb", x"eb", x"ee", x"ed", x"eb", 
        x"ef", x"ef", x"eb", x"ed", x"ed", x"ef", x"eb", x"ea", x"ee", x"ed", x"ea", x"ee", x"e9", x"ea", x"ee", 
        x"ec", x"e9", x"ea", x"ef", x"ec", x"eb", x"e9", x"ea", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ed", 
        x"eb", x"eb", x"ec", x"e8", x"e8", x"eb", x"ed", x"ee", x"ed", x"ec", x"ed", x"ee", x"eb", x"eb", x"ea", 
        x"ea", x"ec", x"df", x"da", x"eb", x"ef", x"eb", x"ec", x"ed", x"ec", x"ea", x"ec", x"ed", x"ec", x"ed", 
        x"eb", x"eb", x"e9", x"e8", x"e8", x"eb", x"eb", x"e9", x"ea", x"ef", x"f1", x"ef", x"ed", x"ec", x"eb", 
        x"e8", x"e9", x"e9", x"eb", x"ec", x"e9", x"ea", x"ec", x"eb", x"eb", x"ec", x"eb", x"ea", x"eb", x"e9", 
        x"ea", x"ee", x"ef", x"ec", x"e8", x"e8", x"ea", x"ea", x"e8", x"eb", x"ed", x"ef", x"ef", x"ee", x"ee", 
        x"eb", x"eb", x"ee", x"ef", x"ed", x"ed", x"ef", x"eb", x"e9", x"ea", x"eb", x"ed", x"ed", x"ec", x"ec", 
        x"ee", x"e7", x"e8", x"ef", x"ee", x"ee", x"ee", x"ef", x"ee", x"ec", x"ed", x"ed", x"ed", x"ef", x"f0", 
        x"ef", x"ee", x"ed", x"ec", x"ef", x"ef", x"f1", x"f4", x"f3", x"ee", x"ec", x"f0", x"ef", x"f1", x"f0", 
        x"f1", x"f0", x"ee", x"f0", x"ee", x"ec", x"f0", x"ef", x"ef", x"f1", x"f2", x"f4", x"f5", x"f6", x"f3", 
        x"f0", x"f0", x"ee", x"ee", x"f0", x"f2", x"f0", x"f1", x"f3", x"f0", x"f0", x"ee", x"eb", x"ee", x"ee", 
        x"eb", x"f0", x"f1", x"f2", x"e8", x"ed", x"ef", x"f0", x"f0", x"f1", x"ee", x"f1", x"f1", x"f0", x"f1", 
        x"ed", x"ee", x"f1", x"ee", x"ee", x"f0", x"f1", x"f0", x"ef", x"f1", x"f1", x"f2", x"f2", x"f0", x"ef", 
        x"f0", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", x"f3", x"f8", x"f4", x"f0", x"ef", x"f1", x"f0", x"ef", 
        x"f0", x"ee", x"ee", x"f0", x"f1", x"ef", x"f0", x"ed", x"ef", x"f0", x"ef", x"ee", x"ec", x"e7", x"ec", 
        x"ef", x"ef", x"ed", x"ef", x"ef", x"ef", x"f1", x"ee", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"f0", 
        x"f0", x"ef", x"f0", x"f0", x"f0", x"f3", x"f2", x"f0", x"f1", x"f0", x"f0", x"f2", x"f1", x"ec", x"ec", 
        x"ef", x"f1", x"f0", x"ee", x"ee", x"ef", x"f2", x"f2", x"da", x"89", x"83", x"91", x"a1", x"89", x"9d", 
        x"8c", x"78", x"71", x"7a", x"b8", x"ba", x"9f", x"a1", x"e1", x"f1", x"ef", x"eb", x"ec", x"ee", x"eb", 
        x"ea", x"ee", x"c1", x"87", x"b4", x"cd", x"cb", x"d0", x"cc", x"d5", x"dd", x"f0", x"ec", x"eb", x"e9", 
        x"e5", x"e4", x"e8", x"e7", x"e6", x"ec", x"e4", x"df", x"e8", x"e0", x"79", x"3c", x"68", x"9c", x"97", 
        x"8f", x"88", x"7f", x"77", x"58", x"5f", x"6b", x"56", x"4c", x"44", x"61", x"b3", x"a6", x"4a", x"32", 
        x"57", x"5e", x"61", x"60", x"64", x"68", x"6d", x"78", x"78", x"71", x"74", x"79", x"73", x"75", x"3a", 
        x"08", x"0a", x"19", x"48", x"b6", x"cf", x"6a", x"0e", x"05", x"05", x"04", x"03", x"01", x"03", x"08", 
        x"07", x"23", x"90", x"6b", x"13", x"05", x"07", x"1c", x"62", x"8e", x"7b", x"69", x"88", x"59", x"22", 
        x"1d", x"1a", x"18", x"1a", x"1e", x"15", x"15", x"2c", x"12", x"05", x"05", x"03", x"13", x"5c", x"61", 
        x"3b", x"1f", x"0e", x"0a", x"34", x"5b", x"52", x"68", x"39", x"23", x"17", x"2c", x"6f", x"98", x"b3", 
        x"d1", x"78", x"23", x"34", x"37", x"31", x"3a", x"3e", x"41", x"54", x"5c", x"62", x"6e", x"63", x"4e", 
        x"50", x"6d", x"aa", x"b7", x"67", x"50", x"b1", x"ab", x"bf", x"90", x"51", x"52", x"4d", x"49", x"46", 
        x"4b", x"49", x"47", x"41", x"3a", x"36", x"3b", x"3a", x"40", x"3c", x"32", x"30", x"30", x"2a", x"20", 
        x"15", x"12", x"0c", x"3b", x"a4", x"8f", x"2e", x"3b", x"47", x"23", x"2b", x"32", x"32", x"23", x"32", 
        x"3e", x"2b", x"1f", x"76", x"d7", x"c2", x"d3", x"e3", x"cd", x"c4", x"d2", x"e0", x"de", x"dc", x"e1", 
        x"e5", x"e3", x"de", x"e2", x"e5", x"e1", x"e3", x"e1", x"e1", x"e6", x"e3", x"d3", x"da", x"e4", x"df", 
        x"db", x"e5", x"e6", x"e1", x"e3", x"e2", x"ea", x"ec", x"ea", x"eb", x"e4", x"e7", x"ea", x"e5", x"e2", 
        x"e2", x"e6", x"e5", x"e3", x"e6", x"e5", x"e8", x"e8", x"e5", x"e9", x"eb", x"e5", x"e6", x"e6", x"e6", 
        x"e9", x"e3", x"e2", x"e4", x"e1", x"df", x"e5", x"e4", x"e6", x"e5", x"e1", x"e4", x"e9", x"e9", x"e6", 
        x"e6", x"e9", x"e9", x"e7", x"e6", x"e4", x"e2", x"e8", x"e8", x"e8", x"e8", x"e7", x"e8", x"e5", x"e8", 
        x"ea", x"ec", x"eb", x"e4", x"e2", x"e2", x"e6", x"e8", x"e9", x"e6", x"e8", x"e6", x"e2", x"e7", x"e9", 
        x"e6", x"eb", x"ed", x"e8", x"e6", x"ec", x"e9", x"ea", x"eb", x"ea", x"ee", x"ed", x"e8", x"e9", x"ea", 
        x"e7", x"ea", x"e9", x"eb", x"ec", x"ec", x"f0", x"ed", x"e8", x"e6", x"e5", x"e6", x"e6", x"e3", x"e6", 
        x"e7", x"e7", x"e8", x"e9", x"e5", x"e9", x"ed", x"ea", x"e9", x"e5", x"e2", x"eb", x"ea", x"e9", x"ea", 
        x"eb", x"ec", x"e8", x"e6", x"e8", x"e2", x"e3", x"e6", x"e7", x"e8", x"ea", x"e8", x"e9", x"e9", x"e7", 
        x"e8", x"e9", x"eb", x"ea", x"e9", x"de", x"ea", x"e9", x"e6", x"eb", x"eb", x"e8", x"eb", x"eb", x"ed", 
        x"ec", x"e6", x"e8", x"eb", x"e7", x"e6", x"ec", x"e9", x"ea", x"eb", x"e7", x"e9", x"ec", x"eb", x"e8", 
        x"e8", x"e9", x"e8", x"eb", x"e8", x"eb", x"eb", x"e3", x"e7", x"ee", x"e6", x"e1", x"ef", x"ee", x"ea", 
        x"ed", x"eb", x"eb", x"eb", x"ec", x"ea", x"e7", x"ec", x"ec", x"e7", x"e8", x"ea", x"eb", x"e8", x"e9", 
        x"ec", x"eb", x"ec", x"ee", x"ea", x"ea", x"ed", x"ee", x"ee", x"eb", x"e7", x"e9", x"ea", x"ec", x"e7", 
        x"e8", x"ee", x"ea", x"ed", x"ed", x"eb", x"ea", x"e9", x"eb", x"ea", x"e7", x"eb", x"e8", x"e8", x"e9", 
        x"ee", x"ed", x"ee", x"ef", x"ed", x"eb", x"ec", x"e9", x"ea", x"ed", x"ea", x"ed", x"ed", x"ee", x"f0", 
        x"ed", x"f0", x"ed", x"e7", x"ec", x"ed", x"ec", x"ed", x"ed", x"ed", x"eb", x"eb", x"ec", x"ec", x"ea", 
        x"e9", x"e9", x"e0", x"dd", x"e9", x"ee", x"ee", x"eb", x"e9", x"eb", x"eb", x"ea", x"eb", x"ea", x"ee", 
        x"ee", x"ed", x"eb", x"eb", x"eb", x"ea", x"e9", x"e9", x"e7", x"e9", x"eb", x"eb", x"eb", x"ec", x"ec", 
        x"ed", x"ea", x"ea", x"ea", x"ea", x"e8", x"eb", x"ec", x"eb", x"eb", x"ec", x"ec", x"ec", x"ed", x"ec", 
        x"eb", x"ed", x"ed", x"ec", x"ea", x"e9", x"ea", x"ef", x"ec", x"ed", x"ed", x"ec", x"ed", x"eb", x"eb", 
        x"ea", x"eb", x"ec", x"ec", x"ed", x"ed", x"ee", x"eb", x"ec", x"ee", x"ec", x"ed", x"ef", x"ec", x"eb", 
        x"f0", x"e7", x"e4", x"ef", x"ee", x"ef", x"ef", x"f1", x"ee", x"eb", x"ec", x"ee", x"ee", x"ee", x"ee", 
        x"ee", x"ea", x"ec", x"f0", x"ee", x"ee", x"ef", x"ef", x"ef", x"ee", x"ef", x"f1", x"ef", x"f1", x"ee", 
        x"ee", x"f1", x"ef", x"ef", x"ee", x"f0", x"f3", x"f2", x"f0", x"f1", x"f3", x"f6", x"f5", x"f5", x"f3", 
        x"ef", x"ef", x"ee", x"f0", x"f0", x"f1", x"f2", x"f3", x"f2", x"ef", x"ec", x"ed", x"ef", x"ef", x"ee", 
        x"ee", x"ef", x"ed", x"ef", x"e5", x"eb", x"eb", x"ef", x"ef", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ed", x"ee", x"ee", x"ec", x"ee", x"ee", x"ef", x"f2", x"f0", x"f3", x"f2", x"f2", x"f1", x"f0", x"f0", 
        x"f1", x"f2", x"f2", x"f1", x"f1", x"f2", x"f4", x"f6", x"f7", x"f2", x"f1", x"f1", x"f0", x"ef", x"f0", 
        x"f1", x"f2", x"ee", x"f1", x"f3", x"ed", x"f0", x"f2", x"ef", x"ee", x"ee", x"ec", x"ea", x"ec", x"ef", 
        x"f1", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f1", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", 
        x"f2", x"f0", x"f0", x"ef", x"f0", x"f5", x"f4", x"ef", x"ee", x"f0", x"f1", x"f1", x"f1", x"ef", x"f0", 
        x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"f3", x"da", x"8c", x"90", x"95", x"b5", x"95", x"95", 
        x"95", x"7b", x"7b", x"67", x"a6", x"c2", x"9e", x"a0", x"ce", x"ef", x"ee", x"eb", x"ec", x"ec", x"eb", 
        x"eb", x"f0", x"bd", x"83", x"ae", x"c4", x"cf", x"cb", x"c9", x"d3", x"de", x"f1", x"f1", x"f0", x"f1", 
        x"ee", x"ea", x"ec", x"e7", x"e0", x"e2", x"d6", x"d3", x"be", x"7d", x"38", x"21", x"28", x"3c", x"65", 
        x"6c", x"50", x"16", x"09", x"08", x"10", x"36", x"5d", x"73", x"37", x"3f", x"7d", x"5b", x"27", x"2a", 
        x"62", x"6d", x"66", x"62", x"60", x"54", x"50", x"49", x"49", x"46", x"43", x"44", x"42", x"3d", x"1a", 
        x"06", x"03", x"1a", x"79", x"d8", x"d1", x"7e", x"16", x"04", x"05", x"06", x"03", x"01", x"02", x"04", 
        x"05", x"25", x"9f", x"8f", x"22", x"28", x"55", x"8e", x"b7", x"af", x"a8", x"8c", x"a3", x"bd", x"76", 
        x"35", x"20", x"1f", x"22", x"27", x"28", x"2c", x"47", x"37", x"2e", x"33", x"36", x"3c", x"51", x"44", 
        x"30", x"2c", x"37", x"3f", x"48", x"4f", x"5a", x"71", x"5e", x"4b", x"42", x"4b", x"75", x"88", x"aa", 
        x"c9", x"5d", x"23", x"30", x"4a", x"5e", x"5d", x"50", x"3d", x"40", x"46", x"41", x"40", x"3f", x"36", 
        x"2e", x"55", x"98", x"b1", x"9c", x"4c", x"aa", x"b2", x"c3", x"8d", x"2a", x"15", x"16", x"13", x"10", 
        x"0e", x"10", x"14", x"0e", x"0d", x"11", x"12", x"1c", x"2c", x"27", x"25", x"27", x"22", x"1d", x"1f", 
        x"18", x"1b", x"11", x"55", x"cf", x"99", x"2a", x"30", x"4a", x"32", x"2f", x"24", x"1f", x"19", x"25", 
        x"2f", x"36", x"24", x"87", x"dd", x"cd", x"d3", x"e0", x"cc", x"c4", x"d0", x"df", x"dd", x"de", x"e4", 
        x"e3", x"df", x"e3", x"e1", x"dd", x"e4", x"e2", x"dd", x"e0", x"e7", x"e3", x"c9", x"d6", x"e7", x"e1", 
        x"df", x"e4", x"e5", x"e2", x"e4", x"dd", x"e1", x"e6", x"e3", x"e5", x"e6", x"e7", x"e7", x"e6", x"e2", 
        x"e2", x"e5", x"e3", x"e6", x"e7", x"e4", x"e5", x"e9", x"e8", x"ea", x"e9", x"e2", x"e7", x"e9", x"e3", 
        x"e5", x"e2", x"df", x"e3", x"e0", x"e5", x"e2", x"e4", x"e4", x"e0", x"e3", x"dc", x"e1", x"e5", x"e2", 
        x"e3", x"e7", x"e6", x"e8", x"e6", x"e4", x"e6", x"e7", x"e6", x"e7", x"e9", x"e6", x"e4", x"e5", x"e6", 
        x"e6", x"e9", x"e8", x"e5", x"e8", x"e5", x"e7", x"e7", x"e5", x"e5", x"e3", x"df", x"e2", x"ea", x"e8", 
        x"e6", x"e9", x"ea", x"e7", x"e7", x"e9", x"e6", x"e8", x"ec", x"e8", x"eb", x"eb", x"e6", x"e7", x"e9", 
        x"ea", x"ea", x"e7", x"ea", x"eb", x"eb", x"ef", x"ec", x"e8", x"e8", x"e6", x"e8", x"eb", x"e9", x"e7", 
        x"e5", x"e9", x"ee", x"eb", x"e5", x"e6", x"e6", x"ec", x"e9", x"e5", x"e1", x"e8", x"e8", x"e5", x"e2", 
        x"e8", x"eb", x"e7", x"e3", x"e6", x"e6", x"e4", x"e5", x"e6", x"e7", x"e9", x"e7", x"e9", x"ec", x"ea", 
        x"ea", x"ec", x"ec", x"ea", x"e8", x"e0", x"e9", x"e8", x"e6", x"ed", x"e8", x"ea", x"ed", x"ea", x"ed", 
        x"eb", x"e6", x"e8", x"eb", x"eb", x"ed", x"ee", x"eb", x"e9", x"e7", x"e5", x"e8", x"ea", x"ea", x"e8", 
        x"e9", x"ea", x"e9", x"eb", x"e7", x"ea", x"eb", x"e6", x"e7", x"e9", x"e3", x"e1", x"ed", x"ec", x"e9", 
        x"eb", x"ea", x"eb", x"eb", x"eb", x"eb", x"ea", x"eb", x"e9", x"e9", x"ed", x"ee", x"ef", x"ea", x"eb", 
        x"ed", x"ec", x"ee", x"ee", x"eb", x"ea", x"eb", x"eb", x"eb", x"eb", x"ea", x"ea", x"ea", x"ef", x"ec", 
        x"eb", x"ee", x"eb", x"ea", x"ea", x"eb", x"ea", x"ec", x"ec", x"e8", x"e9", x"ec", x"eb", x"ec", x"ec", 
        x"ed", x"ec", x"ec", x"ec", x"ed", x"ea", x"ea", x"ea", x"ee", x"ed", x"eb", x"eb", x"ea", x"eb", x"ea", 
        x"eb", x"ee", x"ee", x"ea", x"ed", x"ed", x"ec", x"ea", x"ea", x"ea", x"e8", x"ea", x"ec", x"eb", x"eb", 
        x"eb", x"eb", x"e2", x"de", x"e8", x"ec", x"ec", x"ea", x"e9", x"ee", x"ee", x"eb", x"ea", x"e9", x"ea", 
        x"ea", x"ed", x"ed", x"eb", x"ea", x"eb", x"ec", x"ea", x"e8", x"e9", x"ea", x"ea", x"ea", x"eb", x"ed", 
        x"ed", x"ea", x"ea", x"ea", x"ec", x"ea", x"ee", x"ed", x"eb", x"eb", x"eb", x"ec", x"ed", x"ed", x"ee", 
        x"ee", x"ee", x"ec", x"ec", x"ec", x"ec", x"ed", x"ef", x"ee", x"ec", x"ec", x"ec", x"ec", x"ec", x"ec", 
        x"eb", x"ea", x"ea", x"eb", x"ed", x"ee", x"ed", x"eb", x"ee", x"ef", x"eb", x"eb", x"ed", x"ec", x"eb", 
        x"ee", x"e5", x"e2", x"ed", x"ed", x"ee", x"ec", x"ee", x"ee", x"ee", x"f0", x"f1", x"f0", x"f1", x"f0", 
        x"f0", x"ed", x"ef", x"f2", x"f0", x"ef", x"ed", x"ed", x"ef", x"ef", x"ef", x"f1", x"ef", x"f0", x"f0", 
        x"f1", x"f2", x"f1", x"f1", x"f1", x"f2", x"f3", x"f0", x"ee", x"f0", x"f2", x"f5", x"f6", x"f6", x"f3", 
        x"ef", x"ef", x"ee", x"f0", x"f0", x"f0", x"f1", x"f2", x"f1", x"ef", x"ee", x"ef", x"ef", x"ed", x"ed", 
        x"ef", x"f0", x"ec", x"eb", x"e5", x"ed", x"ee", x"ef", x"ed", x"ee", x"ef", x"ee", x"ef", x"f0", x"ef", 
        x"ee", x"ed", x"ed", x"ec", x"ee", x"ee", x"ee", x"f1", x"ef", x"f1", x"f1", x"f2", x"f1", x"f0", x"ef", 
        x"f1", x"f2", x"f5", x"f3", x"f1", x"f2", x"f2", x"f5", x"f6", x"f1", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"f0", x"f2", x"ef", x"f1", x"f2", x"ed", x"f0", x"f1", x"ee", x"ee", x"ee", x"ec", x"eb", x"eb", x"ed", 
        x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"ef", x"ef", 
        x"f0", x"ef", x"f0", x"f1", x"f3", x"f7", x"f4", x"f0", x"ef", x"f0", x"f1", x"f1", x"f0", x"ee", x"ef", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", x"f1", x"e3", x"98", x"94", x"a3", x"bb", x"9c", x"9d", 
        x"a4", x"7e", x"84", x"61", x"8d", x"c5", x"ab", x"a5", x"ce", x"f1", x"ee", x"ea", x"ed", x"ec", x"ec", 
        x"ec", x"e4", x"b1", x"7c", x"a9", x"c3", x"cf", x"cb", x"ca", x"ce", x"d4", x"ca", x"c4", x"c0", x"bb", 
        x"b8", x"af", x"a7", x"9e", x"94", x"91", x"89", x"88", x"59", x"20", x"14", x"14", x"2a", x"66", x"6d", 
        x"60", x"3f", x"0f", x"05", x"08", x"04", x"0a", x"2a", x"54", x"28", x"1d", x"29", x"20", x"19", x"16", 
        x"1b", x"1c", x"1f", x"2a", x"30", x"1a", x"16", x"15", x"12", x"14", x"12", x"10", x"12", x"0c", x"05", 
        x"07", x"03", x"10", x"53", x"a2", x"82", x"45", x"0d", x"05", x"08", x"07", x"03", x"02", x"01", x"04", 
        x"06", x"29", x"9e", x"97", x"48", x"83", x"bd", x"d6", x"d3", x"ca", x"c6", x"a0", x"92", x"c6", x"c6", 
        x"6e", x"38", x"40", x"46", x"45", x"4c", x"4f", x"59", x"56", x"4d", x"4d", x"55", x"53", x"49", x"3c", 
        x"32", x"2f", x"39", x"3f", x"3a", x"49", x"65", x"6c", x"62", x"3b", x"2c", x"44", x"7e", x"7e", x"a3", 
        x"c3", x"4c", x"23", x"30", x"32", x"31", x"21", x"16", x"0f", x"12", x"18", x"1e", x"1d", x"1b", x"12", 
        x"14", x"4a", x"92", x"a2", x"af", x"5a", x"a3", x"b0", x"c3", x"92", x"2a", x"0d", x"10", x"0e", x"0e", 
        x"0f", x"15", x"1a", x"15", x"11", x"1b", x"23", x"3d", x"52", x"3b", x"38", x"3c", x"3c", x"40", x"42", 
        x"2a", x"2a", x"1b", x"51", x"cd", x"a1", x"2b", x"15", x"34", x"2d", x"23", x"1a", x"22", x"27", x"25", 
        x"38", x"3c", x"27", x"78", x"d1", x"c7", x"c8", x"dd", x"cf", x"c2", x"c9", x"e0", x"de", x"df", x"e1", 
        x"dd", x"d9", x"e3", x"de", x"d6", x"e5", x"e5", x"dd", x"e2", x"e4", x"e6", x"d8", x"df", x"e8", x"e1", 
        x"e5", x"e5", x"e7", x"e1", x"e1", x"e1", x"e4", x"e8", x"e3", x"e1", x"e7", x"e8", x"e6", x"e8", x"e3", 
        x"e3", x"e5", x"e1", x"e5", x"e5", x"e6", x"e7", x"ec", x"e8", x"e6", x"e9", x"e4", x"e3", x"e9", x"e5", 
        x"e4", x"e2", x"e0", x"e6", x"e2", x"e2", x"d9", x"e0", x"d2", x"cc", x"e2", x"df", x"e3", x"e7", x"e4", 
        x"e4", x"e7", x"e6", x"e9", x"e6", x"e5", x"e7", x"e6", x"e3", x"e3", x"e8", x"e8", x"e8", x"e9", x"e5", 
        x"e4", x"eb", x"eb", x"e4", x"e7", x"e9", x"ea", x"e9", x"e9", x"e3", x"e6", x"e3", x"e7", x"ea", x"e4", 
        x"e4", x"e7", x"e8", x"e8", x"e8", x"e9", x"e5", x"e6", x"e9", x"e9", x"ea", x"e8", x"ea", x"ea", x"e6", 
        x"e8", x"ea", x"ea", x"eb", x"e7", x"e5", x"e9", x"e8", x"e8", x"ee", x"eb", x"ea", x"eb", x"ea", x"eb", 
        x"e9", x"e8", x"ee", x"ec", x"e7", x"e5", x"e4", x"ef", x"e9", x"e9", x"ea", x"ec", x"eb", x"e9", x"e5", 
        x"ea", x"ea", x"ea", x"e5", x"e5", x"ea", x"e9", x"e9", x"e9", x"eb", x"ea", x"e4", x"e5", x"e9", x"e7", 
        x"e6", x"eb", x"e9", x"ec", x"eb", x"e9", x"eb", x"ea", x"eb", x"ed", x"ea", x"ed", x"e8", x"e8", x"ec", 
        x"ef", x"eb", x"e8", x"eb", x"ec", x"eb", x"ec", x"ea", x"e9", x"e9", x"eb", x"eb", x"e7", x"e6", x"e7", 
        x"e9", x"ea", x"ea", x"e8", x"e2", x"e9", x"ed", x"ea", x"eb", x"e9", x"e8", x"ea", x"ef", x"ed", x"e9", 
        x"ea", x"ea", x"e9", x"e7", x"e7", x"e9", x"e7", x"e8", x"e9", x"ec", x"ec", x"e9", x"ec", x"e7", x"e8", 
        x"ea", x"e9", x"ea", x"eb", x"ed", x"ed", x"ec", x"ea", x"eb", x"ec", x"ee", x"ec", x"e8", x"eb", x"ea", 
        x"ec", x"ed", x"e8", x"e4", x"e3", x"e7", x"e7", x"ec", x"ed", x"e9", x"ea", x"eb", x"eb", x"ec", x"ec", 
        x"ec", x"ea", x"e9", x"ec", x"f0", x"ec", x"e9", x"ef", x"f1", x"eb", x"ed", x"eb", x"ec", x"eb", x"e9", 
        x"eb", x"ed", x"ec", x"eb", x"ed", x"ee", x"ed", x"e9", x"e8", x"e8", x"e8", x"eb", x"ec", x"ea", x"ea", 
        x"eb", x"ec", x"e4", x"db", x"e5", x"ed", x"ec", x"e4", x"e2", x"ee", x"ef", x"ed", x"ed", x"eb", x"ed", 
        x"ed", x"ee", x"ed", x"e9", x"e7", x"e8", x"e9", x"e7", x"e9", x"ea", x"e9", x"e8", x"e8", x"eb", x"ef", 
        x"ee", x"e9", x"e8", x"e8", x"ec", x"eb", x"ee", x"ec", x"ec", x"ec", x"ec", x"ec", x"eb", x"eb", x"ec", 
        x"ef", x"ed", x"eb", x"eb", x"ed", x"ee", x"ef", x"f1", x"ef", x"ea", x"eb", x"ee", x"ec", x"eb", x"ea", 
        x"ea", x"eb", x"ed", x"ed", x"ed", x"ec", x"ec", x"eb", x"ea", x"eb", x"eb", x"ed", x"ed", x"ed", x"ec", 
        x"ef", x"e7", x"e4", x"ee", x"ef", x"f0", x"ed", x"ec", x"eb", x"ec", x"f0", x"f0", x"ee", x"f0", x"ef", 
        x"ef", x"ed", x"ee", x"f0", x"f0", x"ee", x"ec", x"ee", x"f2", x"f2", x"ef", x"ef", x"ee", x"f0", x"f2", 
        x"f2", x"f2", x"f1", x"f3", x"f2", x"f1", x"f1", x"ee", x"ee", x"f2", x"f4", x"f6", x"f6", x"f7", x"f4", 
        x"f0", x"f0", x"ef", x"f0", x"ee", x"ef", x"f0", x"f0", x"f0", x"f0", x"f0", x"ee", x"ef", x"ee", x"ed", 
        x"ed", x"f0", x"ef", x"eb", x"e6", x"ee", x"f0", x"f0", x"ee", x"ee", x"ed", x"ec", x"ed", x"ef", x"f1", 
        x"f0", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"f1", 
        x"f4", x"f6", x"f7", x"f5", x"f2", x"f1", x"f2", x"f4", x"f4", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", 
        x"f0", x"f1", x"ee", x"f0", x"f1", x"ed", x"f0", x"f1", x"ef", x"ee", x"ee", x"ec", x"ec", x"ea", x"ea", 
        x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"ed", x"ee", x"ef", x"f0", x"f0", x"ef", 
        x"ed", x"ed", x"ef", x"f1", x"f3", x"f5", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"ee", x"ed", x"ee", 
        x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ed", x"ef", x"ed", x"a4", x"87", x"b3", x"bb", x"94", x"93", 
        x"ac", x"7c", x"82", x"6a", x"7d", x"c3", x"ba", x"b6", x"db", x"ef", x"ea", x"ee", x"dd", x"ac", x"95", 
        x"85", x"81", x"78", x"74", x"a9", x"cb", x"cf", x"c7", x"cd", x"d4", x"bf", x"6a", x"3c", x"39", x"35", 
        x"37", x"36", x"31", x"2e", x"29", x"26", x"2a", x"2b", x"15", x"0f", x"18", x"1d", x"39", x"8c", x"59", 
        x"23", x"0e", x"06", x"05", x"05", x"03", x"0f", x"18", x"14", x"1b", x"50", x"5e", x"3c", x"1c", x"11", 
        x"0e", x"08", x"14", x"27", x"32", x"1e", x"21", x"2c", x"2c", x"32", x"32", x"2f", x"2e", x"10", x"02", 
        x"05", x"03", x"09", x"15", x"2c", x"18", x"06", x"05", x"08", x"05", x"03", x"03", x"05", x"03", x"09", 
        x"08", x"26", x"8b", x"89", x"80", x"b6", x"c5", x"c8", x"cb", x"cf", x"cb", x"ab", x"90", x"b2", x"db", 
        x"9e", x"3d", x"27", x"2c", x"28", x"27", x"28", x"24", x"22", x"1d", x"1f", x"1d", x"29", x"61", x"5a", 
        x"39", x"24", x"18", x"13", x"0f", x"22", x"4c", x"70", x"6f", x"2d", x"07", x"31", x"7e", x"85", x"a7", 
        x"c6", x"48", x"25", x"35", x"32", x"27", x"17", x"0d", x"0f", x"13", x"16", x"22", x"21", x"21", x"22", 
        x"28", x"50", x"71", x"80", x"b4", x"7f", x"83", x"8a", x"b0", x"a4", x"4f", x"41", x"49", x"46", x"50", 
        x"54", x"58", x"5b", x"56", x"4b", x"53", x"61", x"6d", x"72", x"5b", x"5d", x"5e", x"5e", x"5e", x"59", 
        x"3f", x"44", x"30", x"57", x"c5", x"9d", x"26", x"14", x"35", x"3d", x"27", x"1b", x"1d", x"17", x"1a", 
        x"40", x"2c", x"1e", x"7f", x"d8", x"cc", x"ca", x"dd", x"d1", x"c3", x"cc", x"e5", x"df", x"dd", x"e2", 
        x"e0", x"df", x"e6", x"e5", x"e1", x"e7", x"e1", x"de", x"e2", x"e1", x"e5", x"e3", x"e1", x"e3", x"dd", 
        x"e4", x"e1", x"e5", x"e3", x"e3", x"dc", x"dd", x"e6", x"e6", x"e2", x"e5", x"e6", x"e3", x"e6", x"e4", 
        x"e6", x"e5", x"e2", x"e6", x"e6", x"ea", x"e4", x"e5", x"e5", x"e5", x"e4", x"e0", x"e1", x"e2", x"e6", 
        x"e5", x"e5", x"e7", x"e6", x"e2", x"e3", x"df", x"e4", x"d2", x"cf", x"e3", x"e9", x"ea", x"e9", x"e6", 
        x"e3", x"e4", x"e7", x"e3", x"e1", x"e1", x"e0", x"e4", x"e2", x"df", x"dc", x"da", x"e2", x"e2", x"e2", 
        x"df", x"de", x"e6", x"e9", x"e7", x"e8", x"e8", x"ea", x"ed", x"e6", x"e8", x"e9", x"e9", x"eb", x"ea", 
        x"e7", x"e7", x"e6", x"e8", x"eb", x"ed", x"ec", x"e9", x"e3", x"e6", x"ee", x"ec", x"ea", x"e7", x"e3", 
        x"e4", x"e2", x"e5", x"e9", x"e8", x"e9", x"ec", x"eb", x"eb", x"ee", x"ea", x"e6", x"e6", x"eb", x"ed", 
        x"ec", x"e7", x"e7", x"ec", x"e9", x"e8", x"ea", x"ef", x"e8", x"ea", x"ed", x"eb", x"eb", x"eb", x"e8", 
        x"ea", x"e6", x"ed", x"ee", x"e7", x"e6", x"ea", x"eb", x"e8", x"ec", x"ec", x"e5", x"e5", x"e7", x"e8", 
        x"e7", x"ec", x"e9", x"ea", x"eb", x"ed", x"ec", x"ed", x"ec", x"e6", x"e7", x"e8", x"e8", x"ec", x"eb", 
        x"e9", x"ea", x"eb", x"e9", x"e9", x"eb", x"ed", x"ec", x"e9", x"e9", x"ea", x"e9", x"e9", x"eb", x"ea", 
        x"e9", x"e9", x"e9", x"ec", x"e7", x"ea", x"ea", x"e5", x"e5", x"e4", x"e7", x"e8", x"e9", x"eb", x"e9", 
        x"e9", x"ea", x"e7", x"e5", x"e5", x"e6", x"e9", x"eb", x"ec", x"e9", x"e7", x"e7", x"ed", x"ea", x"ec", 
        x"ee", x"ed", x"ee", x"ee", x"ed", x"ec", x"ec", x"e9", x"e8", x"e9", x"eb", x"ed", x"eb", x"ea", x"ea", 
        x"ed", x"ee", x"ea", x"e8", x"e6", x"e9", x"ea", x"ea", x"ed", x"ed", x"eb", x"ea", x"e8", x"e8", x"ec", 
        x"ed", x"eb", x"e9", x"ec", x"f0", x"ef", x"f0", x"f1", x"ed", x"ed", x"eb", x"e8", x"ea", x"ec", x"eb", 
        x"ed", x"ed", x"ec", x"e9", x"e6", x"e7", x"e8", x"e8", x"eb", x"ea", x"e9", x"ed", x"ec", x"e9", x"e9", 
        x"e9", x"ea", x"e3", x"d9", x"e4", x"ee", x"ee", x"e5", x"e1", x"eb", x"ed", x"ea", x"eb", x"eb", x"ed", 
        x"ed", x"eb", x"ea", x"ea", x"eb", x"eb", x"e9", x"e9", x"ea", x"ea", x"ea", x"e9", x"e8", x"eb", x"ee", 
        x"ee", x"ea", x"ea", x"e8", x"eb", x"eb", x"eb", x"ea", x"ea", x"ea", x"eb", x"eb", x"ec", x"ed", x"ed", 
        x"ed", x"eb", x"ea", x"ec", x"ed", x"ed", x"ed", x"ee", x"ef", x"eb", x"eb", x"ed", x"ec", x"ed", x"ed", 
        x"ec", x"ea", x"ea", x"ea", x"ec", x"ed", x"ec", x"ea", x"e8", x"e8", x"e9", x"e9", x"e6", x"ea", x"ee", 
        x"f1", x"e7", x"e2", x"ed", x"f0", x"f2", x"ee", x"ed", x"eb", x"ec", x"ef", x"ee", x"ea", x"ee", x"ee", 
        x"ed", x"ed", x"ee", x"ed", x"ef", x"f0", x"ed", x"ed", x"ef", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", 
        x"f0", x"ee", x"ef", x"f2", x"f2", x"f2", x"f1", x"ee", x"ee", x"f2", x"f5", x"f6", x"f6", x"f7", x"f4", 
        x"f0", x"f0", x"ef", x"f0", x"ee", x"ef", x"ef", x"ef", x"ef", x"f1", x"f2", x"f0", x"f2", x"f1", x"ed", 
        x"eb", x"ec", x"ec", x"ed", x"e7", x"ea", x"f0", x"f1", x"ef", x"ef", x"f1", x"f1", x"ef", x"ee", x"ef", 
        x"ed", x"eb", x"ec", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"f1", x"f4", x"f7", x"f4", x"f1", x"f1", x"f3", x"f4", x"f4", x"f0", x"f0", x"f0", x"ef", x"ee", x"ee", 
        x"ef", x"ef", x"ee", x"ee", x"ef", x"ee", x"f1", x"f2", x"ef", x"ef", x"ee", x"ed", x"ed", x"e9", x"e8", 
        x"ed", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ef", x"f0", x"ef", x"ef", 
        x"f1", x"ef", x"f0", x"f2", x"f4", x"f6", x"f2", x"f0", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ef", 
        x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"ee", x"f0", x"c1", x"8f", x"a9", x"c2", x"95", x"79", 
        x"98", x"75", x"70", x"6c", x"7c", x"b9", x"b4", x"b0", x"cc", x"ec", x"ec", x"dd", x"79", x"34", x"2c", 
        x"28", x"2f", x"4d", x"71", x"a4", x"c8", x"d4", x"c6", x"d0", x"e0", x"d2", x"70", x"18", x"1d", x"1f", 
        x"1f", x"1c", x"19", x"1a", x"1f", x"1e", x"1b", x"23", x"16", x"09", x"20", x"5b", x"77", x"a4", x"59", 
        x"1e", x"10", x"07", x"07", x"06", x"07", x"0b", x"13", x"0e", x"13", x"63", x"b5", x"a9", x"56", x"12", 
        x"10", x"0d", x"18", x"4d", x"63", x"59", x"5c", x"60", x"60", x"5e", x"5b", x"50", x"48", x"1e", x"06", 
        x"03", x"01", x"04", x"06", x"04", x"04", x"04", x"04", x"04", x"03", x"03", x"02", x"02", x"03", x"07", 
        x"07", x"21", x"8d", x"8c", x"99", x"ad", x"a9", x"b8", x"c9", x"cb", x"d0", x"b7", x"8f", x"9e", x"d5", 
        x"c0", x"49", x"05", x"09", x"0f", x"0d", x"0a", x"0d", x"0d", x"0b", x"0c", x"0d", x"32", x"6b", x"48", 
        x"33", x"2c", x"1e", x"1b", x"1f", x"20", x"2a", x"49", x"75", x"46", x"07", x"30", x"72", x"90", x"a2", 
        x"a9", x"42", x"28", x"2f", x"49", x"6a", x"5e", x"4d", x"4f", x"52", x"55", x"5e", x"5d", x"60", x"6b", 
        x"67", x"6d", x"89", x"97", x"9f", x"9d", x"8b", x"7c", x"a0", x"af", x"5f", x"4b", x"54", x"53", x"54", 
        x"50", x"4c", x"4a", x"49", x"3d", x"3c", x"37", x"2d", x"29", x"2d", x"2a", x"22", x"1f", x"1e", x"19", 
        x"4d", x"56", x"29", x"4a", x"b5", x"84", x"1c", x"12", x"2d", x"3f", x"2c", x"26", x"2a", x"22", x"1b", 
        x"36", x"2b", x"1c", x"80", x"d8", x"cc", x"cb", x"da", x"c9", x"bb", x"c5", x"e0", x"e1", x"df", x"de", 
        x"e0", x"e2", x"e4", x"e6", x"e6", x"e5", x"e5", x"e6", x"e2", x"e4", x"e4", x"e0", x"e1", x"e1", x"de", 
        x"e8", x"e4", x"e8", x"e6", x"e6", x"e4", x"e5", x"e8", x"e7", x"e4", x"e2", x"e3", x"e2", x"e3", x"e4", 
        x"e7", x"e5", x"e5", x"e8", x"e4", x"e5", x"e2", x"e2", x"e6", x"e9", x"e7", x"e6", x"e5", x"e1", x"e7", 
        x"e3", x"e0", x"e4", x"e3", x"e7", x"e6", x"e2", x"e7", x"e2", x"e4", x"e8", x"e8", x"e6", x"e4", x"e3", 
        x"e3", x"e4", x"e7", x"e4", x"e4", x"e3", x"e0", x"e7", x"e6", x"e2", x"e3", x"e5", x"e9", x"e3", x"e4", 
        x"df", x"d6", x"de", x"ea", x"e6", x"e4", x"e8", x"e8", x"e6", x"e5", x"ec", x"eb", x"e6", x"e8", x"ee", 
        x"ed", x"eb", x"e6", x"e7", x"e9", x"e9", x"ed", x"eb", x"e6", x"e7", x"ed", x"ea", x"ea", x"eb", x"e9", 
        x"ee", x"ea", x"e9", x"ea", x"e9", x"ea", x"e9", x"e6", x"e0", x"dc", x"e5", x"eb", x"ec", x"ee", x"e9", 
        x"e8", x"ea", x"e7", x"eb", x"ea", x"e9", x"ea", x"e9", x"e7", x"e7", x"e9", x"e7", x"ec", x"ed", x"e9", 
        x"e8", x"e7", x"ed", x"e9", x"e3", x"e7", x"eb", x"ea", x"e6", x"eb", x"ed", x"e7", x"e6", x"e8", x"eb", 
        x"eb", x"ee", x"eb", x"e8", x"eb", x"ec", x"e8", x"ed", x"ea", x"e8", x"e8", x"e8", x"ed", x"ee", x"ec", 
        x"e8", x"ea", x"eb", x"e8", x"ea", x"ec", x"ed", x"ef", x"ee", x"ea", x"e6", x"e2", x"e6", x"ed", x"ea", 
        x"e8", x"e7", x"e7", x"e8", x"e4", x"ea", x"ed", x"e7", x"e6", x"e6", x"ea", x"e8", x"e6", x"e9", x"e8", 
        x"e8", x"ea", x"e7", x"e8", x"e9", x"e9", x"ec", x"ec", x"eb", x"e9", x"e7", x"ea", x"e8", x"e5", x"e8", 
        x"eb", x"e8", x"e8", x"e9", x"eb", x"ed", x"ed", x"ea", x"e8", x"e8", x"ea", x"ec", x"eb", x"eb", x"eb", 
        x"ec", x"eb", x"ec", x"ea", x"e5", x"e6", x"e9", x"e7", x"ec", x"ef", x"ec", x"ec", x"e9", x"e9", x"ed", 
        x"ef", x"ef", x"ea", x"e6", x"e7", x"ec", x"f0", x"ea", x"e1", x"ee", x"ef", x"eb", x"eb", x"eb", x"ea", 
        x"e8", x"e6", x"ec", x"ed", x"ea", x"ea", x"e8", x"eb", x"ec", x"e8", x"ea", x"ec", x"ec", x"ea", x"e9", 
        x"e9", x"eb", x"e5", x"dc", x"e8", x"ef", x"ee", x"ed", x"ee", x"ee", x"ee", x"ec", x"ec", x"ec", x"ee", 
        x"ed", x"e8", x"e7", x"ea", x"ed", x"ea", x"e4", x"e3", x"e9", x"ec", x"ed", x"ed", x"eb", x"eb", x"ec", 
        x"ec", x"ec", x"ed", x"ea", x"ec", x"eb", x"ec", x"ea", x"ea", x"ea", x"ea", x"eb", x"eb", x"ec", x"eb", 
        x"ea", x"ea", x"eb", x"ec", x"ed", x"ed", x"ec", x"e9", x"ed", x"ed", x"ed", x"eb", x"ed", x"f1", x"ef", 
        x"ed", x"ec", x"eb", x"ec", x"ec", x"ee", x"ec", x"ed", x"ef", x"ee", x"ed", x"ea", x"e8", x"eb", x"ed", 
        x"ef", x"e2", x"dc", x"ea", x"ef", x"f1", x"ec", x"ee", x"ee", x"f0", x"f2", x"ef", x"ea", x"ef", x"ef", 
        x"ee", x"ef", x"ef", x"ed", x"f0", x"f2", x"f1", x"ef", x"ed", x"ee", x"ee", x"ef", x"f1", x"f0", x"f0", 
        x"ee", x"ec", x"ef", x"f1", x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f5", x"f8", x"f6", x"f6", x"f4", 
        x"ef", x"ef", x"ee", x"f0", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"f2", x"f1", x"f1", x"ef", x"ed", 
        x"ee", x"ee", x"eb", x"ee", x"e8", x"e8", x"ef", x"f0", x"f0", x"ef", x"ef", x"ee", x"ed", x"ed", x"ef", 
        x"ef", x"f0", x"ef", x"f0", x"ef", x"ef", x"ef", x"ee", x"f0", x"ef", x"f0", x"f0", x"ef", x"ef", x"ef", 
        x"f2", x"f6", x"f7", x"f4", x"f1", x"f2", x"f4", x"f4", x"f3", x"f0", x"f0", x"f0", x"f0", x"ee", x"ef", 
        x"f0", x"f0", x"ee", x"ee", x"ef", x"f0", x"f1", x"f2", x"ef", x"ef", x"ee", x"ee", x"ef", x"e9", x"e7", 
        x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"f0", x"f1", x"ef", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"f2", x"f0", x"f0", x"f1", x"f4", x"f6", x"f1", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"f0", 
        x"f0", x"ef", x"ed", x"ed", x"ee", x"ee", x"f1", x"ee", x"f0", x"e2", x"a9", x"a8", x"c0", x"ab", x"90", 
        x"a3", x"98", x"79", x"6a", x"75", x"a3", x"b5", x"b8", x"c0", x"e6", x"ef", x"e2", x"5c", x"1f", x"1f", 
        x"1e", x"2c", x"54", x"78", x"a5", x"c5", x"d7", x"cc", x"d1", x"d9", x"d9", x"9a", x"3e", x"3f", x"45", 
        x"4a", x"50", x"51", x"52", x"53", x"4f", x"57", x"5d", x"40", x"20", x"40", x"7d", x"ab", x"a1", x"52", 
        x"1d", x"11", x"08", x"03", x"06", x"14", x"16", x"17", x"10", x"1d", x"65", x"b8", x"c3", x"66", x"10", 
        x"0c", x"09", x"0f", x"2a", x"34", x"2b", x"2c", x"26", x"24", x"22", x"20", x"20", x"24", x"0f", x"04", 
        x"04", x"06", x"03", x"03", x"07", x"06", x"03", x"05", x"08", x"05", x"02", x"02", x"05", x"07", x"05", 
        x"11", x"27", x"71", x"94", x"9b", x"92", x"9b", x"ba", x"c4", x"c9", x"c9", x"ba", x"90", x"8e", x"c3", 
        x"d9", x"7a", x"25", x"2c", x"32", x"38", x"40", x"4f", x"53", x"4f", x"4b", x"51", x"65", x"5d", x"3c", 
        x"34", x"3c", x"5a", x"5e", x"5f", x"58", x"3c", x"30", x"57", x"55", x"11", x"49", x"83", x"9a", x"b8", 
        x"a7", x"3c", x"30", x"36", x"43", x"57", x"4f", x"3e", x"3b", x"3c", x"46", x"46", x"40", x"3d", x"41", 
        x"3c", x"31", x"5b", x"9e", x"aa", x"b4", x"98", x"8d", x"ab", x"b4", x"45", x"13", x"16", x"1a", x"16", 
        x"13", x"12", x"13", x"14", x"10", x"0d", x"0f", x"15", x"16", x"1c", x"06", x"05", x"07", x"0a", x"08", 
        x"3a", x"36", x"17", x"53", x"c1", x"88", x"1f", x"20", x"2e", x"38", x"2c", x"29", x"2b", x"25", x"20", 
        x"32", x"35", x"21", x"8f", x"d6", x"c4", x"c6", x"d7", x"c3", x"c2", x"d2", x"dc", x"dd", x"e1", x"e1", 
        x"e3", x"e2", x"e2", x"e6", x"e9", x"e7", x"e1", x"e0", x"db", x"de", x"de", x"de", x"e3", x"e0", x"e0", 
        x"e9", x"e5", x"e7", x"e5", x"e3", x"e3", x"e6", x"e2", x"df", x"e1", x"df", x"df", x"e2", x"e3", x"e7", 
        x"e7", x"e4", x"e6", x"e8", x"e1", x"e4", x"e9", x"e4", x"e7", x"ea", x"e7", x"e8", x"e1", x"de", x"e5", 
        x"e4", x"e3", x"e5", x"e8", x"e5", x"e6", x"e7", x"e5", x"e5", x"e9", x"ed", x"e8", x"e4", x"e5", x"e5", 
        x"e5", x"e4", x"e3", x"e7", x"e9", x"e8", x"e6", x"eb", x"e9", x"e6", x"e9", x"e7", x"e7", x"e2", x"e3", 
        x"e3", x"e1", x"e6", x"eb", x"ec", x"ec", x"f1", x"ec", x"e8", x"ea", x"e7", x"e7", x"e8", x"e8", x"e9", 
        x"eb", x"e8", x"e9", x"ec", x"eb", x"e7", x"eb", x"ed", x"ed", x"e9", x"ea", x"e7", x"e8", x"e3", x"da", 
        x"e4", x"e8", x"eb", x"e9", x"e8", x"ed", x"ed", x"ec", x"e7", x"e1", x"e8", x"ea", x"e6", x"e8", x"e8", 
        x"e9", x"ea", x"e6", x"e8", x"e8", x"ea", x"ea", x"ea", x"e7", x"e5", x"e9", x"e7", x"ec", x"ec", x"ea", 
        x"e9", x"ea", x"ea", x"e3", x"e1", x"ea", x"eb", x"e9", x"e5", x"eb", x"ed", x"e8", x"e7", x"e8", x"e9", 
        x"e8", x"e9", x"eb", x"ea", x"ef", x"ef", x"e8", x"e9", x"ea", x"ea", x"e8", x"e9", x"eb", x"e9", x"eb", 
        x"ea", x"ea", x"e9", x"e7", x"e9", x"e7", x"e8", x"ee", x"ec", x"e9", x"e9", x"e7", x"e9", x"ee", x"ec", 
        x"eb", x"ec", x"ec", x"eb", x"e3", x"e8", x"ec", x"e8", x"e7", x"e7", x"e8", x"e5", x"e6", x"e8", x"e9", 
        x"e8", x"eb", x"e7", x"ea", x"ed", x"eb", x"ec", x"e7", x"e5", x"e7", x"e9", x"ec", x"ea", x"e8", x"ee", 
        x"f0", x"ea", x"e9", x"ea", x"ec", x"ed", x"ef", x"ec", x"ea", x"eb", x"ed", x"ee", x"ed", x"ec", x"ee", 
        x"ed", x"eb", x"ee", x"ef", x"ed", x"ec", x"eb", x"eb", x"ee", x"ee", x"eb", x"ed", x"ed", x"ed", x"ee", 
        x"ed", x"ee", x"ec", x"e9", x"ec", x"ec", x"e9", x"e4", x"db", x"e5", x"ea", x"ea", x"e8", x"ea", x"ec", 
        x"eb", x"ea", x"e9", x"e6", x"e8", x"e9", x"e3", x"e5", x"e1", x"df", x"ea", x"eb", x"ec", x"ec", x"eb", 
        x"eb", x"ee", x"e9", x"e0", x"e9", x"ed", x"ea", x"ea", x"ee", x"ec", x"eb", x"e9", x"e9", x"e9", x"eb", 
        x"e9", x"e3", x"e4", x"e8", x"e9", x"e7", x"e5", x"e6", x"ea", x"ec", x"ed", x"ec", x"ea", x"e9", x"e9", 
        x"e9", x"eb", x"ee", x"eb", x"ec", x"ec", x"ed", x"eb", x"eb", x"eb", x"eb", x"eb", x"ea", x"eb", x"ea", 
        x"e9", x"e9", x"eb", x"ed", x"ed", x"ed", x"ed", x"eb", x"eb", x"ee", x"ee", x"ed", x"ed", x"ed", x"ed", 
        x"ed", x"ef", x"ef", x"ef", x"ee", x"ec", x"eb", x"ef", x"ef", x"ec", x"eb", x"e7", x"e7", x"e9", x"eb", 
        x"f0", x"e0", x"d9", x"e9", x"ef", x"ee", x"ec", x"ef", x"f0", x"f1", x"f2", x"ef", x"eb", x"ef", x"ef", 
        x"ef", x"f1", x"f0", x"ed", x"f0", x"ee", x"f0", x"ef", x"ed", x"ef", x"f2", x"f1", x"f1", x"ef", x"ef", 
        x"ef", x"ed", x"f0", x"f2", x"f0", x"ee", x"ee", x"f0", x"ef", x"ef", x"f4", x"f9", x"f5", x"f6", x"f3", 
        x"ef", x"ef", x"ee", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"f1", x"f0", x"ed", x"ee", x"ed", x"ee", 
        x"f0", x"f0", x"ed", x"ed", x"e9", x"e8", x"ef", x"ee", x"f0", x"f0", x"ee", x"ee", x"ef", x"ef", x"ee", 
        x"ee", x"ee", x"ee", x"ef", x"ee", x"ef", x"f0", x"ee", x"f1", x"ef", x"ef", x"f0", x"ef", x"ef", x"f1", 
        x"f5", x"f8", x"f7", x"f4", x"f2", x"f4", x"f5", x"f3", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", 
        x"f0", x"f1", x"f1", x"ef", x"ef", x"f1", x"f1", x"f0", x"ee", x"ef", x"ed", x"ee", x"f1", x"ea", x"e7", 
        x"ef", x"f0", x"f0", x"f0", x"ef", x"ef", x"ef", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ee", x"ed", 
        x"f0", x"ee", x"ee", x"f0", x"f3", x"f5", x"f0", x"ef", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", 
        x"ef", x"ef", x"ee", x"ef", x"ee", x"ed", x"ee", x"eb", x"ef", x"ef", x"a5", x"a1", x"b4", x"b0", x"9b", 
        x"a7", x"ad", x"88", x"7a", x"74", x"97", x"ad", x"ac", x"ab", x"d3", x"dd", x"cf", x"73", x"59", x"61", 
        x"64", x"66", x"6f", x"74", x"a8", x"c5", x"d8", x"d0", x"d3", x"d5", x"dd", x"ba", x"6c", x"61", x"62", 
        x"63", x"64", x"5e", x"57", x"55", x"4e", x"53", x"61", x"60", x"73", x"93", x"82", x"93", x"66", x"31", 
        x"29", x"0f", x"07", x"03", x"08", x"0f", x"15", x"20", x"11", x"3b", x"8c", x"c9", x"d8", x"7c", x"13", 
        x"0d", x"0e", x"0c", x"0e", x"1c", x"1b", x"1d", x"1b", x"21", x"24", x"1f", x"29", x"28", x"0c", x"05", 
        x"03", x"05", x"03", x"02", x"04", x"03", x"05", x"08", x"05", x"05", x"04", x"01", x"03", x"03", x"11", 
        x"52", x"81", x"87", x"97", x"8a", x"78", x"95", x"b4", x"ba", x"c2", x"c7", x"ba", x"9b", x"90", x"aa", 
        x"d1", x"aa", x"58", x"60", x"67", x"64", x"62", x"5c", x"52", x"52", x"56", x"53", x"57", x"4c", x"3c", 
        x"3a", x"40", x"3e", x"3e", x"3d", x"2a", x"19", x"2d", x"41", x"5c", x"17", x"51", x"8e", x"97", x"b9", 
        x"84", x"26", x"32", x"33", x"25", x"15", x"10", x"11", x"10", x"0e", x"21", x"15", x"0f", x"0d", x"0e", 
        x"0e", x"16", x"42", x"6b", x"7d", x"b4", x"b5", x"8a", x"aa", x"bf", x"45", x"0d", x"0e", x"15", x"0d", 
        x"0d", x"15", x"14", x"0c", x"0e", x"0e", x"14", x"13", x"1e", x"27", x"0f", x"0f", x"10", x"0c", x"0e", 
        x"7c", x"49", x"27", x"40", x"83", x"63", x"2b", x"30", x"2f", x"32", x"32", x"32", x"32", x"2c", x"2a", 
        x"2a", x"27", x"24", x"8e", x"e0", x"d0", x"ce", x"dd", x"d1", x"cf", x"d4", x"d7", x"dc", x"e4", x"e1", 
        x"e3", x"e2", x"e4", x"e5", x"e5", x"e6", x"e9", x"e6", x"e6", x"e3", x"e0", x"e4", x"e4", x"e2", x"e3", 
        x"e8", x"e5", x"e6", x"e7", x"e9", x"e6", x"e5", x"df", x"df", x"eb", x"eb", x"e6", x"e6", x"e6", x"e9", 
        x"e7", x"e4", x"e7", x"e5", x"e1", x"e4", x"e6", x"df", x"e5", x"ea", x"e4", x"e3", x"dc", x"d9", x"e0", 
        x"e6", x"e8", x"e5", x"e6", x"df", x"e7", x"e9", x"e4", x"e8", x"e7", x"e6", x"e2", x"e3", x"e7", x"e9", 
        x"ea", x"e9", x"e4", x"e6", x"e4", x"e4", x"e8", x"e9", x"e8", x"e7", x"e9", x"e6", x"e6", x"e5", x"e3", 
        x"e1", x"e5", x"e8", x"e5", x"e2", x"e6", x"e6", x"e3", x"e8", x"ea", x"e2", x"e3", x"e9", x"e5", x"de", 
        x"e6", x"e9", x"e6", x"ed", x"ef", x"e7", x"e9", x"ea", x"eb", x"e6", x"ea", x"e5", x"e8", x"ea", x"e7", 
        x"e7", x"e6", x"e9", x"e8", x"ea", x"ef", x"eb", x"e8", x"e8", x"e9", x"eb", x"ea", x"e9", x"ee", x"eb", 
        x"e8", x"ea", x"eb", x"e8", x"e7", x"ea", x"e6", x"ea", x"e7", x"e9", x"ed", x"e8", x"e7", x"e5", x"e5", 
        x"eb", x"e9", x"ea", x"eb", x"ec", x"e7", x"e7", x"ea", x"e4", x"e9", x"ec", x"e9", x"ea", x"ea", x"eb", 
        x"eb", x"ea", x"ee", x"ea", x"ec", x"e9", x"e4", x"eb", x"ef", x"e9", x"e7", x"ec", x"e7", x"ea", x"ec", 
        x"e8", x"ec", x"ef", x"eb", x"e7", x"e5", x"ed", x"ee", x"e7", x"e4", x"ec", x"ee", x"ec", x"ec", x"eb", 
        x"e9", x"e8", x"eb", x"ec", x"e5", x"e6", x"e8", x"e8", x"e8", x"e7", x"e7", x"e5", x"e8", x"eb", x"eb", 
        x"e9", x"ea", x"e6", x"e8", x"ed", x"e7", x"ed", x"e7", x"e1", x"e4", x"e7", x"eb", x"e9", x"e9", x"ed", 
        x"ee", x"e9", x"e7", x"e8", x"e9", x"ea", x"eb", x"ea", x"e9", x"ea", x"eb", x"eb", x"e9", x"e7", x"ea", 
        x"ec", x"ea", x"ea", x"eb", x"ee", x"ec", x"ea", x"ed", x"ee", x"ec", x"eb", x"ea", x"ee", x"ef", x"ee", 
        x"e9", x"eb", x"ec", x"eb", x"f1", x"ed", x"e7", x"ef", x"ed", x"ea", x"eb", x"eb", x"e9", x"ea", x"ee", 
        x"ed", x"ef", x"ec", x"e9", x"eb", x"ec", x"e7", x"eb", x"e9", x"e5", x"ec", x"ea", x"ec", x"ec", x"ea", 
        x"ea", x"eb", x"e4", x"dc", x"e8", x"ef", x"ee", x"ed", x"ef", x"ed", x"ec", x"eb", x"eb", x"e9", x"ec", 
        x"ec", x"eb", x"ed", x"ec", x"e9", x"ea", x"ed", x"ee", x"ef", x"ef", x"ed", x"ed", x"eb", x"eb", x"ec", 
        x"ea", x"ea", x"ec", x"e9", x"ea", x"eb", x"ec", x"ea", x"e9", x"ea", x"eb", x"eb", x"ec", x"ec", x"ea", 
        x"ea", x"eb", x"ec", x"ed", x"ec", x"ee", x"f0", x"f0", x"ec", x"ed", x"ee", x"f0", x"ee", x"e7", x"eb", 
        x"ee", x"ee", x"ee", x"ed", x"ec", x"ec", x"ed", x"ed", x"e8", x"e7", x"eb", x"ec", x"ed", x"eb", x"ea", 
        x"f1", x"e5", x"dd", x"ee", x"ee", x"ec", x"eb", x"ed", x"ee", x"ed", x"ee", x"ec", x"ea", x"ef", x"ee", 
        x"ed", x"f0", x"f0", x"ec", x"ee", x"ef", x"f2", x"ef", x"eb", x"ed", x"f2", x"f2", x"f1", x"ef", x"ef", 
        x"f0", x"ef", x"f2", x"f2", x"f1", x"ef", x"ef", x"f2", x"ef", x"eb", x"f1", x"f6", x"f5", x"f5", x"f2", 
        x"ee", x"ee", x"ed", x"f0", x"f0", x"f0", x"f0", x"f1", x"f2", x"f2", x"ef", x"ec", x"ee", x"ef", x"ef", 
        x"ee", x"ed", x"ee", x"ed", x"ea", x"e9", x"f1", x"ee", x"ef", x"f0", x"ef", x"ef", x"f0", x"f0", x"ef", 
        x"ed", x"ec", x"ed", x"f0", x"ee", x"ef", x"f0", x"ed", x"f0", x"f0", x"f2", x"f2", x"f1", x"f0", x"f1", 
        x"f4", x"f6", x"f7", x"f4", x"f2", x"f2", x"f3", x"f2", x"ef", x"ef", x"f1", x"f1", x"f0", x"f0", x"f0", 
        x"f0", x"f2", x"f2", x"f0", x"ef", x"f0", x"f0", x"ef", x"ed", x"ed", x"ed", x"ef", x"f1", x"eb", x"e8", 
        x"f0", x"f0", x"f0", x"ef", x"f0", x"ef", x"ef", x"ee", x"ec", x"eb", x"ed", x"f0", x"ee", x"ed", x"ed", 
        x"ef", x"ee", x"ef", x"f0", x"f3", x"f6", x"f1", x"ef", x"ef", x"ee", x"ee", x"ee", x"ef", x"f0", x"ef", 
        x"ed", x"f0", x"f0", x"f0", x"ee", x"ee", x"ed", x"f0", x"f0", x"ee", x"b4", x"aa", x"bc", x"ae", x"9b", 
        x"a5", x"a8", x"81", x"89", x"6c", x"94", x"aa", x"bc", x"a4", x"6f", x"56", x"54", x"5c", x"5d", x"54", 
        x"4b", x"5b", x"6c", x"5b", x"95", x"b5", x"d2", x"d0", x"d4", x"d6", x"df", x"bb", x"49", x"1b", x"22", 
        x"24", x"26", x"1f", x"20", x"25", x"24", x"51", x"77", x"69", x"77", x"98", x"7b", x"3a", x"2e", x"38", 
        x"3f", x"21", x"19", x"0d", x"06", x"11", x"1e", x"1d", x"08", x"27", x"a0", x"ed", x"ea", x"8c", x"13", 
        x"1b", x"43", x"35", x"1e", x"49", x"59", x"5c", x"5e", x"61", x"59", x"57", x"69", x"49", x"17", x"08", 
        x"06", x"1d", x"1d", x"13", x"22", x"13", x"08", x"08", x"05", x"04", x"02", x"02", x"03", x"02", x"17", 
        x"65", x"80", x"7e", x"78", x"73", x"75", x"9d", x"b1", x"b4", x"c2", x"c6", x"b9", x"9c", x"8c", x"af", 
        x"cb", x"9d", x"32", x"1d", x"1f", x"16", x"17", x"16", x"0f", x"10", x"13", x"11", x"1f", x"44", x"41", 
        x"3d", x"32", x"17", x"09", x"09", x"06", x"0a", x"2c", x"37", x"53", x"33", x"62", x"9e", x"9d", x"9c", 
        x"56", x"27", x"3f", x"25", x"0f", x"0b", x"10", x"12", x"10", x"16", x"30", x"1d", x"16", x"19", x"1d", 
        x"17", x"1d", x"45", x"87", x"81", x"92", x"c1", x"9f", x"a4", x"b8", x"4f", x"25", x"2b", x"3b", x"3f", 
        x"43", x"53", x"55", x"46", x"46", x"44", x"42", x"45", x"63", x"6a", x"5a", x"5c", x"5a", x"4d", x"4f", 
        x"8d", x"52", x"39", x"65", x"ae", x"71", x"27", x"32", x"33", x"3e", x"45", x"36", x"38", x"31", x"36", 
        x"32", x"2b", x"22", x"79", x"dd", x"ca", x"c9", x"dc", x"ca", x"c8", x"d4", x"d5", x"d9", x"e4", x"da", 
        x"dc", x"e2", x"e5", x"e5", x"e2", x"e1", x"e5", x"e3", x"e1", x"e7", x"e5", x"e6", x"e6", x"de", x"dd", 
        x"e3", x"e8", x"e1", x"e1", x"e3", x"e6", x"e1", x"de", x"e0", x"ea", x"ea", x"e5", x"e4", x"e4", x"e7", 
        x"e2", x"e7", x"eb", x"e1", x"e0", x"e4", x"e5", x"e5", x"e5", x"e6", x"e5", x"e6", x"e1", x"e5", x"e6", 
        x"e6", x"e5", x"e9", x"ea", x"e3", x"e8", x"e6", x"e5", x"e4", x"e5", x"e3", x"df", x"e2", x"e3", x"e5", 
        x"e6", x"e9", x"e9", x"e7", x"e5", x"e6", x"e7", x"ea", x"e6", x"e4", x"e5", x"e6", x"e7", x"e3", x"e5", 
        x"e4", x"e6", x"e6", x"e5", x"dc", x"d8", x"db", x"e5", x"e9", x"e8", x"ea", x"ec", x"ec", x"e1", x"db", 
        x"e3", x"e5", x"e4", x"e7", x"e8", x"e4", x"e8", x"ee", x"e8", x"e1", x"eb", x"e9", x"e5", x"e6", x"e5", 
        x"e1", x"e7", x"e6", x"e6", x"e9", x"ec", x"e8", x"e7", x"e8", x"e7", x"ea", x"e9", x"e7", x"ec", x"ef", 
        x"ea", x"e8", x"ea", x"eb", x"e8", x"eb", x"e8", x"e9", x"e9", x"ed", x"ef", x"eb", x"e9", x"e6", x"e4", 
        x"ea", x"e8", x"ee", x"eb", x"ec", x"e5", x"e4", x"eb", x"e8", x"e9", x"eb", x"e8", x"eb", x"e9", x"e4", 
        x"e8", x"ea", x"ea", x"e8", x"e8", x"eb", x"eb", x"e5", x"e6", x"eb", x"e7", x"e9", x"ea", x"ec", x"e8", 
        x"e7", x"e7", x"ea", x"ec", x"e9", x"e5", x"eb", x"e8", x"e5", x"e7", x"eb", x"ea", x"e6", x"e9", x"ed", 
        x"ec", x"e8", x"e9", x"e9", x"e3", x"e7", x"e9", x"e8", x"e8", x"e9", x"e8", x"e3", x"e7", x"ec", x"eb", 
        x"e9", x"e9", x"e8", x"e5", x"ec", x"e8", x"ea", x"eb", x"e9", x"ec", x"e9", x"e5", x"e7", x"ea", x"e7", 
        x"e7", x"e9", x"e8", x"ea", x"e9", x"e9", x"ea", x"ea", x"ed", x"ee", x"e9", x"e8", x"e9", x"ec", x"ea", 
        x"eb", x"ec", x"ea", x"ed", x"ee", x"ec", x"ee", x"ec", x"eb", x"ee", x"ec", x"e8", x"e8", x"eb", x"ec", 
        x"ea", x"ea", x"eb", x"eb", x"ee", x"ee", x"ec", x"ee", x"ed", x"eb", x"ed", x"e9", x"ea", x"eb", x"ea", 
        x"e9", x"e9", x"e9", x"ea", x"eb", x"eb", x"e9", x"e9", x"e9", x"ec", x"ed", x"e8", x"e8", x"ec", x"ec", 
        x"ea", x"e8", x"e5", x"df", x"e9", x"ed", x"eb", x"ea", x"ee", x"f0", x"eb", x"ed", x"e9", x"e5", x"ea", 
        x"ea", x"eb", x"eb", x"e9", x"ea", x"ee", x"ec", x"eb", x"ec", x"ec", x"e7", x"ed", x"eb", x"ed", x"ee", 
        x"ee", x"ec", x"ea", x"e9", x"ea", x"ea", x"e9", x"e6", x"e7", x"ec", x"ec", x"ec", x"ee", x"ec", x"e8", 
        x"ec", x"ed", x"ec", x"ef", x"eb", x"eb", x"ee", x"ec", x"ef", x"ee", x"eb", x"ef", x"ed", x"ed", x"ea", 
        x"eb", x"ed", x"ef", x"ee", x"eb", x"e8", x"ed", x"ee", x"ea", x"ea", x"ea", x"e9", x"ea", x"ea", x"e9", 
        x"eb", x"e7", x"dd", x"ee", x"ed", x"ec", x"e9", x"ed", x"ef", x"ed", x"ec", x"ec", x"ee", x"f2", x"ef", 
        x"ee", x"f0", x"f0", x"ee", x"ed", x"ef", x"ef", x"ef", x"ee", x"ef", x"ef", x"ef", x"ee", x"f1", x"f1", 
        x"f1", x"ef", x"ef", x"ef", x"f1", x"f1", x"f0", x"f3", x"f0", x"f2", x"f5", x"f6", x"f5", x"f3", x"f0", 
        x"ed", x"ec", x"ed", x"ee", x"f1", x"ef", x"ed", x"ec", x"ee", x"f1", x"f1", x"ef", x"ed", x"ec", x"f1", 
        x"ed", x"eb", x"ed", x"ef", x"eb", x"e7", x"f1", x"f0", x"ef", x"ef", x"f0", x"ef", x"ee", x"ef", x"ef", 
        x"ee", x"ef", x"f0", x"f0", x"ee", x"ee", x"f0", x"ed", x"ed", x"f1", x"f0", x"f1", x"f1", x"f1", x"f1", 
        x"f4", x"f7", x"f7", x"f5", x"ef", x"ed", x"ef", x"f1", x"ef", x"ef", x"f1", x"f1", x"ef", x"f0", x"ef", 
        x"ee", x"ee", x"ee", x"ed", x"ee", x"ef", x"f0", x"f0", x"ee", x"eb", x"eb", x"ee", x"ec", x"ec", x"ea", 
        x"ee", x"ee", x"f0", x"ed", x"f1", x"ee", x"ee", x"f1", x"ed", x"ed", x"f0", x"f1", x"ee", x"ed", x"f0", 
        x"ed", x"ef", x"ef", x"ed", x"ee", x"f1", x"f1", x"f0", x"f1", x"f1", x"ef", x"ef", x"f0", x"f0", x"f0", 
        x"ec", x"ee", x"ec", x"ef", x"ec", x"ee", x"ef", x"f3", x"ef", x"ed", x"aa", x"9d", x"bf", x"a6", x"ab", 
        x"b4", x"b1", x"73", x"7d", x"62", x"99", x"a4", x"bb", x"88", x"2d", x"34", x"26", x"21", x"25", x"24", 
        x"1f", x"3b", x"67", x"4f", x"86", x"c0", x"c6", x"d1", x"d8", x"da", x"e2", x"ce", x"64", x"2f", x"34", 
        x"36", x"3a", x"33", x"31", x"33", x"41", x"63", x"6d", x"67", x"68", x"68", x"63", x"44", x"41", x"56", 
        x"55", x"4a", x"52", x"47", x"16", x"10", x"16", x"11", x"07", x"32", x"a4", x"db", x"d8", x"93", x"17", 
        x"1a", x"25", x"19", x"15", x"33", x"39", x"35", x"30", x"2d", x"26", x"23", x"22", x"15", x"0e", x"05", 
        x"13", x"69", x"67", x"32", x"46", x"22", x"07", x"05", x"01", x"03", x"03", x"03", x"03", x"04", x"1b", 
        x"67", x"85", x"77", x"64", x"5c", x"87", x"ac", x"b7", x"bf", x"c5", x"c8", x"bb", x"96", x"7d", x"ac", 
        x"d8", x"8f", x"1d", x"0a", x"0e", x"0d", x"16", x"1c", x"10", x"11", x"10", x"0d", x"24", x"4a", x"46", 
        x"4a", x"34", x"1e", x"14", x"13", x"15", x"13", x"2f", x"38", x"5e", x"7c", x"6a", x"a3", x"bb", x"8e", 
        x"48", x"4c", x"77", x"57", x"35", x"43", x"48", x"4a", x"4a", x"4c", x"59", x"54", x"4f", x"5c", x"60", 
        x"5a", x"61", x"5d", x"70", x"81", x"9a", x"bb", x"ac", x"9f", x"bd", x"73", x"5c", x"63", x"6d", x"71", 
        x"5f", x"56", x"52", x"4d", x"4c", x"4d", x"51", x"46", x"46", x"43", x"41", x"3b", x"3b", x"47", x"3f", 
        x"5d", x"49", x"55", x"9a", x"cd", x"69", x"27", x"32", x"2f", x"47", x"4f", x"2f", x"33", x"36", x"3b", 
        x"31", x"23", x"19", x"6f", x"d8", x"c9", x"c9", x"de", x"c6", x"bc", x"c9", x"d4", x"dc", x"e4", x"dd", 
        x"e0", x"e2", x"e6", x"e0", x"dc", x"e9", x"e4", x"e3", x"e3", x"e8", x"e5", x"e4", x"e4", x"de", x"dc", 
        x"e5", x"e7", x"df", x"e4", x"e1", x"e2", x"e6", x"e7", x"e3", x"e1", x"e0", x"e4", x"e7", x"e5", x"e8", 
        x"e3", x"e6", x"e8", x"e3", x"e4", x"e4", x"e5", x"e4", x"e2", x"e2", x"e1", x"e3", x"e6", x"ea", x"e4", 
        x"e1", x"e3", x"e8", x"e7", x"e1", x"e4", x"e5", x"e5", x"e3", x"e4", x"e1", x"e3", x"e6", x"e7", x"e8", 
        x"e7", x"ea", x"eb", x"e6", x"e7", x"e6", x"e7", x"e9", x"e6", x"e4", x"e3", x"e6", x"ea", x"e7", x"e4", 
        x"e3", x"e8", x"e8", x"e7", x"e4", x"e3", x"e5", x"ea", x"ea", x"e9", x"ea", x"ea", x"e8", x"df", x"d8", 
        x"e1", x"e8", x"e8", x"e4", x"e7", x"e9", x"ea", x"ee", x"e8", x"e3", x"ea", x"ed", x"e5", x"e2", x"e3", 
        x"e0", x"e9", x"e8", x"e7", x"e9", x"e9", x"e7", x"e5", x"e8", x"e5", x"e6", x"e7", x"e6", x"e8", x"ea", 
        x"e9", x"e8", x"e6", x"e8", x"e8", x"e9", x"e9", x"eb", x"e5", x"e9", x"e8", x"e7", x"e6", x"e6", x"ea", 
        x"e7", x"d9", x"e5", x"e9", x"e7", x"e5", x"e7", x"e9", x"e9", x"e9", x"ea", x"e8", x"eb", x"ea", x"e3", 
        x"e5", x"e8", x"ea", x"e7", x"e7", x"eb", x"ed", x"ea", x"e7", x"e8", x"e6", x"e9", x"ea", x"ea", x"e8", 
        x"e9", x"eb", x"ee", x"ef", x"ea", x"e5", x"e9", x"e9", x"e8", x"e9", x"ec", x"eb", x"e4", x"e8", x"eb", 
        x"eb", x"eb", x"e9", x"e7", x"e3", x"e9", x"eb", x"e8", x"e8", x"ea", x"e9", x"e5", x"e7", x"eb", x"eb", 
        x"e8", x"e8", x"e8", x"e6", x"e9", x"e7", x"e9", x"e9", x"e7", x"eb", x"eb", x"eb", x"e8", x"e8", x"e6", 
        x"e7", x"ea", x"e9", x"ea", x"e9", x"ea", x"eb", x"ec", x"ee", x"ed", x"e9", x"e9", x"eb", x"ec", x"e8", 
        x"e9", x"ef", x"eb", x"eb", x"ed", x"ed", x"ee", x"eb", x"ea", x"eb", x"ea", x"e9", x"e8", x"eb", x"ed", 
        x"e9", x"e7", x"e8", x"ee", x"ee", x"ed", x"ec", x"ee", x"ee", x"e9", x"ec", x"e9", x"ec", x"ed", x"eb", 
        x"ea", x"e8", x"e9", x"eb", x"eb", x"ec", x"ec", x"eb", x"e8", x"ea", x"ed", x"eb", x"e9", x"eb", x"eb", 
        x"e7", x"e6", x"e9", x"e1", x"ea", x"ed", x"e9", x"e8", x"ed", x"ed", x"eb", x"eb", x"e8", x"e7", x"ed", 
        x"eb", x"ea", x"e9", x"e9", x"ea", x"ec", x"ea", x"e7", x"ec", x"ec", x"e7", x"ec", x"eb", x"ed", x"ee", 
        x"eb", x"ea", x"ea", x"ea", x"e9", x"e9", x"ea", x"e9", x"e9", x"ed", x"eb", x"ea", x"ed", x"ea", x"e7", 
        x"ec", x"ee", x"ec", x"ee", x"ea", x"e9", x"ec", x"ec", x"ee", x"ec", x"eb", x"f0", x"ed", x"ec", x"ec", 
        x"ec", x"ee", x"ef", x"ef", x"ed", x"ec", x"ec", x"ea", x"e8", x"ea", x"eb", x"ea", x"eb", x"ec", x"ea", 
        x"eb", x"e7", x"dc", x"ee", x"ee", x"ef", x"ed", x"ef", x"ef", x"ee", x"ed", x"ee", x"ef", x"ee", x"ed", 
        x"ee", x"ef", x"ed", x"ec", x"ef", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ef", x"ee", x"f0", x"ee", 
        x"ef", x"ef", x"ef", x"f0", x"f1", x"f1", x"ef", x"f0", x"f2", x"f3", x"f6", x"f7", x"f4", x"ee", x"ec", 
        x"ef", x"f0", x"ef", x"ef", x"f1", x"ee", x"ed", x"ee", x"ed", x"ed", x"f0", x"ef", x"ee", x"ed", x"f1", 
        x"ee", x"ed", x"ee", x"f0", x"ed", x"e8", x"f1", x"f1", x"f0", x"f0", x"f0", x"ee", x"ee", x"f0", x"ef", 
        x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"f1", x"ef", x"ed", x"f0", x"f0", x"f1", x"f0", x"f0", x"f1", 
        x"f6", x"f7", x"f4", x"f2", x"ef", x"ee", x"f0", x"f1", x"ee", x"ed", x"ee", x"ef", x"f0", x"f0", x"ef", 
        x"ed", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ed", x"ee", x"ee", x"ec", x"ee", x"ec", x"ec", x"e7", 
        x"ec", x"ec", x"ee", x"ee", x"f3", x"ec", x"ed", x"ee", x"ef", x"f3", x"f1", x"f0", x"f1", x"f2", x"ef", 
        x"ea", x"ed", x"ef", x"ef", x"f2", x"f3", x"f1", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"f0", x"f1", 
        x"eb", x"ef", x"ea", x"ee", x"ef", x"eb", x"ef", x"f3", x"f0", x"ef", x"ba", x"9d", x"b1", x"8f", x"95", 
        x"ac", x"b3", x"7b", x"78", x"68", x"9b", x"ad", x"b4", x"7d", x"37", x"52", x"45", x"38", x"40", x"3f", 
        x"3f", x"45", x"63", x"64", x"90", x"c3", x"ca", x"d7", x"db", x"d5", x"cd", x"c6", x"8e", x"6a", x"6a", 
        x"70", x"6d", x"70", x"69", x"66", x"61", x"5e", x"5d", x"65", x"6e", x"68", x"75", x"78", x"72", x"77", 
        x"6a", x"63", x"67", x"61", x"22", x"05", x"0a", x"08", x"0b", x"3f", x"99", x"af", x"b1", x"86", x"15", 
        x"17", x"15", x"0a", x"05", x"0d", x"0e", x"0e", x"0a", x"0c", x"0c", x"08", x"08", x"04", x"03", x"09", 
        x"1c", x"51", x"3e", x"13", x"12", x"09", x"04", x"02", x"01", x"02", x"04", x"06", x"02", x"02", x"1a", 
        x"5b", x"77", x"5a", x"45", x"62", x"9a", x"b4", x"b6", x"bf", x"c7", x"c9", x"c1", x"a3", x"6f", x"95", 
        x"ce", x"89", x"2e", x"2e", x"31", x"2f", x"40", x"45", x"2e", x"2f", x"2d", x"31", x"43", x"51", x"4f", 
        x"54", x"4d", x"50", x"4b", x"47", x"4d", x"45", x"48", x"3e", x"79", x"b1", x"65", x"8c", x"c2", x"99", 
        x"3d", x"6e", x"a3", x"84", x"69", x"71", x"6d", x"68", x"66", x"5a", x"54", x"4e", x"4b", x"49", x"4b", 
        x"4d", x"52", x"54", x"4e", x"5f", x"8f", x"b9", x"b8", x"a9", x"bc", x"65", x"36", x"3f", x"34", x"28", 
        x"1d", x"1b", x"19", x"14", x"1a", x"19", x"11", x"0e", x"11", x"0d", x"0b", x"09", x"19", x"28", x"10", 
        x"52", x"54", x"4c", x"8e", x"c8", x"64", x"2a", x"2c", x"28", x"46", x"54", x"3e", x"3e", x"3a", x"36", 
        x"2b", x"2d", x"2b", x"78", x"cf", x"c6", x"cd", x"e0", x"ca", x"c1", x"d1", x"e2", x"e0", x"e1", x"e0", 
        x"df", x"de", x"e3", x"d1", x"c6", x"e1", x"e0", x"e3", x"e3", x"e5", x"e4", x"e6", x"e4", x"e0", x"e1", 
        x"e5", x"e0", x"dd", x"ec", x"e6", x"e4", x"e5", x"e6", x"e6", x"e4", x"dd", x"df", x"e4", x"e6", x"e7", 
        x"e4", x"e3", x"e5", x"e8", x"ea", x"e4", x"e6", x"e5", x"e3", x"e4", x"e4", x"e5", x"e5", x"e6", x"e7", 
        x"e9", x"e6", x"e5", x"e4", x"e7", x"e6", x"e7", x"e7", x"e4", x"e7", x"e4", x"e5", x"e6", x"e5", x"e4", 
        x"e2", x"e3", x"e5", x"e1", x"e4", x"e4", x"e5", x"e8", x"e9", x"eb", x"e8", x"e7", x"e7", x"e3", x"e0", 
        x"e3", x"e9", x"e7", x"e4", x"e2", x"e3", x"e5", x"e9", x"ea", x"ec", x"ec", x"e5", x"e2", x"e5", x"e8", 
        x"eb", x"e9", x"e8", x"e9", x"ee", x"eb", x"e7", x"ea", x"eb", x"e7", x"e8", x"ee", x"e8", x"e3", x"e7", 
        x"e7", x"eb", x"e7", x"e8", x"e9", x"e6", x"e6", x"e8", x"ec", x"e9", x"e7", x"e8", x"e7", x"e8", x"ec", 
        x"ec", x"e9", x"e8", x"e8", x"e6", x"e5", x"e9", x"ec", x"e8", x"e9", x"e8", x"eb", x"ec", x"ed", x"eb", 
        x"e4", x"d5", x"e0", x"e6", x"e8", x"e7", x"e9", x"e6", x"e7", x"e9", x"e9", x"e6", x"e5", x"e8", x"e9", 
        x"e5", x"e7", x"eb", x"ea", x"e4", x"e6", x"ef", x"ec", x"eb", x"eb", x"e8", x"e8", x"e9", x"ea", x"e8", 
        x"e7", x"eb", x"ee", x"ec", x"e9", x"e9", x"eb", x"ed", x"ea", x"e8", x"ec", x"ec", x"e4", x"e9", x"ec", 
        x"ea", x"ec", x"e8", x"e5", x"e4", x"ea", x"eb", x"e7", x"e7", x"ea", x"ea", x"e7", x"e8", x"ea", x"e9", 
        x"e6", x"e6", x"e7", x"e8", x"e5", x"e2", x"ea", x"ee", x"ec", x"ea", x"e9", x"ec", x"ed", x"ed", x"eb", 
        x"ec", x"ee", x"ec", x"e9", x"eb", x"ed", x"ee", x"ed", x"ec", x"eb", x"e9", x"ea", x"eb", x"ec", x"e9", 
        x"e9", x"eb", x"eb", x"ea", x"e8", x"ec", x"ec", x"e9", x"eb", x"ed", x"ed", x"ed", x"eb", x"ed", x"f1", 
        x"ef", x"ec", x"ea", x"ed", x"ef", x"f0", x"ef", x"ee", x"ec", x"e9", x"eb", x"ea", x"ee", x"f0", x"f0", 
        x"ee", x"ec", x"e6", x"e6", x"ea", x"ec", x"eb", x"e9", x"e9", x"eb", x"ef", x"ee", x"ec", x"eb", x"eb", 
        x"e7", x"e5", x"e8", x"e0", x"ea", x"ee", x"e9", x"e9", x"ee", x"eb", x"ea", x"e8", x"e8", x"eb", x"ee", 
        x"ed", x"ec", x"e8", x"e9", x"ea", x"eb", x"ed", x"eb", x"e8", x"e8", x"e8", x"ee", x"ed", x"ed", x"ec", 
        x"ec", x"ec", x"eb", x"ea", x"ec", x"ee", x"ef", x"ed", x"ea", x"ed", x"ea", x"ea", x"ec", x"eb", x"e9", 
        x"ef", x"f0", x"ef", x"ef", x"ec", x"ec", x"ed", x"ed", x"ec", x"eb", x"eb", x"f0", x"ed", x"ea", x"ec", 
        x"ec", x"ec", x"ec", x"ed", x"ed", x"ee", x"ef", x"ed", x"ec", x"ee", x"ee", x"ec", x"ec", x"ed", x"ec", 
        x"ed", x"e9", x"dd", x"ee", x"ef", x"f2", x"f1", x"f0", x"ee", x"ed", x"ee", x"ef", x"f0", x"ee", x"ec", 
        x"ec", x"ee", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"f1", x"ed", 
        x"ee", x"ef", x"f0", x"ef", x"ef", x"f2", x"ef", x"ef", x"f5", x"f5", x"f5", x"f7", x"f3", x"ed", x"ed", 
        x"f0", x"ef", x"ee", x"f0", x"ef", x"eb", x"ee", x"f1", x"ee", x"ed", x"f1", x"f0", x"f1", x"ef", x"ef", 
        x"ee", x"ee", x"ec", x"ee", x"eb", x"e6", x"ef", x"ef", x"ee", x"ef", x"f0", x"ee", x"ef", x"f1", x"f0", 
        x"ee", x"ee", x"ec", x"eb", x"ec", x"ee", x"f2", x"f0", x"ee", x"f0", x"f0", x"f1", x"ef", x"f0", x"f3", 
        x"f7", x"f8", x"f3", x"f1", x"ef", x"f0", x"f2", x"ef", x"ec", x"ef", x"ef", x"f0", x"f1", x"ee", x"eb", 
        x"ea", x"eb", x"ec", x"ec", x"ee", x"ef", x"ef", x"ee", x"ee", x"ee", x"eb", x"ec", x"ee", x"ed", x"e7", 
        x"ed", x"ed", x"ef", x"ef", x"f0", x"e8", x"ef", x"f1", x"f1", x"f0", x"ed", x"ee", x"f1", x"f3", x"ee", 
        x"ed", x"ef", x"f2", x"f3", x"f3", x"f1", x"ed", x"ee", x"ef", x"f0", x"ef", x"f0", x"f1", x"f2", x"f3", 
        x"f1", x"f2", x"ec", x"ed", x"eb", x"f0", x"f0", x"e9", x"e8", x"e6", x"cb", x"9c", x"99", x"85", x"76", 
        x"a3", x"ae", x"7e", x"84", x"7b", x"88", x"bd", x"ba", x"9c", x"6d", x"69", x"64", x"65", x"70", x"73", 
        x"6e", x"73", x"80", x"72", x"66", x"8b", x"c5", x"c9", x"9d", x"72", x"4d", x"54", x"5b", x"52", x"53", 
        x"47", x"47", x"46", x"49", x"56", x"59", x"68", x"6a", x"64", x"68", x"6a", x"7f", x"67", x"34", x"34", 
        x"24", x"1a", x"1b", x"1a", x"0b", x"04", x"04", x"05", x"09", x"2f", x"9a", x"d1", x"d2", x"9f", x"1b", 
        x"18", x"14", x"08", x"08", x"05", x"04", x"06", x"04", x"09", x"08", x"03", x"07", x"11", x"0d", x"0c", 
        x"23", x"44", x"2a", x"0c", x"0b", x"0a", x"0c", x"0f", x"0c", x"05", x"05", x"05", x"04", x"07", x"0a", 
        x"22", x"3b", x"32", x"3b", x"4a", x"5e", x"91", x"b8", x"c7", x"c8", x"c8", x"c2", x"ae", x"87", x"8d", 
        x"c8", x"a3", x"67", x"6d", x"6a", x"67", x"6d", x"72", x"6b", x"69", x"64", x"5f", x"5f", x"4e", x"48", 
        x"57", x"4f", x"47", x"44", x"40", x"44", x"43", x"3c", x"27", x"6a", x"a6", x"68", x"85", x"b4", x"8b", 
        x"38", x"67", x"ae", x"6d", x"31", x"31", x"2c", x"29", x"29", x"1c", x"12", x"17", x"2b", x"1b", x"0f", 
        x"13", x"1b", x"40", x"2d", x"46", x"74", x"b3", x"bb", x"bb", x"b6", x"47", x"19", x"30", x"1f", x"1a", 
        x"14", x"0a", x"05", x"05", x"19", x"18", x"08", x"06", x"07", x"04", x"02", x"03", x"1c", x"2f", x"0f", 
        x"47", x"4b", x"44", x"8f", x"c1", x"64", x"34", x"3a", x"2f", x"34", x"37", x"36", x"38", x"33", x"32", 
        x"2d", x"2e", x"29", x"82", x"d6", x"c2", x"c9", x"e1", x"cf", x"c9", x"d4", x"e3", x"e3", x"e4", x"df", 
        x"e1", x"df", x"e2", x"dd", x"d4", x"e0", x"df", x"e3", x"e1", x"e3", x"e3", x"e6", x"e5", x"e4", x"e3", 
        x"e4", x"e4", x"e2", x"e4", x"e3", x"e7", x"e6", x"e2", x"e5", x"e8", x"e3", x"e4", x"e8", x"e7", x"e4", 
        x"e8", x"e9", x"e7", x"e8", x"e6", x"e2", x"e4", x"e4", x"e2", x"e3", x"e3", x"e4", x"e4", x"e6", x"e6", 
        x"e9", x"e9", x"e9", x"e5", x"ea", x"e6", x"e8", x"e6", x"e3", x"e9", x"e8", x"e6", x"e7", x"e8", x"e8", 
        x"e6", x"e5", x"e4", x"e6", x"e7", x"e3", x"da", x"da", x"e3", x"e8", x"e8", x"e6", x"e4", x"e4", x"e5", 
        x"e9", x"e7", x"e1", x"e2", x"df", x"e2", x"e7", x"eb", x"ea", x"ea", x"e7", x"e9", x"e7", x"e8", x"e9", 
        x"ec", x"ea", x"e5", x"e8", x"e8", x"e5", x"e8", x"eb", x"ea", x"eb", x"e9", x"e9", x"e9", x"e5", x"e9", 
        x"e9", x"eb", x"e9", x"eb", x"eb", x"e6", x"e6", x"ea", x"eb", x"e9", x"ea", x"e9", x"e7", x"ea", x"ee", 
        x"eb", x"e9", x"eb", x"ea", x"e7", x"e8", x"e9", x"ea", x"ea", x"e9", x"ea", x"e4", x"df", x"ea", x"eb", 
        x"e9", x"e4", x"e8", x"e8", x"eb", x"e9", x"e7", x"e6", x"e9", x"e7", x"e9", x"e9", x"e1", x"e6", x"ec", 
        x"e9", x"ea", x"eb", x"e8", x"e6", x"e6", x"ea", x"e6", x"e8", x"ea", x"e9", x"e7", x"e8", x"e9", x"e9", 
        x"e7", x"e7", x"e9", x"e7", x"e8", x"ea", x"ea", x"e8", x"e6", x"e8", x"ec", x"ee", x"ec", x"ea", x"eb", 
        x"eb", x"eb", x"e6", x"e7", x"e7", x"e8", x"e9", x"e4", x"e4", x"e9", x"eb", x"eb", x"eb", x"ed", x"eb", 
        x"e7", x"e7", x"e9", x"ed", x"e8", x"e8", x"ea", x"ea", x"ec", x"ec", x"e9", x"e9", x"ea", x"e8", x"e9", 
        x"eb", x"ec", x"ea", x"e6", x"e9", x"eb", x"ec", x"ec", x"eb", x"ec", x"ee", x"ed", x"eb", x"ec", x"ec", 
        x"e9", x"e7", x"ea", x"ec", x"ea", x"ee", x"ec", x"e9", x"eb", x"ec", x"ed", x"eb", x"e8", x"e9", x"ee", 
        x"ee", x"ec", x"ec", x"ec", x"ed", x"ed", x"ec", x"eb", x"ec", x"ef", x"ed", x"ec", x"eb", x"ec", x"ec", 
        x"eb", x"e9", x"e7", x"e9", x"ec", x"eb", x"e7", x"e7", x"ec", x"ed", x"ec", x"ec", x"ed", x"ed", x"ed", 
        x"ee", x"ed", x"e7", x"e0", x"e9", x"ed", x"ea", x"e9", x"eb", x"ec", x"ec", x"e8", x"ea", x"ec", x"eb", 
        x"ec", x"ee", x"e9", x"ea", x"ea", x"ea", x"ee", x"ee", x"eb", x"e9", x"eb", x"ed", x"ee", x"ed", x"ee", 
        x"ed", x"ea", x"e9", x"eb", x"ef", x"f0", x"ee", x"eb", x"ec", x"ee", x"ec", x"ec", x"ee", x"ef", x"ee", 
        x"ef", x"f1", x"f1", x"f0", x"ef", x"f0", x"f0", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ed", x"ea", 
        x"ea", x"ea", x"eb", x"eb", x"eb", x"eb", x"ee", x"ee", x"ed", x"ee", x"ee", x"ea", x"e8", x"e9", x"ea", 
        x"ec", x"e9", x"dd", x"ec", x"ec", x"ef", x"f0", x"ee", x"ec", x"ed", x"ee", x"ed", x"ed", x"f0", x"ec", 
        x"eb", x"ef", x"ef", x"ed", x"ec", x"ed", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"eb", 
        x"f0", x"f2", x"f2", x"f1", x"ef", x"f1", x"ee", x"ef", x"f5", x"f3", x"f0", x"f3", x"f3", x"f1", x"f1", 
        x"ef", x"eb", x"ed", x"f2", x"ef", x"ee", x"ef", x"f0", x"ee", x"ed", x"ee", x"ee", x"f1", x"ef", x"ed", 
        x"ed", x"ee", x"eb", x"ee", x"ec", x"e6", x"ef", x"f0", x"ef", x"f0", x"f0", x"ee", x"ef", x"f1", x"f1", 
        x"ee", x"ee", x"ec", x"ec", x"ee", x"ee", x"f1", x"f0", x"ee", x"ef", x"ef", x"f1", x"f0", x"f0", x"f4", 
        x"f7", x"f6", x"f4", x"f1", x"f0", x"f0", x"f0", x"ed", x"eb", x"ee", x"ed", x"ed", x"ef", x"ee", x"ec", 
        x"ed", x"ef", x"ef", x"ee", x"ee", x"ef", x"ef", x"ee", x"ee", x"ef", x"eb", x"eb", x"ee", x"ed", x"e6", 
        x"ee", x"ee", x"ef", x"ee", x"ee", x"eb", x"ee", x"eb", x"ee", x"ed", x"f1", x"ee", x"ef", x"f1", x"ee", 
        x"ef", x"f0", x"f2", x"f4", x"f4", x"f1", x"ed", x"f0", x"f1", x"f1", x"f0", x"f0", x"f0", x"ef", x"ef", 
        x"ee", x"ed", x"ef", x"ef", x"e8", x"d8", x"ad", x"8a", x"7f", x"79", x"72", x"92", x"ba", x"ae", x"7b", 
        x"91", x"94", x"7a", x"67", x"56", x"51", x"a7", x"90", x"44", x"41", x"48", x"3e", x"37", x"3c", x"3b", 
        x"36", x"4f", x"89", x"78", x"6b", x"95", x"9c", x"70", x"55", x"4b", x"29", x"1d", x"1e", x"1a", x"22", 
        x"1a", x"1f", x"1d", x"34", x"50", x"5a", x"74", x"76", x"65", x"67", x"66", x"7c", x"6c", x"24", x"2d", 
        x"23", x"1a", x"20", x"1f", x"0b", x"05", x"04", x"07", x"08", x"23", x"92", x"e0", x"e2", x"a5", x"1b", 
        x"19", x"18", x"09", x"0a", x"22", x"35", x"35", x"33", x"3a", x"3d", x"3a", x"40", x"55", x"4e", x"40", 
        x"3f", x"50", x"50", x"48", x"45", x"43", x"45", x"47", x"3c", x"27", x"1c", x"11", x"39", x"6c", x"62", 
        x"53", x"4a", x"42", x"33", x"61", x"73", x"5e", x"83", x"b0", x"c6", x"d0", x"c8", x"af", x"8c", x"92", 
        x"c9", x"a3", x"41", x"2d", x"2a", x"31", x"37", x"2a", x"2c", x"2a", x"25", x"25", x"29", x"3a", x"40", 
        x"4a", x"33", x"16", x"0d", x"0b", x"0c", x"10", x"0d", x"0d", x"2e", x"4c", x"62", x"96", x"af", x"73", 
        x"35", x"3a", x"4e", x"32", x"10", x"0a", x"0a", x"0c", x"0f", x"0c", x"0b", x"13", x"34", x"1f", x"07", 
        x"0c", x"15", x"4c", x"28", x"31", x"48", x"70", x"b1", x"c6", x"ac", x"41", x"1b", x"3c", x"1c", x"1b", 
        x"20", x"1d", x"1a", x"14", x"24", x"27", x"1a", x"19", x"1e", x"20", x"22", x"2a", x"43", x"59", x"45", 
        x"39", x"39", x"36", x"87", x"b4", x"57", x"33", x"37", x"2c", x"2d", x"2f", x"30", x"2d", x"27", x"2b", 
        x"2f", x"2c", x"21", x"84", x"dd", x"c8", x"ce", x"df", x"cf", x"cb", x"d6", x"e3", x"e0", x"e1", x"e0", 
        x"e2", x"df", x"de", x"e3", x"e1", x"df", x"e3", x"e8", x"e7", x"e7", x"e6", x"e8", x"e5", x"e4", x"e6", 
        x"e2", x"e3", x"e4", x"df", x"de", x"e1", x"e4", x"e0", x"e1", x"e9", x"ea", x"ea", x"e7", x"e8", x"e8", 
        x"eb", x"e3", x"db", x"e3", x"e5", x"e3", x"e2", x"e4", x"e4", x"e4", x"e3", x"e5", x"e5", x"e7", x"e4", 
        x"e5", x"e8", x"ea", x"e6", x"e8", x"e3", x"e7", x"e5", x"e2", x"e5", x"e6", x"e7", x"e8", x"e8", x"e3", 
        x"e5", x"e8", x"ec", x"ea", x"e5", x"e2", x"d6", x"d6", x"e2", x"e7", x"e6", x"e2", x"e4", x"e5", x"e5", 
        x"e8", x"e2", x"e0", x"e6", x"e2", x"e6", x"eb", x"ea", x"e6", x"e5", x"e3", x"e9", x"e6", x"e6", x"e9", 
        x"e8", x"e5", x"e8", x"e9", x"e4", x"e5", x"ec", x"ea", x"e6", x"ee", x"ee", x"e8", x"ec", x"e7", x"e9", 
        x"e6", x"e8", x"e7", x"eb", x"eb", x"e5", x"e7", x"eb", x"ea", x"e7", x"eb", x"ed", x"ea", x"ed", x"ee", 
        x"e8", x"ea", x"e6", x"e6", x"eb", x"ed", x"e9", x"eb", x"ed", x"ea", x"eb", x"df", x"d6", x"e8", x"ec", 
        x"ec", x"e8", x"ed", x"eb", x"e9", x"ed", x"e9", x"e6", x"e8", x"df", x"e5", x"ea", x"e2", x"e4", x"ea", 
        x"e9", x"ea", x"ea", x"e8", x"ea", x"e8", x"e9", x"e5", x"e5", x"e5", x"e9", x"e9", x"e8", x"e9", x"ed", 
        x"ea", x"e9", x"e8", x"e6", x"e6", x"e9", x"ed", x"e8", x"e6", x"ea", x"eb", x"eb", x"eb", x"e9", x"eb", 
        x"ed", x"ec", x"e6", x"e8", x"e4", x"e3", x"e7", x"e2", x"e4", x"e8", x"eb", x"ed", x"ec", x"eb", x"e9", 
        x"e7", x"e6", x"e8", x"ec", x"e9", x"eb", x"ec", x"e7", x"ea", x"eb", x"e9", x"ec", x"e9", x"e7", x"e9", 
        x"eb", x"eb", x"eb", x"e8", x"ea", x"ec", x"eb", x"eb", x"eb", x"eb", x"ef", x"ee", x"ec", x"ed", x"eb", 
        x"e9", x"e9", x"e9", x"ec", x"ee", x"ef", x"ec", x"e9", x"e9", x"e9", x"ec", x"ed", x"e9", x"ea", x"ed", 
        x"ed", x"ed", x"ee", x"ed", x"ea", x"e9", x"ea", x"ec", x"ee", x"f0", x"ee", x"ee", x"eb", x"eb", x"ec", 
        x"ee", x"ec", x"ea", x"e9", x"ec", x"ed", x"eb", x"e9", x"e9", x"ea", x"ec", x"ed", x"ee", x"ed", x"eb", 
        x"ee", x"ee", x"e6", x"df", x"e7", x"ec", x"ec", x"ea", x"e9", x"ed", x"ec", x"e9", x"ec", x"eb", x"e7", 
        x"ea", x"ec", x"ea", x"ea", x"ea", x"ea", x"eb", x"ea", x"eb", x"e9", x"eb", x"ea", x"eb", x"eb", x"ec", 
        x"ed", x"eb", x"ea", x"ea", x"eb", x"ec", x"ee", x"ed", x"ec", x"ed", x"ec", x"ec", x"ee", x"f0", x"ef", 
        x"ec", x"ee", x"ef", x"ed", x"ee", x"f0", x"f0", x"ee", x"ee", x"f0", x"f0", x"eb", x"ec", x"ed", x"eb", 
        x"ea", x"eb", x"ed", x"ed", x"ec", x"eb", x"ee", x"ed", x"ec", x"ee", x"ee", x"ea", x"e8", x"e9", x"ea", 
        x"ee", x"ec", x"e0", x"ed", x"ec", x"ee", x"ed", x"ec", x"eb", x"ec", x"ed", x"eb", x"eb", x"f1", x"ef", 
        x"ef", x"f0", x"ee", x"ed", x"ee", x"ee", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"f0", x"f0", x"ee", 
        x"f2", x"f4", x"f1", x"ef", x"ef", x"f2", x"f1", x"f2", x"f6", x"f3", x"f0", x"f1", x"f2", x"f0", x"f1", 
        x"f0", x"ed", x"f0", x"f4", x"ef", x"f0", x"ef", x"ed", x"ee", x"ee", x"eb", x"eb", x"ed", x"ee", x"ec", 
        x"ee", x"f0", x"ee", x"f0", x"ec", x"e6", x"ef", x"f0", x"f0", x"f2", x"f1", x"ef", x"ef", x"f1", x"f1", 
        x"ef", x"ef", x"ee", x"ef", x"f0", x"ee", x"f0", x"f0", x"ef", x"ef", x"ef", x"f2", x"f0", x"f0", x"f5", 
        x"f6", x"f3", x"f2", x"ef", x"ee", x"ef", x"ee", x"ee", x"ee", x"ed", x"eb", x"ec", x"ed", x"ed", x"ed", 
        x"ee", x"f1", x"f0", x"ee", x"ed", x"ed", x"ed", x"ed", x"ee", x"ef", x"eb", x"ec", x"ed", x"ec", x"e6", 
        x"ef", x"ee", x"ec", x"ef", x"f2", x"ef", x"ef", x"ee", x"f1", x"ea", x"ef", x"f0", x"f0", x"f1", x"f0", 
        x"f1", x"f0", x"f2", x"f4", x"f3", x"f0", x"ef", x"ef", x"f0", x"f1", x"f1", x"f1", x"f1", x"f1", x"f0", 
        x"ed", x"ec", x"f1", x"ec", x"e7", x"b1", x"58", x"3c", x"32", x"2d", x"2f", x"60", x"84", x"8e", x"76", 
        x"96", x"a1", x"88", x"45", x"33", x"76", x"c2", x"95", x"1b", x"1a", x"26", x"2c", x"18", x"16", x"16", 
        x"10", x"33", x"69", x"51", x"77", x"aa", x"84", x"53", x"64", x"6b", x"3c", x"22", x"24", x"2d", x"32", 
        x"2d", x"35", x"39", x"42", x"4a", x"5e", x"77", x"73", x"5c", x"63", x"63", x"72", x"7b", x"4e", x"5d", 
        x"5d", x"59", x"60", x"5e", x"21", x"04", x"06", x"06", x"07", x"1a", x"64", x"b5", x"c2", x"8c", x"16", 
        x"19", x"19", x"0b", x"0e", x"42", x"5e", x"58", x"4f", x"52", x"4f", x"50", x"4b", x"4b", x"4b", x"47", 
        x"3b", x"35", x"3a", x"41", x"3c", x"30", x"2f", x"36", x"3c", x"3e", x"3d", x"4c", x"8a", x"c5", x"c1", 
        x"bd", x"b5", x"a7", x"59", x"a7", x"c8", x"91", x"80", x"90", x"8c", x"96", x"b0", x"ad", x"8c", x"93", 
        x"bd", x"9f", x"2e", x"0a", x"08", x"20", x"30", x"08", x"07", x"08", x"09", x"16", x"18", x"26", x"22", 
        x"2f", x"25", x"1b", x"0d", x"09", x"0d", x"10", x"0a", x"09", x"0e", x"16", x"61", x"a7", x"bd", x"65", 
        x"1e", x"1d", x"14", x"13", x"24", x"34", x"38", x"3a", x"37", x"36", x"3d", x"41", x"55", x"45", x"31", 
        x"35", x"3c", x"68", x"4e", x"45", x"4b", x"4e", x"82", x"c3", x"af", x"58", x"46", x"66", x"55", x"57", 
        x"5a", x"5d", x"5e", x"54", x"5c", x"66", x"5d", x"59", x"5e", x"5e", x"59", x"5d", x"68", x"6e", x"68", 
        x"39", x"30", x"37", x"9d", x"c1", x"59", x"2e", x"2d", x"31", x"2e", x"32", x"36", x"41", x"47", x"43", 
        x"40", x"3b", x"2e", x"8d", x"dc", x"c9", x"cf", x"dc", x"cf", x"c9", x"d0", x"df", x"dd", x"e2", x"e2", 
        x"e0", x"e1", x"de", x"df", x"e1", x"e2", x"e4", x"e7", x"e4", x"e5", x"e3", x"e3", x"e0", x"e2", x"e2", 
        x"e2", x"e7", x"e6", x"dc", x"da", x"e4", x"e7", x"de", x"db", x"e0", x"e5", x"e8", x"e7", x"e8", x"e2", 
        x"e4", x"de", x"da", x"e4", x"e4", x"e3", x"e0", x"e4", x"e7", x"e6", x"e4", x"e7", x"e5", x"e4", x"e5", 
        x"e7", x"e5", x"e5", x"e5", x"e9", x"e7", x"ea", x"e6", x"e3", x"e3", x"e7", x"e3", x"e5", x"e9", x"e4", 
        x"e6", x"e7", x"e6", x"e5", x"e6", x"e8", x"e3", x"e0", x"e6", x"e7", x"e6", x"e9", x"e9", x"e2", x"e0", 
        x"e4", x"e2", x"e5", x"e5", x"e1", x"e5", x"e9", x"e6", x"e5", x"e9", x"e6", x"ed", x"e9", x"e8", x"e9", 
        x"e9", x"eb", x"e8", x"e7", x"e9", x"ea", x"eb", x"ec", x"e7", x"ec", x"ea", x"e6", x"ea", x"e6", x"e6", 
        x"e3", x"e5", x"e2", x"e7", x"ea", x"e5", x"e9", x"ec", x"e9", x"e5", x"ea", x"ec", x"ea", x"ea", x"e7", 
        x"e3", x"ea", x"e2", x"e1", x"ea", x"e9", x"e6", x"e9", x"ed", x"e7", x"e6", x"e5", x"e0", x"e7", x"e7", 
        x"ea", x"e7", x"ee", x"ed", x"ec", x"f1", x"f0", x"e8", x"e3", x"d9", x"e0", x"ea", x"e6", x"e7", x"e9", 
        x"e8", x"e7", x"e9", x"eb", x"ea", x"e5", x"e9", x"e7", x"e5", x"e2", x"e7", x"e8", x"e7", x"e6", x"ee", 
        x"ed", x"ea", x"e9", x"e7", x"e7", x"e8", x"ed", x"e8", x"e7", x"ec", x"eb", x"e8", x"e8", x"e9", x"ec", 
        x"ec", x"ed", x"e6", x"e6", x"e1", x"e1", x"e9", x"e2", x"e5", x"e9", x"ea", x"ec", x"ea", x"e8", x"e7", 
        x"ea", x"e8", x"e8", x"e9", x"e9", x"ec", x"ea", x"e4", x"ed", x"ef", x"ea", x"eb", x"ea", x"e8", x"eb", 
        x"ec", x"ea", x"eb", x"e9", x"e9", x"e8", x"ea", x"ec", x"ec", x"ec", x"ef", x"ee", x"eb", x"ed", x"eb", 
        x"ea", x"eb", x"e8", x"e9", x"ec", x"ed", x"eb", x"ec", x"e9", x"e8", x"ec", x"ee", x"ec", x"ec", x"ee", 
        x"ed", x"ed", x"ee", x"ed", x"ea", x"eb", x"ee", x"ee", x"eb", x"ea", x"ed", x"f0", x"ea", x"e8", x"e9", 
        x"ea", x"e8", x"e9", x"e8", x"e7", x"e8", x"e9", x"ea", x"e9", x"e6", x"e5", x"ea", x"ee", x"ec", x"ea", 
        x"ec", x"ee", x"e7", x"dd", x"e6", x"ee", x"ee", x"eb", x"e9", x"ec", x"ec", x"eb", x"ec", x"ea", x"e9", 
        x"ea", x"e8", x"e9", x"ea", x"eb", x"eb", x"ea", x"e9", x"ea", x"e8", x"ee", x"ed", x"ee", x"ec", x"ed", 
        x"ec", x"ed", x"ee", x"ef", x"ee", x"ed", x"ec", x"eb", x"ec", x"eb", x"eb", x"ec", x"ed", x"ed", x"ee", 
        x"ec", x"ed", x"ef", x"ec", x"ee", x"f0", x"ef", x"ef", x"ee", x"f0", x"f1", x"eb", x"ec", x"ec", x"ed", 
        x"ee", x"ee", x"ef", x"ef", x"ed", x"ed", x"ee", x"ed", x"ec", x"ef", x"ef", x"ed", x"ec", x"ed", x"ee", 
        x"f2", x"f0", x"e3", x"f0", x"ef", x"f0", x"ed", x"ec", x"ed", x"ee", x"ee", x"ed", x"ed", x"f0", x"ef", 
        x"f0", x"f0", x"ed", x"ed", x"ef", x"ee", x"ee", x"ee", x"ee", x"ef", x"ef", x"ef", x"f0", x"f1", x"ee", 
        x"f3", x"f4", x"f2", x"f1", x"f2", x"f4", x"f3", x"f5", x"f5", x"f4", x"f4", x"f3", x"f0", x"ef", x"ee", 
        x"ef", x"f0", x"f2", x"f2", x"ed", x"ef", x"ed", x"ec", x"ef", x"f0", x"ed", x"ed", x"ed", x"f0", x"ee", 
        x"f1", x"f0", x"ef", x"ef", x"ea", x"e4", x"ed", x"ee", x"ef", x"f1", x"f2", x"f0", x"ef", x"f0", x"f0", 
        x"ef", x"f0", x"ef", x"f1", x"f1", x"ee", x"f0", x"f1", x"ef", x"f0", x"f1", x"f3", x"f0", x"ef", x"f5", 
        x"f6", x"f1", x"ef", x"ed", x"ed", x"ef", x"ed", x"ed", x"ee", x"e9", x"e9", x"eb", x"ed", x"ef", x"ef", 
        x"ef", x"ef", x"ef", x"ed", x"ee", x"ef", x"ef", x"ef", x"ef", x"ed", x"eb", x"ed", x"eb", x"ec", x"e8", 
        x"ed", x"ec", x"f4", x"d4", x"a2", x"91", x"a9", x"ce", x"e9", x"f0", x"ef", x"f3", x"f2", x"f1", x"f2", 
        x"f2", x"f1", x"f2", x"f4", x"f1", x"ee", x"ee", x"ed", x"ed", x"ef", x"ef", x"ef", x"ef", x"ed", x"ee", 
        x"ec", x"ec", x"f1", x"ec", x"f0", x"ba", x"4f", x"33", x"36", x"32", x"41", x"40", x"2d", x"48", x"70", 
        x"94", x"af", x"9e", x"63", x"8b", x"cb", x"e6", x"bc", x"50", x"56", x"5f", x"69", x"65", x"61", x"67", 
        x"69", x"76", x"7f", x"52", x"6a", x"92", x"70", x"57", x"5c", x"5b", x"71", x"79", x"79", x"7f", x"75", 
        x"74", x"76", x"66", x"53", x"42", x"63", x"79", x"71", x"53", x"5e", x"64", x"69", x"7a", x"5b", x"59", 
        x"56", x"58", x"60", x"54", x"23", x"04", x"05", x"07", x"0d", x"0e", x"33", x"9f", x"bb", x"83", x"14", 
        x"14", x"15", x"0b", x"0d", x"34", x"2e", x"34", x"2d", x"24", x"28", x"43", x"35", x"19", x"25", x"28", 
        x"23", x"1b", x"13", x"0f", x"09", x"04", x"06", x"20", x"30", x"23", x"5b", x"95", x"ac", x"c0", x"c5", 
        x"d3", x"dd", x"a6", x"64", x"b9", x"ce", x"bd", x"a7", x"bb", x"b8", x"9d", x"8c", x"88", x"8e", x"9e", 
        x"cf", x"ac", x"30", x"0a", x"0d", x"34", x"4e", x"1a", x"15", x"14", x"0e", x"0e", x"17", x"20", x"0c", 
        x"0e", x"1d", x"38", x"33", x"2b", x"2e", x"30", x"25", x"13", x"19", x"35", x"55", x"81", x"a3", x"6a", 
        x"1c", x"1c", x"36", x"2c", x"51", x"7d", x"76", x"72", x"6c", x"67", x"6b", x"69", x"68", x"61", x"5a", 
        x"54", x"5c", x"6b", x"67", x"5e", x"6b", x"a0", x"89", x"99", x"b7", x"63", x"40", x"41", x"48", x"49", 
        x"45", x"43", x"3e", x"37", x"46", x"51", x"43", x"38", x"38", x"36", x"33", x"32", x"27", x"21", x"24", 
        x"3f", x"23", x"3b", x"a4", x"a9", x"53", x"4f", x"45", x"4b", x"31", x"28", x"35", x"4c", x"4b", x"46", 
        x"46", x"4b", x"3e", x"93", x"e1", x"ca", x"ce", x"df", x"ce", x"c7", x"d1", x"e3", x"de", x"df", x"e1", 
        x"e2", x"e8", x"e5", x"e2", x"e6", x"e9", x"e4", x"e3", x"df", x"df", x"df", x"e2", x"e1", x"e8", x"e6", 
        x"e6", x"e4", x"e4", x"e2", x"dd", x"e5", x"e9", x"e2", x"e4", x"e4", x"e3", x"e9", x"e8", x"e5", x"e3", 
        x"e7", x"e4", x"e1", x"e8", x"e6", x"e4", x"df", x"e2", x"e6", x"e3", x"df", x"e2", x"e2", x"e2", x"e2", 
        x"e3", x"e3", x"e6", x"e4", x"e7", x"e6", x"e7", x"e3", x"e2", x"e4", x"e9", x"e4", x"e7", x"eb", x"e3", 
        x"e2", x"e2", x"df", x"e2", x"e7", x"e7", x"e8", x"e6", x"e7", x"e6", x"e4", x"e9", x"e7", x"e0", x"e1", 
        x"e4", x"e2", x"e5", x"e6", x"e4", x"e9", x"eb", x"e6", x"e5", x"e9", x"e6", x"ee", x"ec", x"ea", x"e5", 
        x"e2", x"e9", x"ea", x"e4", x"e7", x"e8", x"e9", x"ed", x"dc", x"de", x"e1", x"e4", x"e8", x"e7", x"e9", 
        x"e9", x"e9", x"df", x"e3", x"e8", x"e5", x"e8", x"ea", x"e7", x"e9", x"eb", x"ed", x"ea", x"e7", x"e7", 
        x"e6", x"ed", x"ea", x"e8", x"ea", x"e7", x"eb", x"ee", x"ec", x"e9", x"e7", x"ec", x"e8", x"e4", x"e7", 
        x"e8", x"e8", x"e8", x"e9", x"e9", x"e1", x"e8", x"ea", x"ea", x"e5", x"e7", x"ea", x"e7", x"e9", x"e9", 
        x"ea", x"eb", x"e8", x"ea", x"eb", x"e3", x"e4", x"e8", x"ea", x"e6", x"e9", x"e7", x"e5", x"e6", x"ea", 
        x"eb", x"e9", x"e7", x"e8", x"eb", x"ea", x"ec", x"e8", x"e6", x"e9", x"e9", x"e8", x"e9", x"eb", x"e8", 
        x"e6", x"eb", x"e7", x"e6", x"e6", x"e6", x"eb", x"e5", x"e7", x"ea", x"ea", x"ec", x"eb", x"e9", x"ea", 
        x"f0", x"ee", x"ec", x"ea", x"eb", x"ec", x"eb", x"e6", x"eb", x"eb", x"e9", x"eb", x"e9", x"e8", x"eb", 
        x"ec", x"eb", x"ed", x"ec", x"ea", x"e9", x"ea", x"ed", x"ed", x"eb", x"ed", x"ec", x"e9", x"ee", x"ee", 
        x"eb", x"e7", x"e8", x"ea", x"e9", x"ea", x"ea", x"ed", x"eb", x"e8", x"eb", x"ec", x"eb", x"ed", x"ed", 
        x"eb", x"eb", x"ed", x"ec", x"ec", x"ed", x"ed", x"e9", x"e7", x"e9", x"ed", x"f1", x"eb", x"ea", x"eb", 
        x"eb", x"ea", x"eb", x"eb", x"ea", x"ea", x"e9", x"e9", x"e9", x"e3", x"e0", x"e9", x"ed", x"eb", x"e9", 
        x"e8", x"eb", x"eb", x"de", x"e6", x"ef", x"ed", x"ea", x"e9", x"e9", x"eb", x"eb", x"ea", x"eb", x"ec", 
        x"ea", x"e8", x"e9", x"e9", x"eb", x"ee", x"ed", x"ee", x"eb", x"e6", x"ec", x"e9", x"ed", x"ed", x"f0", 
        x"f0", x"ec", x"eb", x"eb", x"ed", x"ec", x"ea", x"e9", x"eb", x"eb", x"eb", x"eb", x"ea", x"ea", x"ec", 
        x"ed", x"ee", x"f0", x"ec", x"ef", x"f0", x"ef", x"ee", x"ec", x"ec", x"ef", x"ea", x"eb", x"e9", x"ec", 
        x"ee", x"ee", x"ee", x"ee", x"ed", x"ed", x"ed", x"ec", x"eb", x"ed", x"ed", x"ec", x"eb", x"eb", x"ec", 
        x"ef", x"eb", x"de", x"ed", x"ed", x"f0", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ec", 
        x"ec", x"ef", x"ef", x"ee", x"ed", x"ed", x"ed", x"ee", x"ee", x"ee", x"ef", x"ef", x"f2", x"f3", x"f0", 
        x"f3", x"f3", x"f1", x"f1", x"f1", x"ee", x"ee", x"f0", x"ef", x"f0", x"f2", x"f2", x"f1", x"f1", x"f0", 
        x"ef", x"f0", x"f1", x"f1", x"ef", x"f0", x"ee", x"ec", x"ee", x"ef", x"ee", x"f0", x"f0", x"f2", x"f0", 
        x"f0", x"ef", x"ef", x"f0", x"eb", x"e5", x"ef", x"ef", x"f0", x"f2", x"f3", x"f0", x"ef", x"f0", x"f0", 
        x"ef", x"f0", x"f0", x"f1", x"f2", x"ef", x"f1", x"f1", x"f0", x"f0", x"f3", x"f3", x"ef", x"ee", x"f3", 
        x"f5", x"f1", x"ef", x"ef", x"ef", x"ef", x"ec", x"ec", x"ed", x"eb", x"ee", x"ef", x"ef", x"ee", x"ed", 
        x"ea", x"ee", x"ee", x"ee", x"ef", x"ef", x"ee", x"ec", x"ee", x"ef", x"ee", x"ee", x"ea", x"ea", x"e7", 
        x"eb", x"ee", x"e3", x"88", x"2f", x"21", x"2b", x"48", x"9f", x"eb", x"f2", x"f2", x"f2", x"f1", x"ec", 
        x"ec", x"ee", x"f1", x"f4", x"f2", x"ef", x"f1", x"ee", x"ef", x"f3", x"f0", x"ea", x"ea", x"e7", x"e4", 
        x"e1", x"d8", x"d6", x"d2", x"ce", x"b2", x"7e", x"51", x"2f", x"21", x"21", x"1d", x"13", x"14", x"21", 
        x"2a", x"5c", x"90", x"86", x"b3", x"ce", x"e2", x"c0", x"6d", x"73", x"74", x"70", x"71", x"6d", x"71", 
        x"74", x"6e", x"63", x"39", x"29", x"2e", x"21", x"19", x"18", x"20", x"46", x"57", x"54", x"42", x"3c", 
        x"3b", x"39", x"39", x"4a", x"38", x"63", x"73", x"74", x"57", x"5c", x"67", x"6b", x"6e", x"35", x"1f", 
        x"1b", x"28", x"3b", x"20", x"0e", x"03", x"03", x"04", x"0a", x"18", x"59", x"ac", x"bc", x"7f", x"12", 
        x"12", x"18", x"0d", x"15", x"38", x"20", x"29", x"23", x"17", x"20", x"42", x"36", x"15", x"1f", x"1d", 
        x"1b", x"16", x"12", x"12", x"14", x"14", x"13", x"2c", x"3a", x"26", x"77", x"aa", x"9d", x"a9", x"bb", 
        x"c6", x"ce", x"7b", x"58", x"c2", x"cd", x"bf", x"ae", x"bd", x"c8", x"c4", x"b0", x"a3", x"8a", x"89", 
        x"c8", x"b3", x"3d", x"24", x"27", x"31", x"40", x"2d", x"40", x"52", x"46", x"33", x"22", x"17", x"12", 
        x"17", x"1e", x"29", x"26", x"26", x"24", x"24", x"1d", x"15", x"16", x"1d", x"2b", x"5d", x"9b", x"84", 
        x"25", x"0b", x"1a", x"28", x"33", x"3c", x"38", x"32", x"33", x"2c", x"29", x"27", x"1f", x"20", x"21", 
        x"1a", x"1e", x"26", x"2b", x"29", x"37", x"90", x"a4", x"ab", x"a6", x"43", x"22", x"14", x"12", x"13", 
        x"13", x"13", x"11", x"1b", x"29", x"1f", x"17", x"10", x"10", x"13", x"1b", x"1e", x"0f", x"09", x"0e", 
        x"1c", x"33", x"53", x"a0", x"c4", x"6a", x"54", x"58", x"4e", x"29", x"22", x"45", x"5b", x"3a", x"3a", 
        x"37", x"36", x"34", x"87", x"e2", x"c6", x"c4", x"dd", x"c4", x"ba", x"ce", x"e3", x"dd", x"e0", x"e2", 
        x"e2", x"e5", x"ea", x"e5", x"e6", x"e3", x"e1", x"e1", x"e4", x"dc", x"e1", x"eb", x"e5", x"df", x"e5", 
        x"e5", x"e1", x"e4", x"e3", x"e1", x"e3", x"e9", x"e7", x"e5", x"e2", x"e8", x"ea", x"e7", x"e1", x"e6", 
        x"e0", x"e1", x"e6", x"e5", x"e2", x"e5", x"e2", x"e2", x"e7", x"e3", x"df", x"e0", x"e0", x"dc", x"e3", 
        x"e6", x"e3", x"e1", x"e1", x"e1", x"e0", x"e3", x"e0", x"e3", x"e8", x"e3", x"e3", x"e8", x"eb", x"e5", 
        x"dd", x"e1", x"e5", x"e6", x"e4", x"e6", x"e5", x"eb", x"e8", x"db", x"dc", x"e7", x"df", x"de", x"e7", 
        x"e5", x"e2", x"e4", x"e3", x"e4", x"e4", x"e9", x"ec", x"e9", x"e7", x"e9", x"e8", x"e6", x"e8", x"e7", 
        x"e4", x"e8", x"ea", x"e3", x"e8", x"ec", x"e9", x"eb", x"e2", x"e0", x"e4", x"e9", x"eb", x"eb", x"ec", 
        x"ee", x"eb", x"db", x"d8", x"e5", x"ea", x"ed", x"ea", x"e5", x"e3", x"e5", x"eb", x"ec", x"e6", x"e8", 
        x"e9", x"e9", x"e7", x"ed", x"ed", x"ea", x"ea", x"ec", x"e6", x"e8", x"e5", x"e4", x"ec", x"eb", x"ec", 
        x"ea", x"ea", x"eb", x"eb", x"e3", x"d3", x"e5", x"eb", x"ea", x"ea", x"ea", x"ec", x"ea", x"e7", x"e8", 
        x"ec", x"ed", x"e7", x"ec", x"e8", x"e4", x"eb", x"e9", x"ea", x"eb", x"eb", x"eb", x"ea", x"e8", x"e3", 
        x"e9", x"ea", x"e8", x"e8", x"e8", x"e5", x"e9", x"e6", x"e4", x"e6", x"e8", x"ea", x"ec", x"ea", x"ec", 
        x"eb", x"ea", x"ea", x"e5", x"e0", x"e6", x"ea", x"e5", x"e5", x"e8", x"eb", x"ec", x"ed", x"ed", x"eb", 
        x"ef", x"ed", x"ea", x"ea", x"ea", x"ea", x"eb", x"ea", x"e9", x"e9", x"eb", x"e9", x"e8", x"ea", x"eb", 
        x"ee", x"ec", x"ec", x"e9", x"ea", x"e9", x"e9", x"ea", x"ec", x"ed", x"ef", x"eb", x"e9", x"ee", x"ec", 
        x"ea", x"ea", x"eb", x"eb", x"ed", x"ef", x"ec", x"ec", x"ee", x"ec", x"ec", x"ea", x"eb", x"f1", x"eb", 
        x"e9", x"eb", x"ec", x"e9", x"e9", x"e8", x"eb", x"e7", x"e8", x"ed", x"ee", x"f0", x"ec", x"e9", x"eb", 
        x"ea", x"eb", x"ec", x"e8", x"e7", x"ec", x"ee", x"ea", x"e8", x"e8", x"e5", x"e6", x"eb", x"ee", x"ec", 
        x"e7", x"e8", x"ea", x"e1", x"e4", x"ed", x"eb", x"ee", x"ec", x"eb", x"e9", x"ea", x"ed", x"eb", x"e9", 
        x"e8", x"ec", x"ea", x"ed", x"ed", x"eb", x"eb", x"eb", x"e9", x"ec", x"ee", x"e8", x"ed", x"ea", x"e7", 
        x"e9", x"ec", x"ea", x"e8", x"e8", x"eb", x"ed", x"eb", x"ea", x"eb", x"eb", x"ea", x"e8", x"e7", x"ea", 
        x"ed", x"ed", x"ef", x"ee", x"ee", x"ef", x"ed", x"ec", x"f2", x"ed", x"ec", x"ec", x"e9", x"e9", x"ec", 
        x"ea", x"ee", x"ed", x"f0", x"ee", x"ed", x"ec", x"ec", x"ef", x"ed", x"ec", x"ec", x"ec", x"eb", x"ec", 
        x"ed", x"e7", x"db", x"ec", x"ed", x"f2", x"f0", x"f0", x"f0", x"ef", x"ee", x"ed", x"ed", x"ed", x"ee", 
        x"ec", x"f0", x"f0", x"ef", x"ee", x"ed", x"f0", x"f1", x"f0", x"f1", x"f2", x"f1", x"f1", x"f2", x"f2", 
        x"f3", x"f3", x"f2", x"f1", x"f0", x"f0", x"f1", x"f0", x"f0", x"f2", x"f1", x"ef", x"f0", x"f0", x"f0", 
        x"f1", x"f1", x"f0", x"ef", x"ef", x"f1", x"f1", x"f0", x"ee", x"ee", x"ee", x"f0", x"ee", x"f1", x"ed", 
        x"ed", x"f1", x"ef", x"ef", x"ec", x"e2", x"ed", x"ee", x"ed", x"f1", x"f1", x"f0", x"f1", x"f1", x"f0", 
        x"ef", x"f0", x"f1", x"f0", x"f0", x"f2", x"f3", x"f1", x"f0", x"f2", x"f2", x"ef", x"ef", x"f3", x"f3", 
        x"f3", x"f1", x"f1", x"ee", x"ec", x"ed", x"ef", x"ef", x"ee", x"ed", x"f1", x"f2", x"f1", x"ee", x"ef", 
        x"f1", x"ef", x"ec", x"ec", x"ef", x"ef", x"f0", x"ee", x"ec", x"ee", x"ef", x"ee", x"f0", x"ec", x"e8", 
        x"ee", x"f0", x"c0", x"47", x"16", x"15", x"26", x"58", x"95", x"e7", x"f0", x"ee", x"f0", x"f2", x"ef", 
        x"ed", x"ed", x"ed", x"f1", x"ed", x"ec", x"ee", x"ed", x"ec", x"e9", x"c2", x"9b", x"97", x"8a", x"7d", 
        x"76", x"72", x"67", x"61", x"59", x"5d", x"5b", x"36", x"1c", x"0f", x"0e", x"0e", x"0b", x"10", x"0e", 
        x"11", x"42", x"77", x"7a", x"af", x"c8", x"e0", x"b2", x"2f", x"20", x"3f", x"3a", x"25", x"21", x"25", 
        x"2a", x"18", x"15", x"0f", x"0b", x"0b", x"10", x"0e", x"0b", x"13", x"32", x"46", x"42", x"23", x"21", 
        x"20", x"1e", x"30", x"4c", x"30", x"61", x"73", x"75", x"50", x"5e", x"67", x"6b", x"6e", x"36", x"1c", 
        x"1e", x"2a", x"37", x"21", x"0d", x"07", x"04", x"03", x"05", x"1f", x"67", x"a1", x"ad", x"76", x"11", 
        x"0e", x"0d", x"0f", x"2c", x"51", x"47", x"44", x"4d", x"4d", x"5c", x"70", x"6c", x"60", x"5f", x"52", 
        x"52", x"55", x"59", x"5c", x"61", x"60", x"64", x"68", x"62", x"5e", x"85", x"ac", x"99", x"a8", x"b5", 
        x"a0", x"a5", x"7e", x"73", x"cd", x"c4", x"c3", x"a6", x"ab", x"bf", x"c3", x"b0", x"a4", x"8b", x"80", 
        x"c7", x"b4", x"36", x"15", x"17", x"0f", x"10", x"18", x"2e", x"3f", x"34", x"25", x"12", x"0b", x"0c", 
        x"0b", x"08", x"0a", x"07", x"0a", x"0a", x"06", x"06", x"06", x"05", x"06", x"18", x"45", x"77", x"7a", 
        x"34", x"0d", x"09", x"14", x"1a", x"17", x"13", x"0d", x"0d", x"0d", x"19", x"0e", x"07", x"09", x"0e", 
        x"0a", x"1f", x"53", x"67", x"64", x"47", x"46", x"5f", x"74", x"69", x"2d", x"22", x"17", x"0e", x"0d", 
        x"10", x"13", x"0c", x"17", x"25", x"13", x"0e", x"09", x"0a", x"0c", x"18", x"1a", x"11", x"0c", x"0c", 
        x"17", x"38", x"45", x"9c", x"cf", x"66", x"30", x"46", x"32", x"2e", x"3a", x"3a", x"41", x"38", x"40", 
        x"34", x"29", x"2d", x"88", x"db", x"c2", x"c9", x"dc", x"c8", x"c4", x"d5", x"e6", x"df", x"e2", x"e3", 
        x"e2", x"e2", x"e6", x"e2", x"e4", x"e4", x"e4", x"e3", x"e3", x"e1", x"e7", x"e8", x"e1", x"df", x"e7", 
        x"e9", x"df", x"df", x"e4", x"e3", x"df", x"e2", x"e2", x"e1", x"df", x"e4", x"e4", x"e2", x"e2", x"e5", 
        x"df", x"e5", x"e5", x"e1", x"e3", x"e6", x"e5", x"e4", x"e4", x"e4", x"e6", x"e0", x"e0", x"df", x"e5", 
        x"e9", x"e7", x"e1", x"df", x"e6", x"e3", x"e8", x"e3", x"e1", x"e4", x"e1", x"e4", x"df", x"dd", x"de", 
        x"e1", x"e6", x"e4", x"e7", x"e5", x"e5", x"e4", x"e8", x"e7", x"e5", x"e3", x"e9", x"ec", x"ea", x"eb", 
        x"e6", x"e7", x"e8", x"e5", x"e6", x"e3", x"e5", x"e9", x"e7", x"e7", x"eb", x"ea", x"e7", x"e9", x"eb", 
        x"ea", x"ec", x"e5", x"e1", x"e5", x"e9", x"e6", x"e8", x"ea", x"eb", x"ea", x"e9", x"e9", x"e9", x"e9", 
        x"ed", x"eb", x"e7", x"e2", x"e2", x"ea", x"e8", x"e4", x"e9", x"e8", x"e4", x"e6", x"e8", x"e5", x"e9", 
        x"eb", x"ea", x"e5", x"e9", x"ee", x"eb", x"e9", x"eb", x"e5", x"e8", x"e4", x"e1", x"ea", x"e9", x"e9", 
        x"e9", x"e7", x"e6", x"ea", x"eb", x"e6", x"e9", x"e6", x"e7", x"e8", x"e7", x"e9", x"e7", x"e5", x"ec", 
        x"eb", x"e8", x"ec", x"ef", x"eb", x"ea", x"e9", x"eb", x"ec", x"ed", x"ed", x"ed", x"eb", x"e9", x"e7", 
        x"e9", x"ea", x"e9", x"e8", x"e8", x"e8", x"ec", x"ea", x"e9", x"e9", x"ea", x"eb", x"ed", x"e9", x"e9", 
        x"eb", x"eb", x"ea", x"e7", x"e5", x"eb", x"ed", x"eb", x"ea", x"e9", x"ea", x"eb", x"eb", x"ec", x"ed", 
        x"ed", x"e8", x"e8", x"ed", x"ec", x"ea", x"eb", x"ec", x"ea", x"eb", x"ed", x"e8", x"e7", x"e9", x"e9", 
        x"ec", x"eb", x"ea", x"e7", x"ed", x"ec", x"e8", x"e8", x"ec", x"ee", x"ee", x"ec", x"e8", x"ed", x"ed", 
        x"e9", x"ec", x"ec", x"e9", x"ec", x"ee", x"ed", x"ee", x"ee", x"ed", x"ed", x"ec", x"ee", x"ee", x"e8", 
        x"eb", x"ec", x"eb", x"ed", x"eb", x"e8", x"ec", x"ea", x"ec", x"ed", x"e8", x"ec", x"eb", x"e4", x"ea", 
        x"ef", x"ed", x"ec", x"e9", x"e9", x"eb", x"ed", x"ec", x"e8", x"e8", x"e8", x"e8", x"ec", x"ee", x"eb", 
        x"e9", x"ea", x"ec", x"e1", x"e1", x"ec", x"ed", x"ee", x"ea", x"eb", x"e8", x"e8", x"ec", x"ea", x"e9", 
        x"e8", x"eb", x"e8", x"ea", x"e9", x"e8", x"e8", x"e8", x"e8", x"eb", x"ee", x"ec", x"f0", x"ee", x"ec", 
        x"ea", x"eb", x"ea", x"e9", x"e9", x"eb", x"ec", x"eb", x"eb", x"ea", x"ec", x"ec", x"ea", x"ec", x"ef", 
        x"eb", x"eb", x"ed", x"ed", x"ed", x"ec", x"ec", x"ec", x"ef", x"ea", x"eb", x"f1", x"ec", x"ec", x"f0", 
        x"ec", x"eb", x"ea", x"ee", x"ef", x"ed", x"ed", x"ed", x"ee", x"eb", x"eb", x"ea", x"e8", x"e9", x"eb", 
        x"ed", x"e8", x"dc", x"eb", x"ee", x"f2", x"f2", x"ef", x"ed", x"ec", x"ee", x"ef", x"f0", x"ef", x"f0", 
        x"ee", x"f1", x"f1", x"ef", x"ef", x"f0", x"f1", x"f0", x"ee", x"f1", x"f2", x"ef", x"f1", x"f3", x"f3", 
        x"f3", x"f3", x"f1", x"ef", x"f0", x"f2", x"f2", x"ef", x"f0", x"f1", x"ef", x"ee", x"ef", x"ef", x"ef", 
        x"f0", x"f0", x"ee", x"ed", x"ee", x"f1", x"f2", x"ef", x"ed", x"ee", x"f0", x"f0", x"ef", x"f1", x"ed", 
        x"ec", x"ef", x"ec", x"ec", x"ec", x"e3", x"ee", x"ef", x"ed", x"f0", x"f1", x"f2", x"f2", x"f2", x"f1", 
        x"f0", x"f0", x"f2", x"f3", x"f2", x"f4", x"f3", x"f1", x"f2", x"f4", x"f2", x"ef", x"f1", x"f5", x"f3", 
        x"f3", x"f2", x"f2", x"f0", x"ef", x"f0", x"f1", x"ef", x"ed", x"ee", x"f0", x"ef", x"f0", x"ef", x"ef", 
        x"ef", x"ed", x"ea", x"eb", x"ee", x"ef", x"f1", x"f1", x"ef", x"ef", x"ef", x"ed", x"f1", x"ed", x"ea", 
        x"f0", x"f1", x"b5", x"3a", x"0a", x"14", x"3b", x"9e", x"bb", x"eb", x"ee", x"f2", x"f0", x"e9", x"ed", 
        x"ea", x"eb", x"eb", x"f2", x"ed", x"ec", x"ec", x"ed", x"ea", x"b3", x"4c", x"2f", x"25", x"26", x"1e", 
        x"1b", x"1d", x"1e", x"2b", x"27", x"22", x"26", x"1b", x"0e", x"0d", x"0f", x"1b", x"28", x"0f", x"11", 
        x"0e", x"30", x"5b", x"77", x"aa", x"bd", x"dc", x"b4", x"2f", x"1e", x"43", x"48", x"2c", x"2b", x"2c", 
        x"2a", x"11", x"0f", x"0e", x"0e", x"11", x"0e", x"0d", x"0a", x"1c", x"44", x"4b", x"48", x"36", x"36", 
        x"35", x"37", x"43", x"4a", x"31", x"69", x"78", x"6f", x"40", x"54", x"64", x"69", x"73", x"70", x"6c", 
        x"6e", x"6f", x"75", x"68", x"26", x"05", x"07", x"08", x"06", x"0d", x"4b", x"a0", x"a5", x"74", x"15", 
        x"07", x"09", x"2b", x"69", x"7b", x"71", x"71", x"6a", x"68", x"79", x"6b", x"64", x"64", x"5f", x"60", 
        x"5f", x"5d", x"5e", x"5f", x"54", x"53", x"4e", x"48", x"45", x"44", x"5f", x"a6", x"a7", x"9a", x"b3", 
        x"be", x"b0", x"69", x"73", x"cf", x"c9", x"cb", x"c1", x"93", x"af", x"ca", x"bf", x"ac", x"8a", x"7b", 
        x"c4", x"b1", x"2f", x"08", x"08", x"06", x"0b", x"13", x"1b", x"29", x"21", x"0b", x"04", x"06", x"04", 
        x"03", x"05", x"06", x"07", x"04", x"08", x"03", x"07", x"08", x"05", x"04", x"10", x"36", x"54", x"3f", 
        x"26", x"2a", x"23", x"2e", x"4a", x"3b", x"1f", x"0f", x"0d", x"12", x"1e", x"17", x"0e", x"0c", x"0c", 
        x"13", x"20", x"33", x"3f", x"4c", x"55", x"51", x"49", x"50", x"4a", x"2c", x"2a", x"26", x"23", x"22", 
        x"23", x"22", x"22", x"38", x"3b", x"24", x"1e", x"1f", x"2d", x"3f", x"50", x"50", x"4b", x"3e", x"3a", 
        x"18", x"29", x"33", x"60", x"97", x"6c", x"32", x"2b", x"17", x"2f", x"42", x"35", x"2e", x"39", x"38", 
        x"2d", x"2d", x"32", x"8f", x"df", x"c5", x"d2", x"de", x"c9", x"c6", x"cc", x"dd", x"e0", x"e3", x"e1", 
        x"df", x"e0", x"e6", x"e5", x"e3", x"e1", x"e7", x"e7", x"e3", x"e3", x"e5", x"e2", x"e5", x"e0", x"e7", 
        x"e4", x"dd", x"e5", x"e9", x"e6", x"e4", x"e5", x"e4", x"e7", x"e5", x"e6", x"e4", x"e1", x"e4", x"e5", 
        x"e3", x"eb", x"e4", x"e0", x"e5", x"e7", x"e6", x"e7", x"e3", x"e4", x"ea", x"e5", x"e3", x"e6", x"e0", 
        x"dc", x"de", x"e3", x"e6", x"e2", x"e2", x"e3", x"dd", x"e1", x"da", x"df", x"e6", x"e0", x"de", x"e2", 
        x"e3", x"e6", x"e6", x"e4", x"e0", x"e1", x"e3", x"e4", x"e2", x"e3", x"e3", x"e2", x"e6", x"e9", x"ea", 
        x"e7", x"e7", x"e6", x"e8", x"e9", x"e7", x"e7", x"e9", x"ea", x"eb", x"ea", x"e9", x"e7", x"e8", x"ec", 
        x"ed", x"ee", x"e8", x"ea", x"eb", x"ea", x"e9", x"e9", x"eb", x"ee", x"eb", x"e8", x"ea", x"eb", x"e8", 
        x"e9", x"e0", x"dc", x"e2", x"e1", x"e8", x"e9", x"e6", x"ed", x"ec", x"e0", x"de", x"e4", x"e7", x"e9", 
        x"ea", x"ea", x"e7", x"e7", x"ee", x"e7", x"e6", x"ec", x"e9", x"ec", x"e9", x"e6", x"eb", x"e9", x"e9", 
        x"e9", x"e7", x"e6", x"eb", x"e9", x"ec", x"ea", x"e6", x"e8", x"e8", x"e6", x"e8", x"e7", x"e5", x"e9", 
        x"e9", x"e9", x"ea", x"e6", x"e4", x"eb", x"ec", x"ed", x"eb", x"e8", x"e7", x"e9", x"ec", x"ed", x"ea", 
        x"e9", x"ec", x"ed", x"ec", x"ea", x"ea", x"e9", x"ea", x"eb", x"eb", x"ea", x"ea", x"eb", x"e8", x"e6", 
        x"ea", x"ed", x"ea", x"e7", x"e6", x"e6", x"e8", x"ea", x"ea", x"e7", x"e7", x"e9", x"ea", x"ec", x"ee", 
        x"ea", x"e5", x"e8", x"ed", x"ec", x"ec", x"ee", x"eb", x"e6", x"e8", x"eb", x"e7", x"e8", x"ea", x"eb", 
        x"ec", x"ea", x"e9", x"e7", x"eb", x"ec", x"ec", x"ed", x"ee", x"ed", x"eb", x"ec", x"ed", x"ed", x"eb", 
        x"eb", x"eb", x"e8", x"e9", x"e9", x"ea", x"ed", x"ee", x"ee", x"ef", x"ed", x"ed", x"eb", x"eb", x"eb", 
        x"eb", x"e9", x"ec", x"ef", x"ee", x"ea", x"ec", x"e9", x"e9", x"ea", x"e3", x"e8", x"ea", x"e4", x"e9", 
        x"ee", x"ec", x"e9", x"e8", x"e8", x"ea", x"ed", x"ef", x"ed", x"eb", x"e9", x"ea", x"ed", x"ec", x"ea", 
        x"eb", x"ed", x"ed", x"e2", x"e2", x"eb", x"eb", x"ed", x"ea", x"ec", x"ea", x"e9", x"ec", x"eb", x"eb", 
        x"ea", x"e8", x"ea", x"eb", x"eb", x"ef", x"ed", x"ed", x"ea", x"e9", x"ed", x"ef", x"ee", x"ed", x"ed", 
        x"eb", x"eb", x"ec", x"eb", x"eb", x"ec", x"e9", x"ea", x"eb", x"e9", x"eb", x"ea", x"e6", x"e8", x"eb", 
        x"ec", x"ef", x"ef", x"ee", x"ec", x"ea", x"eb", x"f0", x"ee", x"e9", x"ec", x"f1", x"ed", x"ec", x"ed", 
        x"ea", x"e9", x"ea", x"ed", x"ee", x"ea", x"ec", x"ee", x"ee", x"eb", x"ec", x"ed", x"ea", x"ea", x"ea", 
        x"eb", x"ea", x"dc", x"eb", x"ee", x"f0", x"f0", x"ee", x"ed", x"ed", x"ee", x"f0", x"f0", x"ef", x"ef", 
        x"eb", x"ee", x"ee", x"ed", x"ed", x"f1", x"f1", x"ef", x"ee", x"f2", x"f4", x"f3", x"f3", x"f4", x"f4", 
        x"f4", x"f3", x"f0", x"ef", x"f0", x"f1", x"f0", x"ee", x"ef", x"f1", x"f1", x"f0", x"ef", x"ee", x"ef", 
        x"f0", x"f0", x"ef", x"ed", x"ee", x"f0", x"f1", x"ee", x"ed", x"ef", x"f1", x"f0", x"ee", x"f0", x"ed", 
        x"ee", x"ee", x"ed", x"ee", x"f0", x"e5", x"ed", x"ee", x"ed", x"ee", x"ef", x"f0", x"f1", x"f2", x"f3", 
        x"f3", x"f2", x"f3", x"f4", x"f4", x"f4", x"f2", x"f0", x"f2", x"f5", x"f3", x"f1", x"f2", x"f5", x"f3", 
        x"f3", x"f2", x"f1", x"f1", x"f1", x"f2", x"f2", x"ef", x"ed", x"ef", x"f0", x"ee", x"f1", x"f2", x"f2", 
        x"f1", x"f0", x"ee", x"ee", x"ee", x"ec", x"ed", x"ed", x"ef", x"f1", x"ee", x"eb", x"ed", x"e9", x"e4", 
        x"ec", x"f2", x"d0", x"51", x"33", x"42", x"57", x"9e", x"b0", x"ec", x"f2", x"ec", x"ef", x"f0", x"ed", 
        x"ee", x"ef", x"eb", x"e9", x"e6", x"e5", x"e4", x"e5", x"ed", x"a0", x"26", x"2f", x"2b", x"31", x"30", 
        x"2f", x"2a", x"2c", x"38", x"33", x"2e", x"2f", x"30", x"20", x"0c", x"0e", x"55", x"81", x"27", x"09", 
        x"07", x"1b", x"59", x"88", x"ac", x"ba", x"d6", x"bf", x"62", x"5e", x"6a", x"71", x"6c", x"6f", x"71", 
        x"5b", x"1a", x"0c", x"09", x"32", x"64", x"23", x"0b", x"09", x"24", x"6d", x"80", x"88", x"89", x"8d", 
        x"8b", x"7e", x"6f", x"51", x"2c", x"68", x"7a", x"74", x"3f", x"54", x"63", x"64", x"75", x"76", x"62", 
        x"60", x"59", x"56", x"59", x"3d", x"0e", x"04", x"05", x"07", x"1a", x"61", x"a4", x"ab", x"91", x"3a", 
        x"0f", x"18", x"34", x"41", x"36", x"2c", x"2f", x"24", x"1f", x"23", x"17", x"22", x"1f", x"11", x"13", 
        x"0d", x"0f", x"1b", x"32", x"20", x"20", x"19", x"14", x"15", x"0f", x"25", x"81", x"b2", x"ac", x"bb", 
        x"c0", x"98", x"50", x"6b", x"c0", x"cf", x"cc", x"d0", x"b1", x"a9", x"c4", x"c7", x"b1", x"88", x"7d", 
        x"c8", x"a6", x"27", x"05", x"06", x"07", x"09", x"13", x"1a", x"29", x"20", x"0c", x"0b", x"0c", x"0c", 
        x"0d", x"11", x"0f", x"10", x"12", x"0f", x"0e", x"17", x"13", x"14", x"13", x"11", x"13", x"16", x"18", 
        x"29", x"41", x"44", x"40", x"4d", x"45", x"2b", x"27", x"35", x"3d", x"42", x"44", x"3e", x"3a", x"38", 
        x"39", x"2f", x"22", x"23", x"28", x"2f", x"2c", x"2a", x"38", x"55", x"61", x"66", x"65", x"69", x"6d", 
        x"71", x"74", x"71", x"70", x"66", x"64", x"6d", x"69", x"68", x"6a", x"6b", x"69", x"62", x"5e", x"63", 
        x"22", x"3d", x"45", x"45", x"74", x"65", x"45", x"2b", x"2a", x"48", x"40", x"30", x"2a", x"2c", x"23", 
        x"25", x"27", x"22", x"7d", x"d8", x"c3", x"cd", x"dd", x"c6", x"c2", x"d0", x"df", x"dc", x"e0", x"df", 
        x"e1", x"e2", x"e2", x"e1", x"e1", x"e3", x"e9", x"e7", x"e6", x"e6", x"e3", x"e2", x"e6", x"e4", x"e5", 
        x"ea", x"e3", x"e0", x"e2", x"e1", x"e2", x"e2", x"e1", x"e7", x"e7", x"e8", x"e6", x"e5", x"e6", x"e4", 
        x"e3", x"e6", x"e4", x"e6", x"e7", x"e7", x"e6", x"e8", x"e5", x"e2", x"e4", x"e6", x"e7", x"e7", x"df", 
        x"e0", x"e4", x"e2", x"e1", x"e0", x"e4", x"d3", x"ce", x"e6", x"de", x"e3", x"e6", x"e3", x"e6", x"ea", 
        x"e5", x"e4", x"e3", x"e1", x"de", x"e0", x"e4", x"e5", x"e6", x"e7", x"e8", x"e3", x"e4", x"e8", x"e6", 
        x"e3", x"e4", x"e5", x"e7", x"e9", x"e8", x"e8", x"e9", x"e9", x"eb", x"e5", x"e8", x"e6", x"e7", x"ec", 
        x"ec", x"ea", x"e5", x"e8", x"e8", x"e7", x"e9", x"e8", x"e7", x"ea", x"e6", x"e2", x"e8", x"eb", x"ea", 
        x"eb", x"e5", x"de", x"e6", x"ea", x"e8", x"ed", x"ee", x"ee", x"ee", x"de", x"d9", x"e3", x"e8", x"e7", 
        x"e7", x"e7", x"e9", x"e9", x"ef", x"e5", x"e4", x"ed", x"ea", x"ec", x"eb", x"e8", x"eb", x"e9", x"e9", 
        x"ea", x"ec", x"e9", x"ee", x"e8", x"e9", x"ed", x"ea", x"e8", x"ea", x"e9", x"ec", x"ec", x"e9", x"e9", 
        x"eb", x"ed", x"e5", x"e7", x"e7", x"e9", x"ed", x"ee", x"ed", x"eb", x"ea", x"ea", x"ec", x"ec", x"ec", 
        x"ec", x"ea", x"ea", x"ea", x"ec", x"ec", x"e7", x"e8", x"eb", x"ec", x"ea", x"ea", x"eb", x"ed", x"ec", 
        x"ed", x"ec", x"e9", x"e9", x"e4", x"e3", x"e8", x"e9", x"ea", x"ea", x"ec", x"ed", x"ec", x"eb", x"e9", 
        x"e8", x"e9", x"eb", x"ec", x"ea", x"eb", x"ec", x"e7", x"e3", x"e6", x"eb", x"e9", x"eb", x"ee", x"ed", 
        x"ed", x"ea", x"e9", x"e8", x"e9", x"ec", x"ee", x"ec", x"e9", x"e9", x"eb", x"eb", x"ee", x"ed", x"e8", 
        x"ec", x"ea", x"e8", x"ee", x"eb", x"ec", x"ec", x"ea", x"ed", x"ee", x"eb", x"eb", x"e8", x"eb", x"ed", 
        x"ed", x"ec", x"e7", x"ea", x"ed", x"ea", x"e9", x"e5", x"e7", x"ea", x"e6", x"e8", x"ed", x"ea", x"ea", 
        x"ea", x"ea", x"ea", x"e9", x"e9", x"eb", x"ed", x"ec", x"ec", x"ec", x"eb", x"ec", x"ed", x"ec", x"ec", 
        x"ec", x"ed", x"ee", x"e4", x"e5", x"ea", x"e9", x"ed", x"eb", x"ec", x"eb", x"e8", x"ea", x"e9", x"eb", 
        x"e9", x"e3", x"e7", x"e9", x"ea", x"f0", x"ed", x"eb", x"ea", x"e6", x"ea", x"ed", x"e9", x"eb", x"ed", 
        x"ec", x"e9", x"ea", x"eb", x"ec", x"ed", x"eb", x"ec", x"eb", x"ed", x"ee", x"ee", x"ed", x"ed", x"ed", 
        x"eb", x"ee", x"ec", x"ec", x"eb", x"ea", x"ed", x"f0", x"ed", x"ea", x"ef", x"f0", x"ed", x"f1", x"ef", 
        x"ed", x"ed", x"ed", x"eb", x"ed", x"ed", x"ec", x"ed", x"ed", x"ea", x"e9", x"eb", x"ed", x"ec", x"ea", 
        x"eb", x"ec", x"de", x"ea", x"ee", x"ee", x"ed", x"ef", x"f0", x"f1", x"f0", x"ee", x"ed", x"f1", x"f0", 
        x"ed", x"ee", x"ef", x"ed", x"ee", x"ef", x"f0", x"f0", x"ef", x"f0", x"f0", x"f2", x"f4", x"f5", x"f5", 
        x"f5", x"f4", x"f1", x"f0", x"ee", x"ed", x"ee", x"ee", x"f1", x"f2", x"f2", x"f1", x"ee", x"ee", x"f0", 
        x"f0", x"f1", x"f1", x"ef", x"ee", x"ed", x"ed", x"ee", x"ef", x"f0", x"f0", x"ef", x"ed", x"ee", x"ed", 
        x"ee", x"ef", x"ef", x"f0", x"f0", x"e5", x"eb", x"ed", x"ee", x"f0", x"f1", x"f1", x"f0", x"f1", x"f2", 
        x"f2", x"f1", x"f0", x"f2", x"f4", x"f3", x"f0", x"ee", x"f0", x"f3", x"f2", x"f0", x"f2", x"f4", x"f3", 
        x"f2", x"f1", x"ee", x"ef", x"f0", x"f2", x"f1", x"f0", x"ee", x"ed", x"ee", x"ec", x"ef", x"ef", x"f0", 
        x"f0", x"ef", x"ef", x"ef", x"ee", x"ed", x"ec", x"ec", x"ef", x"ef", x"ee", x"ec", x"ee", x"ea", x"e4", 
        x"e9", x"f0", x"e1", x"68", x"5f", x"91", x"8e", x"ad", x"af", x"e2", x"f2", x"f0", x"ed", x"ee", x"e6", 
        x"e8", x"ea", x"e3", x"d9", x"dc", x"d9", x"d0", x"d3", x"d6", x"a7", x"5b", x"5e", x"5a", x"60", x"60", 
        x"64", x"67", x"6c", x"71", x"6c", x"6e", x"76", x"7a", x"4c", x"15", x"0c", x"32", x"4f", x"1e", x"0c", 
        x"09", x"14", x"64", x"85", x"9c", x"ae", x"ba", x"b4", x"6d", x"71", x"6f", x"72", x"74", x"6a", x"6b", 
        x"59", x"1e", x"11", x"0b", x"40", x"7d", x"2f", x"0f", x"08", x"2d", x"7c", x"5b", x"46", x"4d", x"4d", 
        x"47", x"40", x"55", x"52", x"35", x"67", x"78", x"78", x"3e", x"4c", x"55", x"4f", x"6a", x"5d", x"2c", 
        x"20", x"19", x"1a", x"23", x"34", x"14", x"0d", x"0a", x"0c", x"32", x"58", x"60", x"56", x"54", x"5e", 
        x"2a", x"2d", x"3b", x"22", x"21", x"23", x"1f", x"1d", x"1c", x"1b", x"1c", x"25", x"25", x"1f", x"23", 
        x"1e", x"1e", x"27", x"3a", x"26", x"25", x"22", x"25", x"29", x"25", x"2f", x"5c", x"a9", x"b8", x"b9", 
        x"d2", x"b3", x"61", x"84", x"bd", x"c9", x"be", x"d1", x"ce", x"b2", x"af", x"b9", x"a5", x"79", x"77", 
        x"c5", x"aa", x"4c", x"40", x"42", x"40", x"40", x"43", x"48", x"57", x"52", x"4b", x"4b", x"47", x"4c", 
        x"50", x"57", x"53", x"50", x"51", x"4e", x"4d", x"4f", x"4e", x"53", x"55", x"4e", x"4c", x"4e", x"4c", 
        x"49", x"46", x"50", x"56", x"55", x"5b", x"5e", x"60", x"6b", x"6d", x"68", x"6d", x"65", x"59", x"4f", 
        x"4d", x"4d", x"4f", x"4e", x"51", x"61", x"59", x"4e", x"4f", x"55", x"56", x"52", x"50", x"4d", x"46", 
        x"41", x"46", x"47", x"3c", x"3a", x"3a", x"3b", x"3a", x"34", x"2d", x"2a", x"2a", x"24", x"1d", x"22", 
        x"42", x"58", x"4d", x"6d", x"9f", x"6b", x"44", x"2f", x"40", x"51", x"46", x"3d", x"28", x"23", x"28", 
        x"37", x"34", x"25", x"7a", x"dc", x"c7", x"c6", x"d8", x"ca", x"c8", x"d3", x"e1", x"df", x"e4", x"e0", 
        x"e3", x"e3", x"de", x"df", x"e1", x"e6", x"e9", x"e8", x"eb", x"e7", x"e0", x"e1", x"e2", x"de", x"dd", 
        x"e3", x"e5", x"e2", x"dc", x"de", x"e5", x"e5", x"e1", x"e5", x"e4", x"e4", x"e2", x"e4", x"e6", x"e3", 
        x"e4", x"e2", x"e4", x"ea", x"e5", x"e3", x"e5", x"e2", x"e2", x"e0", x"dc", x"e2", x"e5", x"e7", x"e5", 
        x"e7", x"e8", x"e1", x"df", x"db", x"dd", x"cb", x"c8", x"e7", x"e8", x"e9", x"ec", x"e4", x"e2", x"e5", 
        x"e6", x"e5", x"e0", x"e0", x"e3", x"e6", x"e4", x"e1", x"e5", x"e8", x"e8", x"e2", x"e0", x"e1", x"df", 
        x"e4", x"e6", x"e3", x"e4", x"e7", x"e7", x"e8", x"e7", x"e6", x"e9", x"e6", x"e9", x"e7", x"e8", x"ec", 
        x"eb", x"e9", x"ea", x"ea", x"e8", x"e7", x"ea", x"ea", x"e6", x"eb", x"e7", x"e1", x"e4", x"e7", x"e6", 
        x"e6", x"eb", x"ea", x"eb", x"ed", x"e9", x"eb", x"ec", x"e8", x"e4", x"e1", x"e1", x"e9", x"eb", x"e7", 
        x"e8", x"e6", x"e8", x"e9", x"ef", x"e7", x"e5", x"eb", x"ea", x"ec", x"ec", x"ea", x"eb", x"ea", x"ea", 
        x"e6", x"eb", x"e8", x"eb", x"e9", x"e9", x"ec", x"e9", x"e5", x"e8", x"e9", x"ec", x"eb", x"e8", x"e9", 
        x"ee", x"ea", x"e5", x"ee", x"ee", x"e9", x"ec", x"ef", x"ed", x"ea", x"e8", x"e8", x"ea", x"ec", x"ef", 
        x"ed", x"e8", x"e5", x"e7", x"ec", x"ee", x"ea", x"ea", x"eb", x"e9", x"e7", x"e9", x"ec", x"ee", x"ef", 
        x"ee", x"ea", x"ea", x"eb", x"e0", x"e3", x"eb", x"e9", x"e9", x"e9", x"eb", x"eb", x"ea", x"e8", x"e7", 
        x"e9", x"ed", x"eb", x"ea", x"ec", x"ec", x"ec", x"e7", x"e4", x"e6", x"e8", x"e9", x"eb", x"ee", x"ee", 
        x"ed", x"e8", x"e7", x"e7", x"ec", x"ed", x"ec", x"e8", x"e4", x"e5", x"e9", x"ea", x"ec", x"ed", x"ea", 
        x"ea", x"e8", x"ea", x"ee", x"ed", x"ee", x"eb", x"e6", x"eb", x"ee", x"ea", x"ea", x"ea", x"ed", x"eb", 
        x"eb", x"ec", x"e2", x"e7", x"ea", x"e8", x"e9", x"e8", x"eb", x"ec", x"e8", x"ea", x"f0", x"ed", x"eb", 
        x"ec", x"e9", x"e9", x"e7", x"e7", x"ec", x"ee", x"eb", x"ee", x"ee", x"ec", x"eb", x"eb", x"ec", x"ee", 
        x"ed", x"ec", x"ee", x"e3", x"e4", x"eb", x"ea", x"ed", x"ea", x"ed", x"ed", x"ea", x"ea", x"ea", x"ec", 
        x"ea", x"e6", x"e8", x"e9", x"e9", x"ed", x"eb", x"ea", x"ee", x"eb", x"ea", x"ec", x"e7", x"e8", x"eb", 
        x"ec", x"e9", x"eb", x"ea", x"eb", x"ec", x"ec", x"ed", x"eb", x"ee", x"eb", x"ea", x"ed", x"ee", x"eb", 
        x"e9", x"eb", x"e7", x"e9", x"eb", x"eb", x"ef", x"f0", x"ee", x"ef", x"f0", x"ec", x"ea", x"f0", x"f1", 
        x"ee", x"ef", x"ed", x"e7", x"ea", x"ed", x"ec", x"ed", x"ed", x"e8", x"e6", x"e8", x"eb", x"ec", x"ec", 
        x"ec", x"ed", x"e0", x"ea", x"ef", x"ee", x"ee", x"ef", x"f1", x"f1", x"f0", x"ed", x"ed", x"f2", x"f2", 
        x"ef", x"ef", x"f1", x"ef", x"f0", x"f0", x"f2", x"f3", x"f2", x"ef", x"ef", x"f2", x"f4", x"f5", x"f6", 
        x"f5", x"f4", x"f2", x"f1", x"f0", x"ed", x"ee", x"f0", x"f2", x"f1", x"f0", x"f0", x"ed", x"ed", x"f1", 
        x"f0", x"f2", x"f3", x"f0", x"f0", x"ed", x"ec", x"ef", x"f1", x"f1", x"ee", x"f0", x"ee", x"ee", x"ec", 
        x"ee", x"ec", x"ee", x"ed", x"ed", x"e4", x"ec", x"ef", x"f0", x"f2", x"f0", x"ee", x"ee", x"f0", x"f2", 
        x"f2", x"f1", x"f0", x"f3", x"f5", x"f5", x"f2", x"f0", x"f0", x"f2", x"f2", x"f0", x"f2", x"f3", x"f2", 
        x"f0", x"f1", x"f0", x"f0", x"f1", x"f0", x"ef", x"ef", x"ef", x"eb", x"ed", x"ec", x"ec", x"ea", x"eb", 
        x"ec", x"ed", x"ef", x"ef", x"ef", x"ef", x"ec", x"ea", x"ed", x"ee", x"ed", x"ef", x"f0", x"ed", x"e8", 
        x"ea", x"ed", x"c7", x"60", x"67", x"90", x"82", x"94", x"b6", x"e6", x"f3", x"f0", x"ed", x"d8", x"ad", 
        x"a2", x"a3", x"9a", x"84", x"84", x"7e", x"7b", x"79", x"76", x"7d", x"7a", x"75", x"6f", x"6e", x"69", 
        x"6a", x"68", x"66", x"63", x"5f", x"5f", x"5f", x"5e", x"3b", x"16", x"09", x"06", x"09", x"0b", x"0a", 
        x"09", x"07", x"30", x"48", x"82", x"b4", x"ac", x"8a", x"23", x"27", x"26", x"29", x"2b", x"26", x"1b", 
        x"1c", x"15", x"0d", x"0a", x"10", x"1b", x"0c", x"0f", x"0a", x"33", x"7e", x"3e", x"14", x"25", x"29", 
        x"26", x"21", x"47", x"55", x"3a", x"63", x"75", x"78", x"3e", x"44", x"50", x"49", x"68", x"67", x"3c", 
        x"2f", x"20", x"24", x"21", x"20", x"1c", x"2d", x"36", x"38", x"4c", x"58", x"70", x"6d", x"64", x"6b", 
        x"58", x"64", x"62", x"4b", x"50", x"52", x"3e", x"3c", x"40", x"3f", x"49", x"53", x"58", x"54", x"5c", 
        x"62", x"60", x"67", x"70", x"5d", x"59", x"5c", x"65", x"6b", x"71", x"74", x"6a", x"80", x"b9", x"b6", 
        x"cb", x"b8", x"93", x"a2", x"ae", x"d6", x"b4", x"b8", x"cc", x"cb", x"c1", x"bd", x"ac", x"80", x"73", 
        x"ba", x"bc", x"86", x"86", x"84", x"83", x"84", x"7b", x"74", x"75", x"76", x"77", x"79", x"6f", x"6e", 
        x"6f", x"6f", x"6c", x"66", x"5e", x"57", x"54", x"4a", x"4a", x"49", x"53", x"59", x"55", x"4f", x"45", 
        x"48", x"46", x"42", x"43", x"3f", x"3d", x"3a", x"3a", x"47", x"43", x"36", x"36", x"32", x"2e", x"2a", 
        x"28", x"28", x"2a", x"21", x"26", x"47", x"2c", x"20", x"1f", x"19", x"17", x"14", x"16", x"0b", x"09", 
        x"0b", x"0e", x"0f", x"0a", x"24", x"21", x"09", x"06", x"04", x"02", x"03", x"04", x"04", x"02", x"02", 
        x"5e", x"4c", x"33", x"89", x"c0", x"75", x"25", x"20", x"2a", x"30", x"36", x"36", x"35", x"29", x"21", 
        x"29", x"30", x"31", x"8b", x"e4", x"cb", x"cb", x"dd", x"ca", x"c3", x"cc", x"dc", x"e1", x"e6", x"e1", 
        x"e1", x"e1", x"e1", x"e7", x"e3", x"df", x"dc", x"e4", x"e3", x"df", x"dd", x"e5", x"ea", x"e4", x"e0", 
        x"e9", x"e9", x"e3", x"e1", x"e2", x"e6", x"e5", x"e1", x"e3", x"e1", x"e2", x"e1", x"e3", x"e4", x"e5", 
        x"ea", x"e7", x"e4", x"e3", x"e1", x"e1", x"e6", x"e4", x"e4", x"e6", x"e2", x"e3", x"e3", x"e0", x"df", 
        x"e2", x"e6", x"e7", x"e5", x"e4", x"e7", x"e3", x"e2", x"e8", x"ea", x"ea", x"e7", x"e2", x"e3", x"e7", 
        x"e9", x"e8", x"e2", x"de", x"e2", x"e8", x"e7", x"e1", x"e5", x"e7", x"e6", x"e0", x"e4", x"df", x"d9", 
        x"e0", x"e3", x"e2", x"e4", x"e4", x"e5", x"ea", x"ec", x"ea", x"ec", x"ec", x"eb", x"e9", x"ea", x"ec", 
        x"eb", x"eb", x"ed", x"e8", x"e9", x"ea", x"e9", x"ec", x"ea", x"eb", x"e8", x"e5", x"e6", x"e7", x"e5", 
        x"e3", x"e6", x"e7", x"e8", x"e9", x"ec", x"ec", x"ea", x"e7", x"e2", x"e8", x"ea", x"eb", x"e8", x"e3", 
        x"ea", x"e8", x"e6", x"e9", x"ec", x"ea", x"e9", x"e9", x"e8", x"e9", x"ea", x"e9", x"e8", x"e7", x"e8", 
        x"e7", x"ec", x"ec", x"e9", x"e8", x"ea", x"ec", x"eb", x"eb", x"ec", x"eb", x"ed", x"eb", x"e8", x"ea", 
        x"ec", x"e7", x"ea", x"e9", x"e4", x"e8", x"eb", x"e7", x"e7", x"e7", x"e8", x"e8", x"e8", x"e9", x"eb", 
        x"eb", x"eb", x"ea", x"e9", x"eb", x"ec", x"eb", x"eb", x"e9", x"e5", x"e3", x"e6", x"e9", x"e5", x"e9", 
        x"ec", x"eb", x"ed", x"ea", x"de", x"e1", x"eb", x"e9", x"e6", x"e6", x"e7", x"e8", x"e8", x"e9", x"eb", 
        x"ec", x"ee", x"ea", x"e7", x"eb", x"eb", x"eb", x"e9", x"e9", x"e9", x"e8", x"ea", x"e9", x"eb", x"eb", 
        x"eb", x"e7", x"e7", x"e8", x"ea", x"eb", x"ec", x"eb", x"e8", x"e7", x"e7", x"eb", x"e9", x"ee", x"f1", 
        x"ea", x"e8", x"e8", x"e9", x"eb", x"ee", x"eb", x"e8", x"eb", x"ee", x"ee", x"ef", x"ee", x"ed", x"ef", 
        x"e9", x"e9", x"eb", x"eb", x"ed", x"eb", x"ed", x"ed", x"ee", x"ea", x"e7", x"e8", x"ee", x"ec", x"ec", 
        x"f0", x"ee", x"ea", x"e7", x"e8", x"ed", x"ed", x"ea", x"eb", x"ec", x"ea", x"ec", x"ea", x"eb", x"ed", 
        x"ec", x"eb", x"ee", x"e2", x"e2", x"ed", x"ec", x"ed", x"e8", x"ec", x"ed", x"ea", x"ea", x"e9", x"ec", 
        x"ea", x"ec", x"ea", x"eb", x"ea", x"eb", x"eb", x"ec", x"ef", x"ee", x"eb", x"ec", x"ea", x"eb", x"ec", 
        x"ef", x"eb", x"ee", x"eb", x"e8", x"e8", x"e9", x"ec", x"eb", x"ee", x"eb", x"ea", x"ee", x"f1", x"ef", 
        x"ee", x"ee", x"e9", x"eb", x"ee", x"eb", x"ee", x"ec", x"eb", x"ee", x"ef", x"eb", x"ea", x"ef", x"f0", 
        x"e8", x"ee", x"f1", x"eb", x"ea", x"ea", x"ec", x"ef", x"ee", x"eb", x"ea", x"eb", x"ea", x"eb", x"ee", 
        x"ed", x"ed", x"e2", x"ea", x"ee", x"f0", x"ef", x"ee", x"ee", x"ef", x"ef", x"ef", x"ef", x"ef", x"ee", 
        x"ec", x"eb", x"ef", x"ec", x"ee", x"ef", x"ef", x"ef", x"f0", x"f0", x"f0", x"f4", x"f5", x"f5", x"f5", 
        x"f6", x"f4", x"f2", x"f0", x"f1", x"f0", x"f0", x"f1", x"f2", x"ef", x"ee", x"f0", x"ee", x"ed", x"f1", 
        x"ef", x"f0", x"f2", x"ed", x"ef", x"ee", x"ee", x"f0", x"f1", x"f0", x"ee", x"f0", x"f0", x"ef", x"ef", 
        x"ef", x"ea", x"ec", x"ee", x"ed", x"e4", x"ef", x"ef", x"ed", x"ee", x"ee", x"ef", x"f0", x"f0", x"f1", 
        x"f1", x"f1", x"f2", x"f5", x"f7", x"f5", x"f3", x"f3", x"f2", x"f2", x"f2", x"f1", x"f3", x"f3", x"f2", 
        x"ef", x"f1", x"f1", x"f2", x"f3", x"f1", x"ee", x"ee", x"ef", x"ee", x"f0", x"ee", x"ef", x"ed", x"ed", 
        x"ec", x"ec", x"ed", x"ec", x"ed", x"f0", x"ee", x"ec", x"ed", x"ea", x"eb", x"eb", x"ea", x"e7", x"e3", 
        x"e5", x"ec", x"a0", x"67", x"94", x"9e", x"66", x"9c", x"df", x"ef", x"ef", x"ef", x"cc", x"77", x"4a", 
        x"42", x"3f", x"3f", x"40", x"3e", x"30", x"2e", x"30", x"39", x"41", x"2e", x"2f", x"30", x"37", x"36", 
        x"33", x"2e", x"2d", x"2c", x"37", x"3b", x"33", x"26", x"1b", x"0b", x"05", x"09", x"08", x"09", x"09", 
        x"1c", x"2e", x"37", x"49", x"84", x"bc", x"bf", x"86", x"24", x"36", x"2b", x"1d", x"1b", x"22", x"27", 
        x"1f", x"19", x"08", x"0a", x"09", x"08", x"07", x"07", x"07", x"27", x"61", x"54", x"3d", x"44", x"3d", 
        x"35", x"34", x"4f", x"54", x"3b", x"59", x"76", x"79", x"52", x"56", x"61", x"5f", x"79", x"79", x"66", 
        x"69", x"63", x"68", x"66", x"57", x"31", x"4a", x"5c", x"64", x"67", x"53", x"5c", x"62", x"62", x"75", 
        x"8f", x"8b", x"81", x"84", x"80", x"79", x"76", x"7b", x"7d", x"7a", x"76", x"73", x"77", x"6e", x"66", 
        x"69", x"64", x"66", x"61", x"60", x"5c", x"57", x"58", x"5c", x"5f", x"5b", x"80", x"71", x"97", x"c3", 
        x"c9", x"b9", x"9d", x"af", x"a8", x"d8", x"c8", x"b5", x"b5", x"b4", x"c4", x"bd", x"b3", x"99", x"7f", 
        x"bb", x"9d", x"3e", x"33", x"31", x"31", x"2f", x"2c", x"36", x"2f", x"25", x"27", x"2b", x"23", x"1f", 
        x"1f", x"1e", x"1b", x"31", x"4a", x"1f", x"0d", x"13", x"13", x"13", x"13", x"1a", x"19", x"12", x"11", 
        x"1d", x"22", x"0e", x"0c", x"0b", x"0c", x"09", x"10", x"1f", x"12", x"07", x"07", x"09", x"07", x"05", 
        x"04", x"04", x"06", x"05", x"13", x"41", x"16", x"0b", x"0b", x"0a", x"09", x"0a", x"13", x"0a", x"09", 
        x"0d", x"0c", x"0b", x"08", x"30", x"37", x"14", x"11", x"14", x"15", x"17", x"11", x"11", x"20", x"20", 
        x"5e", x"49", x"2c", x"91", x"d0", x"76", x"17", x"15", x"25", x"28", x"34", x"30", x"2c", x"30", x"33", 
        x"2e", x"28", x"25", x"86", x"e1", x"c7", x"cd", x"db", x"c9", x"c6", x"cc", x"df", x"e3", x"e2", x"e1", 
        x"e3", x"e4", x"e0", x"e5", x"e3", x"e3", x"df", x"e2", x"d7", x"db", x"e2", x"e2", x"de", x"e2", x"e2", 
        x"e9", x"e7", x"e4", x"e7", x"e6", x"e3", x"e2", x"e0", x"e2", x"e1", x"e3", x"e3", x"e5", x"e7", x"e4", 
        x"e8", x"e7", x"e1", x"df", x"e7", x"e3", x"e4", x"e7", x"e4", x"e4", x"e1", x"e1", x"e3", x"e3", x"e5", 
        x"e4", x"e5", x"e7", x"e4", x"e8", x"e5", x"e5", x"eb", x"e8", x"e4", x"e6", x"e5", x"e4", x"e5", x"e5", 
        x"e3", x"e6", x"e7", x"e5", x"e7", x"e8", x"e9", x"e6", x"ea", x"e9", x"e8", x"e3", x"e4", x"e2", x"e1", 
        x"e5", x"e4", x"e5", x"e5", x"e2", x"e3", x"e8", x"ea", x"e8", x"ea", x"ef", x"ec", x"e8", x"e8", x"ea", 
        x"e9", x"eb", x"ea", x"e5", x"ea", x"ea", x"e3", x"e5", x"e4", x"e8", x"e9", x"e6", x"e5", x"e5", x"e7", 
        x"e9", x"ea", x"e9", x"e9", x"e7", x"e8", x"e9", x"e9", x"e9", x"e9", x"ec", x"e9", x"e8", x"e5", x"e0", 
        x"e8", x"e7", x"e7", x"eb", x"e8", x"e9", x"eb", x"eb", x"eb", x"eb", x"ec", x"eb", x"e8", x"e8", x"ea", 
        x"ed", x"eb", x"ec", x"e9", x"e8", x"ec", x"ee", x"ea", x"e9", x"ea", x"ea", x"ec", x"ec", x"ea", x"ea", 
        x"ec", x"ed", x"ef", x"ea", x"e4", x"e9", x"ec", x"e9", x"ea", x"eb", x"ec", x"ec", x"eb", x"ea", x"eb", 
        x"ea", x"ec", x"ed", x"ea", x"e9", x"ed", x"ec", x"ec", x"eb", x"e9", x"e8", x"ea", x"ec", x"e7", x"eb", 
        x"ee", x"eb", x"ed", x"eb", x"e5", x"e3", x"e5", x"e7", x"e8", x"e6", x"e8", x"ed", x"ec", x"ea", x"ec", 
        x"ea", x"ed", x"ee", x"ea", x"e9", x"ec", x"ea", x"e7", x"e8", x"e7", x"e6", x"ea", x"e8", x"eb", x"eb", 
        x"ec", x"e9", x"ea", x"ec", x"e8", x"e9", x"ed", x"ec", x"e9", x"e9", x"ec", x"eb", x"e6", x"eb", x"f0", 
        x"ee", x"eb", x"e8", x"ea", x"ed", x"f0", x"ed", x"eb", x"e9", x"ea", x"ec", x"ed", x"e8", x"de", x"e9", 
        x"ec", x"e8", x"ea", x"e8", x"ed", x"ee", x"ef", x"ed", x"ed", x"ea", x"ea", x"e6", x"eb", x"ec", x"ec", 
        x"ee", x"f0", x"ea", x"e8", x"e9", x"ec", x"ec", x"eb", x"eb", x"e9", x"ea", x"ed", x"ec", x"eb", x"ec", 
        x"ec", x"eb", x"ec", x"e3", x"e4", x"ec", x"eb", x"ed", x"e9", x"eb", x"ed", x"eb", x"e9", x"ea", x"ec", 
        x"eb", x"ea", x"e7", x"eb", x"eb", x"eb", x"ec", x"ec", x"ec", x"ed", x"e9", x"eb", x"ec", x"ec", x"eb", 
        x"ec", x"e9", x"ee", x"eb", x"e8", x"e9", x"ea", x"ef", x"ee", x"ee", x"ed", x"eb", x"eb", x"eb", x"ec", 
        x"ee", x"ee", x"e8", x"ec", x"ef", x"ea", x"ec", x"eb", x"ea", x"ed", x"ef", x"ec", x"ec", x"ee", x"ee", 
        x"e1", x"e9", x"ee", x"ed", x"ed", x"ec", x"ec", x"eb", x"ea", x"eb", x"ee", x"ee", x"e8", x"e9", x"f0", 
        x"ed", x"ed", x"e4", x"e9", x"ed", x"f0", x"ed", x"ee", x"ee", x"ef", x"f0", x"f0", x"ef", x"ee", x"ec", 
        x"eb", x"ea", x"ee", x"ec", x"ef", x"f3", x"ef", x"ed", x"ee", x"f1", x"f1", x"f3", x"f6", x"f7", x"f7", 
        x"f6", x"f4", x"f1", x"ef", x"f1", x"f1", x"ef", x"f1", x"f2", x"f0", x"f0", x"f2", x"ee", x"ed", x"f1", 
        x"ed", x"ed", x"ef", x"eb", x"ee", x"f0", x"f1", x"f1", x"ef", x"ee", x"ed", x"ee", x"ee", x"ef", x"f1", 
        x"f2", x"ea", x"ed", x"ef", x"ed", x"e3", x"ed", x"ee", x"eb", x"ef", x"ef", x"ef", x"f1", x"f1", x"f1", 
        x"f2", x"f3", x"f4", x"f5", x"f5", x"f2", x"f1", x"f2", x"f1", x"f2", x"f3", x"f2", x"f4", x"f3", x"f2", 
        x"ef", x"f1", x"ef", x"f2", x"f3", x"f1", x"ef", x"f0", x"f1", x"ef", x"ed", x"eb", x"ee", x"f1", x"f0", 
        x"ee", x"ee", x"ef", x"ec", x"eb", x"f0", x"ee", x"ec", x"ed", x"ea", x"ea", x"eb", x"e7", x"e5", x"e3", 
        x"eb", x"d6", x"78", x"6e", x"80", x"9a", x"9e", x"bf", x"ec", x"ef", x"e7", x"eb", x"bc", x"48", x"33", 
        x"2c", x"2e", x"3a", x"4f", x"43", x"2d", x"2f", x"2d", x"3b", x"49", x"23", x"28", x"2c", x"31", x"31", 
        x"32", x"36", x"40", x"39", x"3e", x"46", x"45", x"43", x"45", x"46", x"42", x"4b", x"4b", x"46", x"38", 
        x"6a", x"9b", x"74", x"64", x"98", x"ba", x"bb", x"a3", x"5e", x"6b", x"64", x"65", x"61", x"67", x"74", 
        x"75", x"53", x"30", x"1b", x"09", x"0a", x"0a", x"07", x"0f", x"35", x"55", x"71", x"7a", x"7a", x"70", 
        x"69", x"6a", x"64", x"49", x"37", x"54", x"7c", x"7e", x"6e", x"75", x"7d", x"77", x"7f", x"81", x"6a", 
        x"67", x"64", x"68", x"69", x"51", x"2a", x"43", x"5a", x"5c", x"57", x"4f", x"57", x"4b", x"5f", x"79", 
        x"63", x"46", x"45", x"45", x"41", x"36", x"43", x"47", x"3c", x"41", x"40", x"33", x"33", x"36", x"22", 
        x"1f", x"1d", x"1a", x"1c", x"30", x"2b", x"19", x"17", x"19", x"1b", x"35", x"74", x"89", x"72", x"bb", 
        x"d4", x"a5", x"a2", x"bc", x"bb", x"cf", x"d4", x"ba", x"bf", x"b2", x"b2", x"b9", x"ab", x"8a", x"7a", 
        x"b9", x"86", x"18", x"11", x"10", x"0e", x"0c", x"17", x"39", x"30", x"0d", x"0e", x"0f", x"0e", x"12", 
        x"11", x"0c", x"09", x"25", x"48", x"1e", x"0a", x"0d", x"0f", x"11", x"11", x"14", x"14", x"14", x"13", 
        x"2e", x"3a", x"13", x"0f", x"0f", x"11", x"14", x"21", x"32", x"2d", x"35", x"3e", x"3e", x"2f", x"1f", 
        x"13", x"14", x"14", x"12", x"1f", x"56", x"41", x"35", x"3b", x"33", x"24", x"26", x"35", x"2c", x"37", 
        x"3a", x"2f", x"33", x"39", x"55", x"5a", x"40", x"44", x"47", x"42", x"45", x"3c", x"39", x"4d", x"4c", 
        x"6b", x"6d", x"58", x"83", x"d0", x"8f", x"26", x"25", x"27", x"2a", x"24", x"1d", x"19", x"20", x"3a", 
        x"33", x"33", x"26", x"80", x"da", x"c5", x"ca", x"d9", x"c4", x"bf", x"cd", x"d9", x"e0", x"e5", x"e1", 
        x"e1", x"e2", x"e0", x"e5", x"e5", x"df", x"df", x"df", x"da", x"dd", x"e3", x"e2", x"dc", x"e5", x"e7", 
        x"e4", x"e6", x"e9", x"e7", x"e5", x"db", x"df", x"e8", x"e7", x"e4", x"e4", x"e6", x"e8", x"e4", x"e5", 
        x"e7", x"e1", x"e3", x"e7", x"e3", x"df", x"e7", x"e4", x"e3", x"e6", x"d9", x"d9", x"e2", x"e8", x"e8", 
        x"e5", x"e4", x"e4", x"e7", x"e6", x"e3", x"e7", x"ea", x"e8", x"e3", x"e6", x"e8", x"e8", x"e5", x"e9", 
        x"e4", x"e3", x"e3", x"e4", x"e8", x"e7", x"e6", x"ea", x"eb", x"e8", x"e7", x"e3", x"df", x"e1", x"e4", 
        x"e7", x"e4", x"e7", x"e5", x"e4", x"e3", x"e6", x"ea", x"e7", x"ea", x"ec", x"eb", x"e8", x"e3", x"ea", 
        x"eb", x"eb", x"e5", x"e5", x"eb", x"e8", x"e7", x"e7", x"e5", x"ea", x"ed", x"e7", x"ec", x"eb", x"ea", 
        x"e9", x"eb", x"e7", x"e3", x"e7", x"e7", x"e6", x"ea", x"eb", x"e6", x"e9", x"e9", x"eb", x"ec", x"e9", 
        x"e9", x"e7", x"ea", x"eb", x"e7", x"e7", x"eb", x"ea", x"ea", x"e6", x"e8", x"ec", x"ea", x"ec", x"ed", 
        x"eb", x"ed", x"f1", x"f0", x"e6", x"e9", x"ef", x"ed", x"e6", x"e7", x"eb", x"ea", x"eb", x"ea", x"e9", 
        x"e8", x"ea", x"eb", x"eb", x"eb", x"ee", x"ef", x"ee", x"ed", x"ed", x"ef", x"ea", x"eb", x"ea", x"e8", 
        x"e9", x"eb", x"eb", x"e8", x"e8", x"ea", x"f0", x"ec", x"e8", x"ea", x"eb", x"e9", x"ea", x"eb", x"ec", 
        x"ef", x"eb", x"e9", x"ec", x"e8", x"e5", x"e7", x"eb", x"ed", x"eb", x"e9", x"eb", x"eb", x"eb", x"ec", 
        x"e7", x"eb", x"ed", x"ed", x"ec", x"ec", x"ed", x"ea", x"e6", x"e5", x"e5", x"e6", x"e9", x"ed", x"eb", 
        x"ec", x"ed", x"e7", x"eb", x"ec", x"e9", x"ee", x"ec", x"eb", x"ee", x"ed", x"ea", x"e9", x"eb", x"eb", 
        x"ec", x"eb", x"eb", x"ed", x"eb", x"ea", x"ec", x"eb", x"eb", x"ef", x"ee", x"e9", x"e7", x"e4", x"e6", 
        x"eb", x"ed", x"e8", x"e9", x"ec", x"ef", x"f0", x"ed", x"ea", x"ea", x"ea", x"ec", x"ee", x"ec", x"eb", 
        x"ea", x"ef", x"e8", x"ea", x"e8", x"e6", x"ec", x"eb", x"e9", x"eb", x"eb", x"e9", x"ea", x"ee", x"ee", 
        x"ec", x"ea", x"ed", x"e4", x"e2", x"e9", x"eb", x"ec", x"eb", x"ec", x"ec", x"ea", x"e8", x"e7", x"e9", 
        x"ea", x"e8", x"e8", x"eb", x"ec", x"ec", x"ea", x"e9", x"eb", x"ec", x"ea", x"ea", x"ea", x"eb", x"ec", 
        x"eb", x"eb", x"ef", x"ee", x"ea", x"e8", x"e9", x"ef", x"f1", x"ec", x"ea", x"ec", x"ef", x"e9", x"ea", 
        x"ef", x"ed", x"ea", x"eb", x"ec", x"eb", x"ef", x"ee", x"ee", x"ee", x"ed", x"ed", x"ee", x"ed", x"e9", 
        x"e5", x"e9", x"ef", x"ef", x"ed", x"ed", x"ef", x"ed", x"eb", x"ec", x"ee", x"ef", x"ec", x"eb", x"ed", 
        x"ee", x"ed", x"e0", x"e8", x"ee", x"ee", x"ee", x"ef", x"ed", x"ed", x"ed", x"ee", x"ec", x"ef", x"ee", 
        x"ed", x"ef", x"f0", x"ed", x"ec", x"f0", x"ef", x"ef", x"f0", x"f1", x"f2", x"f4", x"f6", x"f6", x"f6", 
        x"f7", x"f4", x"f0", x"f0", x"f0", x"f2", x"f0", x"ef", x"f3", x"f1", x"f0", x"f2", x"f3", x"f2", x"f2", 
        x"f3", x"f1", x"ee", x"ee", x"ef", x"ee", x"ed", x"ed", x"ef", x"ef", x"ee", x"f0", x"ef", x"ee", x"f1", 
        x"f0", x"eb", x"f1", x"ee", x"ed", x"e5", x"eb", x"ef", x"ec", x"ef", x"f2", x"f3", x"f3", x"f1", x"ef", 
        x"f0", x"ef", x"f0", x"f4", x"f5", x"f2", x"f1", x"f1", x"f1", x"f3", x"f2", x"ed", x"ef", x"ee", x"ee", 
        x"ef", x"f0", x"f1", x"f4", x"e6", x"e6", x"f1", x"f1", x"f0", x"ef", x"ef", x"ee", x"ee", x"ed", x"ec", 
        x"ec", x"ee", x"ef", x"ec", x"ea", x"eb", x"ef", x"f0", x"ed", x"eb", x"ec", x"ec", x"eb", x"e6", x"e1", 
        x"e6", x"ab", x"74", x"8a", x"76", x"5f", x"a4", x"7b", x"b7", x"ee", x"ea", x"e6", x"c2", x"6e", x"73", 
        x"70", x"71", x"76", x"88", x"84", x"75", x"6e", x"68", x"6b", x"77", x"75", x"75", x"70", x"71", x"77", 
        x"80", x"8b", x"96", x"91", x"8e", x"93", x"96", x"9a", x"98", x"9c", x"9b", x"9c", x"9d", x"8a", x"6e", 
        x"a0", x"c9", x"ab", x"7a", x"ac", x"b2", x"8e", x"99", x"76", x"7a", x"7c", x"7e", x"7d", x"77", x"6f", 
        x"6f", x"69", x"5e", x"33", x"1d", x"38", x"3e", x"1d", x"14", x"44", x"5b", x"57", x"43", x"46", x"47", 
        x"46", x"4c", x"3d", x"31", x"37", x"50", x"75", x"73", x"55", x"5a", x"74", x"79", x"84", x"8b", x"42", 
        x"27", x"3c", x"24", x"26", x"25", x"2d", x"43", x"59", x"68", x"61", x"3c", x"27", x"33", x"65", x"82", 
        x"38", x"0e", x"13", x"14", x"15", x"12", x"28", x"27", x"0c", x"0e", x"0e", x"0b", x"10", x"29", x"0f", 
        x"0b", x"0d", x"0b", x"12", x"27", x"20", x"0e", x"12", x"14", x"16", x"44", x"59", x"91", x"84", x"81", 
        x"cf", x"9a", x"8a", x"b6", x"bf", x"cb", x"da", x"c8", x"b8", x"c9", x"b2", x"b6", x"b9", x"8d", x"8d", 
        x"c3", x"7b", x"20", x"1a", x"1c", x"20", x"24", x"2a", x"4c", x"55", x"2e", x"25", x"22", x"32", x"37", 
        x"3b", x"44", x"40", x"3f", x"40", x"2b", x"1c", x"21", x"2d", x"3c", x"3d", x"3f", x"3e", x"46", x"46", 
        x"52", x"5c", x"4f", x"4a", x"49", x"51", x"4f", x"50", x"56", x"54", x"57", x"5b", x"5d", x"55", x"4b", 
        x"48", x"4b", x"50", x"58", x"58", x"66", x"65", x"69", x"6d", x"74", x"70", x"6d", x"6d", x"64", x"6c", 
        x"6d", x"60", x"62", x"67", x"64", x"62", x"62", x"64", x"62", x"5a", x"62", x"65", x"61", x"60", x"61"
    );
begin
    -- Port A
    process(i_clk_a)
    begin
        if(rising_edge(i_clk_a)) then 
            if(i_we_a = '1') then
                ram(i_addr_a) := i_data_a;
            end if;
            o_q_a <= ram(i_addr_a);
        end if;
    end process;
    
    -- Port B
    process(i_clk_b)
    begin
        if(rising_edge(i_clk_b)) then
            if(i_we_b = '1') then
                ram(i_addr_b) := i_data_b;
            end if;
            o_q_b <= ram(i_addr_b);
        end if;
    end process;
end rtl;
