��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_A?N��Y�jo���e�YI��#~B�t��@E����2u�@��G^��8�=�Q�Ps�t�N����ꈱX^�1��Fȑt��X���ސ�t\J���6����9*���$�L[P��#L�pfR������N�Gm�IGlr�FUx��盆(0�ܥ�!٨Im]�>��r�J������<{��	,�Y x{��a���T���9P7	����p��(p>��7YN����aD��Z�<�ѭu�W�B#�X�fn�ٿ��f����x�ڦ9B��B߳&B�24��f�����˹'qF�R��nE'��r=	���Tf0��6,p���g&O>Z���^y0�S.��RF����v�����CG<����G}J����y�'b���Q�;�K����ɘ>��سP�̫�Tہ����`J�� ]u�"��Mҧ��Mx�(�Hw�g��qV��8E!/=Н�-�9�E"M�3�n�o�b���� �P�Lc�! n���v�c�>��n�a}���D���(��G���'D�i����}�U��3��;K������Q�&�3����aLxmEQT義46��W������N`�hl���\ �ew!�L1���a���g�]��)<�cG��Ħaý��)�t2��a��_��t�D.���Q6�����̕&H#F�^�(��:��i*F�Y�n�����?������c�E�	Կ\�cb��z:��W,L8����o~��@�F��r�iAds�U	��̺���<�ʹ�m3V3=TH��n��@W	��#���B-�8C�S��nU�H���|����=�,t7s�c�f�4#U�^ :�)�C�+�2�(��a,��:Q�� ����_2�����c�2�U��zMjhHGd@f"jV��:��� �l�Rb���K�#�ƽ���"�}q�D	� ��=D���K�ߊ��3�j�����Z���:�I/s���e@i 5�0��}���Or�Z*���u待%��ia|?E�9?7���v����ƺ�A=uC�����`� 7�n��	��U$!	<D��:�vG�,..����K�.�2[o+����x�͞][�SNb?6��b��R'���w[7*����oh$���V�{��\o�'�A����em�J�ݰ�t���x��,�ͬp��D8�����Y�AP�ߋңi�e=���[�:��*gJ�
Gz�<MT_D�¬hb�qvf�qDbN��j��Պv���+w�AM�*a5��0		W���.�@��]�˔4�\r�2l��y���6� �~=�%0�;X�\8&2gS���aU�;���H�q�F[	E�O/�3h��.�99����OS��-�#��&s���!ijzM�Q\
Fp \�鞇�g�ᣌ����m�r[œ��W�m���Y��%�P'9=E��j�/�0��<pe$���&�G�FM�$7�a>������a�akʛ��]_N���'C\�*��z�Y ҟ�k���e�Ι��>�2�l�>��M�3m��.�T�`CA"�¦ �'v�c?��+�a�nk��B��~�Vv�1 .ڄ�-�N����_7�@�%��7/��6�b�o���/�� �n 9J(�ƺt�̩<'���������oR%���;��p�)42.�ѬF��TY|;�2�[gs�4�;!���2p2���s���`��h�3����Oo�.�Wt����.Brny���^�e����+ �$��[�X��������C�up,�"���Ht�߫�\�:��Ő�����H������n(����dZY��f��~��|"������W�aҔ+&8��8�λ�ͥ^�u��f������1y/r�Ө�XG�w���ņ��y.�Vuml�=����7���R��q��p/<ev����P׎�����O����¢�@7�5�G�8?�-�bG�-~h:i�l)�`|j��R�,
vD;�xr�W��H���*��q�r�,'8
����HU0F(~�r	A��9 �3��5eDh��!0�]�Ntky�i�
q`��+����i��^�z�&e�s�(�˾����/i-U6����>��n�������9}k؟~��@�|��C@EC�i���1��7�\�Ruܠ�6�y���4��b�5�B��!��Ǭ_��#�8�K�a��n}��|���G\v��Ň$�	hʣ�c��ǈbZ�C�@ �e��X+�\qN�͡���-��e�P�E}�|:�{���25ra�nA����6i�3�W��ˢ �@��E����A6.��l���Ѭ~v<�v���VG}䮦��c>h̡3m�A<�$��0��}��}<��
��%���P����`r7E�;�x���h��#-\�y	��H��MfN��Aޯ��u�ӇW����&̛�)��D	L�Ģ9ڧI�b��@۳9E4-����]RC� ;���Csp��n
��Y��ækg�f�b��8��0��]�;jS�